module Reservation_Station(
  input          clock,
  input          reset,
  input          io_i_dispatch_packs_0_valid,
  input  [31:0]  io_i_dispatch_packs_0_pc,
  input  [31:0]  io_i_dispatch_packs_0_inst,
  input  [6:0]   io_i_dispatch_packs_0_func_code,
  input          io_i_dispatch_packs_0_branch_predict_pack_valid,
  input  [63:0]  io_i_dispatch_packs_0_branch_predict_pack_target,
  input  [3:0]   io_i_dispatch_packs_0_branch_predict_pack_branch_type,
  input          io_i_dispatch_packs_0_branch_predict_pack_select,
  input          io_i_dispatch_packs_0_branch_predict_pack_taken,
  input  [6:0]   io_i_dispatch_packs_0_phy_dst,
  input  [6:0]   io_i_dispatch_packs_0_stale_dst,
  input  [4:0]   io_i_dispatch_packs_0_arch_dst,
  input  [2:0]   io_i_dispatch_packs_0_inst_type,
  input          io_i_dispatch_packs_0_regWen,
  input          io_i_dispatch_packs_0_src1_valid,
  input  [6:0]   io_i_dispatch_packs_0_phy_rs1,
  input  [4:0]   io_i_dispatch_packs_0_arch_rs1,
  input          io_i_dispatch_packs_0_src2_valid,
  input  [6:0]   io_i_dispatch_packs_0_phy_rs2,
  input  [4:0]   io_i_dispatch_packs_0_arch_rs2,
  input  [6:0]   io_i_dispatch_packs_0_rob_idx,
  input  [63:0]  io_i_dispatch_packs_0_imm,
  input  [63:0]  io_i_dispatch_packs_0_src1_value,
  input  [63:0]  io_i_dispatch_packs_0_src2_value,
  input  [2:0]   io_i_dispatch_packs_0_op1_sel,
  input  [2:0]   io_i_dispatch_packs_0_op2_sel,
  input  [4:0]   io_i_dispatch_packs_0_alu_sel,
  input  [3:0]   io_i_dispatch_packs_0_branch_type,
  input  [1:0]   io_i_dispatch_packs_0_mem_type,
  input          io_i_dispatch_packs_1_valid,
  input  [31:0]  io_i_dispatch_packs_1_pc,
  input  [31:0]  io_i_dispatch_packs_1_inst,
  input  [6:0]   io_i_dispatch_packs_1_func_code,
  input          io_i_dispatch_packs_1_branch_predict_pack_valid,
  input  [63:0]  io_i_dispatch_packs_1_branch_predict_pack_target,
  input  [3:0]   io_i_dispatch_packs_1_branch_predict_pack_branch_type,
  input          io_i_dispatch_packs_1_branch_predict_pack_select,
  input          io_i_dispatch_packs_1_branch_predict_pack_taken,
  input  [6:0]   io_i_dispatch_packs_1_phy_dst,
  input  [6:0]   io_i_dispatch_packs_1_stale_dst,
  input  [4:0]   io_i_dispatch_packs_1_arch_dst,
  input  [2:0]   io_i_dispatch_packs_1_inst_type,
  input          io_i_dispatch_packs_1_regWen,
  input          io_i_dispatch_packs_1_src1_valid,
  input  [6:0]   io_i_dispatch_packs_1_phy_rs1,
  input  [4:0]   io_i_dispatch_packs_1_arch_rs1,
  input          io_i_dispatch_packs_1_src2_valid,
  input  [6:0]   io_i_dispatch_packs_1_phy_rs2,
  input  [4:0]   io_i_dispatch_packs_1_arch_rs2,
  input  [6:0]   io_i_dispatch_packs_1_rob_idx,
  input  [63:0]  io_i_dispatch_packs_1_imm,
  input  [63:0]  io_i_dispatch_packs_1_src1_value,
  input  [63:0]  io_i_dispatch_packs_1_src2_value,
  input  [2:0]   io_i_dispatch_packs_1_op1_sel,
  input  [2:0]   io_i_dispatch_packs_1_op2_sel,
  input  [4:0]   io_i_dispatch_packs_1_alu_sel,
  input  [3:0]   io_i_dispatch_packs_1_branch_type,
  input  [1:0]   io_i_dispatch_packs_1_mem_type,
  output         io_o_issue_packs_0_valid,
  output [31:0]  io_o_issue_packs_0_pc,
  output [31:0]  io_o_issue_packs_0_inst,
  output [6:0]   io_o_issue_packs_0_func_code,
  output         io_o_issue_packs_0_branch_predict_pack_valid,
  output [63:0]  io_o_issue_packs_0_branch_predict_pack_target,
  output [3:0]   io_o_issue_packs_0_branch_predict_pack_branch_type,
  output         io_o_issue_packs_0_branch_predict_pack_select,
  output         io_o_issue_packs_0_branch_predict_pack_taken,
  output [6:0]   io_o_issue_packs_0_phy_dst,
  output [6:0]   io_o_issue_packs_0_stale_dst,
  output [4:0]   io_o_issue_packs_0_arch_dst,
  output [2:0]   io_o_issue_packs_0_inst_type,
  output         io_o_issue_packs_0_regWen,
  output         io_o_issue_packs_0_src1_valid,
  output [6:0]   io_o_issue_packs_0_phy_rs1,
  output [4:0]   io_o_issue_packs_0_arch_rs1,
  output         io_o_issue_packs_0_src2_valid,
  output [6:0]   io_o_issue_packs_0_phy_rs2,
  output [4:0]   io_o_issue_packs_0_arch_rs2,
  output [6:0]   io_o_issue_packs_0_rob_idx,
  output [63:0]  io_o_issue_packs_0_imm,
  output [63:0]  io_o_issue_packs_0_src1_value,
  output [63:0]  io_o_issue_packs_0_src2_value,
  output [2:0]   io_o_issue_packs_0_op1_sel,
  output [2:0]   io_o_issue_packs_0_op2_sel,
  output [4:0]   io_o_issue_packs_0_alu_sel,
  output [3:0]   io_o_issue_packs_0_branch_type,
  output [1:0]   io_o_issue_packs_0_mem_type,
  output         io_o_issue_packs_1_valid,
  output [31:0]  io_o_issue_packs_1_pc,
  output [31:0]  io_o_issue_packs_1_inst,
  output [6:0]   io_o_issue_packs_1_func_code,
  output         io_o_issue_packs_1_branch_predict_pack_valid,
  output [63:0]  io_o_issue_packs_1_branch_predict_pack_target,
  output [3:0]   io_o_issue_packs_1_branch_predict_pack_branch_type,
  output         io_o_issue_packs_1_branch_predict_pack_select,
  output         io_o_issue_packs_1_branch_predict_pack_taken,
  output [6:0]   io_o_issue_packs_1_phy_dst,
  output [6:0]   io_o_issue_packs_1_stale_dst,
  output [4:0]   io_o_issue_packs_1_arch_dst,
  output [2:0]   io_o_issue_packs_1_inst_type,
  output         io_o_issue_packs_1_regWen,
  output         io_o_issue_packs_1_src1_valid,
  output [6:0]   io_o_issue_packs_1_phy_rs1,
  output [4:0]   io_o_issue_packs_1_arch_rs1,
  output         io_o_issue_packs_1_src2_valid,
  output [6:0]   io_o_issue_packs_1_phy_rs2,
  output [4:0]   io_o_issue_packs_1_arch_rs2,
  output [6:0]   io_o_issue_packs_1_rob_idx,
  output [63:0]  io_o_issue_packs_1_imm,
  output [63:0]  io_o_issue_packs_1_src1_value,
  output [63:0]  io_o_issue_packs_1_src2_value,
  output [2:0]   io_o_issue_packs_1_op1_sel,
  output [2:0]   io_o_issue_packs_1_op2_sel,
  output [4:0]   io_o_issue_packs_1_alu_sel,
  output [3:0]   io_o_issue_packs_1_branch_type,
  output [1:0]   io_o_issue_packs_1_mem_type,
  input  [127:0] io_i_wakeup_port,
  input          io_i_ex_res_packs_0_valid,
  input  [6:0]   io_i_ex_res_packs_0_uop_phy_dst,
  input  [63:0]  io_i_ex_res_packs_0_uop_dst_value,
  input          io_i_ex_res_packs_1_valid,
  input  [6:0]   io_i_ex_res_packs_1_uop_phy_dst,
  input  [63:0]  io_i_ex_res_packs_1_uop_dst_value,
  input          io_i_branch_resolve_pack_valid,
  input          io_i_branch_resolve_pack_mispred,
  input  [6:0]   io_i_branch_resolve_pack_rob_idx,
  output         io_o_full,
  input          io_i_exception,
  input          io_i_rollback_valid,
  input  [1:0]   io_i_available_funcs_0,
  input  [1:0]   io_i_available_funcs_1,
  input  [1:0]   io_i_available_funcs_2,
  input  [1:0]   io_i_available_funcs_3,
  input  [1:0]   io_i_available_funcs_4,
  input  [1:0]   io_i_available_funcs_5,
  input  [6:0]   io_i_ROB_first_entry
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  reservation_station_0_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_0_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_0_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_0_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_0_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_0_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_0_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_0_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_1_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_1_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_1_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_1_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_1_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_1_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_1_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_2_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_2_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_2_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_2_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_2_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_2_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_2_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_3_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_3_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_3_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_3_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_3_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_3_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_3_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_4_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_4_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_4_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_4_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_4_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_4_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_4_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_5_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_5_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_5_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_5_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_5_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_5_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_5_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_6_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_6_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_6_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_6_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_6_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_6_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_6_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_7_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_7_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_7_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_7_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_7_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_7_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_7_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_8_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_8_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_8_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_8_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_8_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_8_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_8_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_9_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_9_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_9_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_9_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_9_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_9_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_9_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_10_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_10_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_10_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_10_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_10_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_10_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_10_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_11_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_11_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_11_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_11_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_11_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_11_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_11_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_12_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_12_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_12_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_12_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_12_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_12_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_12_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_13_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_13_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_13_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_13_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_13_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_13_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_13_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_14_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_14_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_14_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_14_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_14_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_14_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_14_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_15_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_15_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_15_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_15_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_15_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_15_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_15_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_16_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_16_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_16_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_16_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_16_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_16_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_16_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_17_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_17_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_17_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_17_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_17_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_17_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_17_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_18_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_18_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_18_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_18_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_18_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_18_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_18_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_19_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_19_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_19_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_19_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_19_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_19_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_19_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_20_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_20_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_20_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_20_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_20_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_20_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_20_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_21_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_21_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_21_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_21_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_21_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_21_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_21_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_22_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_22_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_22_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_22_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_22_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_22_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_22_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_23_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_23_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_23_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_23_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_23_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_23_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_23_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_24_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_24_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_24_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_24_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_24_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_24_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_24_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_25_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_25_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_25_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_25_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_25_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_25_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_25_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_26_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_26_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_26_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_26_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_26_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_26_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_26_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_27_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_27_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_27_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_27_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_27_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_27_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_27_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_28_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_28_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_28_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_28_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_28_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_28_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_28_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_29_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_29_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_29_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_29_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_29_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_29_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_29_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_30_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_30_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_30_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_30_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_30_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_30_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_30_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_31_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_31_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_31_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_31_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_31_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_31_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_31_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_32_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_32_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_32_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_32_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_32_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_32_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_32_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_33_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_33_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_33_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_33_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_33_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_33_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_33_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_34_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_34_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_34_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_34_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_34_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_34_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_34_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_35_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_35_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_35_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_35_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_35_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_35_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_35_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_36_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_36_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_36_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_36_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_36_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_36_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_36_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_37_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_37_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_37_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_37_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_37_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_37_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_37_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_38_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_38_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_38_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_38_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_38_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_38_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_38_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_39_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_39_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_39_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_39_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_39_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_39_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_39_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_40_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_40_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_40_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_40_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_40_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_40_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_40_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_41_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_41_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_41_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_41_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_41_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_41_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_41_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_42_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_42_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_42_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_42_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_42_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_42_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_42_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_43_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_43_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_43_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_43_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_43_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_43_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_43_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_44_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_44_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_44_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_44_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_44_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_44_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_44_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_45_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_45_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_45_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_45_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_45_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_45_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_45_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_46_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_46_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_46_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_46_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_46_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_46_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_46_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_47_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_47_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_47_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_47_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_47_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_47_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_47_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_48_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_48_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_48_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_48_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_48_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_48_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_48_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_49_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_49_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_49_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_49_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_49_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_49_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_49_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_50_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_50_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_50_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_50_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_50_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_50_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_50_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_51_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_51_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_51_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_51_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_51_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_51_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_51_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_52_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_52_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_52_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_52_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_52_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_52_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_52_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_53_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_53_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_53_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_53_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_53_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_53_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_53_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_54_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_54_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_54_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_54_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_54_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_54_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_54_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_55_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_55_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_55_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_55_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_55_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_55_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_55_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_56_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_56_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_56_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_56_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_56_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_56_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_56_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_57_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_57_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_57_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_57_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_57_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_57_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_57_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_58_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_58_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_58_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_58_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_58_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_58_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_58_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_59_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_59_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_59_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_59_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_59_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_59_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_59_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_60_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_60_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_60_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_60_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_60_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_60_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_60_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_61_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_61_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_61_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_61_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_61_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_61_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_61_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_62_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_62_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_62_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_62_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_62_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_62_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_62_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_allocated_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_63_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_63_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_63_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_age_pack_issue_valid_0; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_age_pack_issue_valid_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_63_io_i_age_pack_max_age; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_63_io_i_age_pack_issued_ages_0; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_63_io_i_age_pack_issued_ages_1; // @[reservation_station.scala 38:51]
  wire [7:0] reservation_station_63_io_o_age; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  temp_1 = reservation_station_1_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_0 = reservation_station_0_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_3 = reservation_station_3_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_2 = reservation_station_2_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_5 = reservation_station_5_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_4 = reservation_station_4_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_7 = reservation_station_7_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_6 = reservation_station_6_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_lo_lo_lo = {temp_7,temp_6,temp_5,temp_4,temp_3,temp_2,temp_1,temp_0}; // @[reservation_station.scala 104:46]
  wire  temp_9 = reservation_station_9_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_8 = reservation_station_8_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_11 = reservation_station_11_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_10 = reservation_station_10_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_13 = reservation_station_13_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_12 = reservation_station_12_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_15 = reservation_station_15_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_14 = reservation_station_14_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [15:0] reservation_station_valid_lo_lo = {temp_15,temp_14,temp_13,temp_12,temp_11,temp_10,temp_9,temp_8,
    reservation_station_valid_lo_lo_lo}; // @[reservation_station.scala 104:46]
  wire  temp_17 = reservation_station_17_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_16 = reservation_station_16_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_19 = reservation_station_19_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_18 = reservation_station_18_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_21 = reservation_station_21_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_20 = reservation_station_20_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_23 = reservation_station_23_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_22 = reservation_station_22_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_lo_hi_lo = {temp_23,temp_22,temp_21,temp_20,temp_19,temp_18,temp_17,temp_16}; // @[reservation_station.scala 104:46]
  wire  temp_25 = reservation_station_25_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_24 = reservation_station_24_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_27 = reservation_station_27_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_26 = reservation_station_26_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_29 = reservation_station_29_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_28 = reservation_station_28_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_31 = reservation_station_31_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_30 = reservation_station_30_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [31:0] reservation_station_valid_lo = {temp_31,temp_30,temp_29,temp_28,temp_27,temp_26,temp_25,temp_24,
    reservation_station_valid_lo_hi_lo,reservation_station_valid_lo_lo}; // @[reservation_station.scala 104:46]
  wire  temp_33 = reservation_station_33_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_32 = reservation_station_32_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_35 = reservation_station_35_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_34 = reservation_station_34_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_37 = reservation_station_37_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_36 = reservation_station_36_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_39 = reservation_station_39_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_38 = reservation_station_38_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_hi_lo_lo = {temp_39,temp_38,temp_37,temp_36,temp_35,temp_34,temp_33,temp_32}; // @[reservation_station.scala 104:46]
  wire  temp_41 = reservation_station_41_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_40 = reservation_station_40_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_43 = reservation_station_43_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_42 = reservation_station_42_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_45 = reservation_station_45_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_44 = reservation_station_44_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_47 = reservation_station_47_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_46 = reservation_station_46_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [15:0] reservation_station_valid_hi_lo = {temp_47,temp_46,temp_45,temp_44,temp_43,temp_42,temp_41,temp_40,
    reservation_station_valid_hi_lo_lo}; // @[reservation_station.scala 104:46]
  wire  temp_49 = reservation_station_49_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_48 = reservation_station_48_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_51 = reservation_station_51_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_50 = reservation_station_50_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_53 = reservation_station_53_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_52 = reservation_station_52_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_55 = reservation_station_55_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_54 = reservation_station_54_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_hi_hi_lo = {temp_55,temp_54,temp_53,temp_52,temp_51,temp_50,temp_49,temp_48}; // @[reservation_station.scala 104:46]
  wire  temp_57 = reservation_station_57_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_56 = reservation_station_56_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_59 = reservation_station_59_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_58 = reservation_station_58_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_61 = reservation_station_61_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_60 = reservation_station_60_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_63 = reservation_station_63_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_62 = reservation_station_62_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [31:0] reservation_station_valid_hi = {temp_63,temp_62,temp_61,temp_60,temp_59,temp_58,temp_57,temp_56,
    reservation_station_valid_hi_hi_lo,reservation_station_valid_hi_lo}; // @[reservation_station.scala 104:46]
  wire [63:0] reservation_station_valid = {reservation_station_valid_hi,reservation_station_valid_lo}; // @[reservation_station.scala 104:46]
  wire [63:0] _write_idx1_T = ~reservation_station_valid; // @[reservation_station.scala 105:34]
  wire [5:0] _write_idx1_T_65 = _write_idx1_T[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_66 = _write_idx1_T[61] ? 6'h3d : _write_idx1_T_65; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_67 = _write_idx1_T[60] ? 6'h3c : _write_idx1_T_66; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_68 = _write_idx1_T[59] ? 6'h3b : _write_idx1_T_67; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_69 = _write_idx1_T[58] ? 6'h3a : _write_idx1_T_68; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_70 = _write_idx1_T[57] ? 6'h39 : _write_idx1_T_69; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_71 = _write_idx1_T[56] ? 6'h38 : _write_idx1_T_70; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_72 = _write_idx1_T[55] ? 6'h37 : _write_idx1_T_71; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_73 = _write_idx1_T[54] ? 6'h36 : _write_idx1_T_72; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_74 = _write_idx1_T[53] ? 6'h35 : _write_idx1_T_73; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_75 = _write_idx1_T[52] ? 6'h34 : _write_idx1_T_74; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_76 = _write_idx1_T[51] ? 6'h33 : _write_idx1_T_75; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_77 = _write_idx1_T[50] ? 6'h32 : _write_idx1_T_76; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_78 = _write_idx1_T[49] ? 6'h31 : _write_idx1_T_77; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_79 = _write_idx1_T[48] ? 6'h30 : _write_idx1_T_78; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_80 = _write_idx1_T[47] ? 6'h2f : _write_idx1_T_79; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_81 = _write_idx1_T[46] ? 6'h2e : _write_idx1_T_80; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_82 = _write_idx1_T[45] ? 6'h2d : _write_idx1_T_81; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_83 = _write_idx1_T[44] ? 6'h2c : _write_idx1_T_82; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_84 = _write_idx1_T[43] ? 6'h2b : _write_idx1_T_83; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_85 = _write_idx1_T[42] ? 6'h2a : _write_idx1_T_84; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_86 = _write_idx1_T[41] ? 6'h29 : _write_idx1_T_85; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_87 = _write_idx1_T[40] ? 6'h28 : _write_idx1_T_86; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_88 = _write_idx1_T[39] ? 6'h27 : _write_idx1_T_87; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_89 = _write_idx1_T[38] ? 6'h26 : _write_idx1_T_88; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_90 = _write_idx1_T[37] ? 6'h25 : _write_idx1_T_89; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_91 = _write_idx1_T[36] ? 6'h24 : _write_idx1_T_90; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_92 = _write_idx1_T[35] ? 6'h23 : _write_idx1_T_91; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_93 = _write_idx1_T[34] ? 6'h22 : _write_idx1_T_92; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_94 = _write_idx1_T[33] ? 6'h21 : _write_idx1_T_93; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_95 = _write_idx1_T[32] ? 6'h20 : _write_idx1_T_94; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_96 = _write_idx1_T[31] ? 6'h1f : _write_idx1_T_95; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_97 = _write_idx1_T[30] ? 6'h1e : _write_idx1_T_96; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_98 = _write_idx1_T[29] ? 6'h1d : _write_idx1_T_97; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_99 = _write_idx1_T[28] ? 6'h1c : _write_idx1_T_98; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_100 = _write_idx1_T[27] ? 6'h1b : _write_idx1_T_99; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_101 = _write_idx1_T[26] ? 6'h1a : _write_idx1_T_100; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_102 = _write_idx1_T[25] ? 6'h19 : _write_idx1_T_101; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_103 = _write_idx1_T[24] ? 6'h18 : _write_idx1_T_102; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_104 = _write_idx1_T[23] ? 6'h17 : _write_idx1_T_103; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_105 = _write_idx1_T[22] ? 6'h16 : _write_idx1_T_104; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_106 = _write_idx1_T[21] ? 6'h15 : _write_idx1_T_105; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_107 = _write_idx1_T[20] ? 6'h14 : _write_idx1_T_106; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_108 = _write_idx1_T[19] ? 6'h13 : _write_idx1_T_107; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_109 = _write_idx1_T[18] ? 6'h12 : _write_idx1_T_108; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_110 = _write_idx1_T[17] ? 6'h11 : _write_idx1_T_109; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_111 = _write_idx1_T[16] ? 6'h10 : _write_idx1_T_110; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_112 = _write_idx1_T[15] ? 6'hf : _write_idx1_T_111; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_113 = _write_idx1_T[14] ? 6'he : _write_idx1_T_112; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_114 = _write_idx1_T[13] ? 6'hd : _write_idx1_T_113; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_115 = _write_idx1_T[12] ? 6'hc : _write_idx1_T_114; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_116 = _write_idx1_T[11] ? 6'hb : _write_idx1_T_115; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_117 = _write_idx1_T[10] ? 6'ha : _write_idx1_T_116; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_118 = _write_idx1_T[9] ? 6'h9 : _write_idx1_T_117; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_119 = _write_idx1_T[8] ? 6'h8 : _write_idx1_T_118; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_120 = _write_idx1_T[7] ? 6'h7 : _write_idx1_T_119; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_121 = _write_idx1_T[6] ? 6'h6 : _write_idx1_T_120; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_122 = _write_idx1_T[5] ? 6'h5 : _write_idx1_T_121; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_123 = _write_idx1_T[4] ? 6'h4 : _write_idx1_T_122; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_124 = _write_idx1_T[3] ? 6'h3 : _write_idx1_T_123; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_125 = _write_idx1_T[2] ? 6'h2 : _write_idx1_T_124; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_126 = _write_idx1_T[1] ? 6'h1 : _write_idx1_T_125; // @[Mux.scala 47:70]
  wire [5:0] write_idx1 = _write_idx1_T[0] ? 6'h0 : _write_idx1_T_126; // @[Mux.scala 47:70]
  wire [63:0] _reservation_station_valid_withmask_T = 64'h1 << write_idx1; // @[OneHot.scala 57:35]
  wire [63:0] reservation_station_valid_withmask = reservation_station_valid | _reservation_station_valid_withmask_T; // @[reservation_station.scala 106:69]
  wire [63:0] _write_idx2_T = ~reservation_station_valid_withmask; // @[reservation_station.scala 107:34]
  wire [5:0] _write_idx2_T_65 = _write_idx2_T[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_66 = _write_idx2_T[61] ? 6'h3d : _write_idx2_T_65; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_67 = _write_idx2_T[60] ? 6'h3c : _write_idx2_T_66; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_68 = _write_idx2_T[59] ? 6'h3b : _write_idx2_T_67; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_69 = _write_idx2_T[58] ? 6'h3a : _write_idx2_T_68; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_70 = _write_idx2_T[57] ? 6'h39 : _write_idx2_T_69; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_71 = _write_idx2_T[56] ? 6'h38 : _write_idx2_T_70; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_72 = _write_idx2_T[55] ? 6'h37 : _write_idx2_T_71; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_73 = _write_idx2_T[54] ? 6'h36 : _write_idx2_T_72; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_74 = _write_idx2_T[53] ? 6'h35 : _write_idx2_T_73; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_75 = _write_idx2_T[52] ? 6'h34 : _write_idx2_T_74; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_76 = _write_idx2_T[51] ? 6'h33 : _write_idx2_T_75; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_77 = _write_idx2_T[50] ? 6'h32 : _write_idx2_T_76; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_78 = _write_idx2_T[49] ? 6'h31 : _write_idx2_T_77; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_79 = _write_idx2_T[48] ? 6'h30 : _write_idx2_T_78; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_80 = _write_idx2_T[47] ? 6'h2f : _write_idx2_T_79; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_81 = _write_idx2_T[46] ? 6'h2e : _write_idx2_T_80; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_82 = _write_idx2_T[45] ? 6'h2d : _write_idx2_T_81; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_83 = _write_idx2_T[44] ? 6'h2c : _write_idx2_T_82; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_84 = _write_idx2_T[43] ? 6'h2b : _write_idx2_T_83; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_85 = _write_idx2_T[42] ? 6'h2a : _write_idx2_T_84; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_86 = _write_idx2_T[41] ? 6'h29 : _write_idx2_T_85; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_87 = _write_idx2_T[40] ? 6'h28 : _write_idx2_T_86; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_88 = _write_idx2_T[39] ? 6'h27 : _write_idx2_T_87; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_89 = _write_idx2_T[38] ? 6'h26 : _write_idx2_T_88; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_90 = _write_idx2_T[37] ? 6'h25 : _write_idx2_T_89; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_91 = _write_idx2_T[36] ? 6'h24 : _write_idx2_T_90; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_92 = _write_idx2_T[35] ? 6'h23 : _write_idx2_T_91; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_93 = _write_idx2_T[34] ? 6'h22 : _write_idx2_T_92; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_94 = _write_idx2_T[33] ? 6'h21 : _write_idx2_T_93; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_95 = _write_idx2_T[32] ? 6'h20 : _write_idx2_T_94; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_96 = _write_idx2_T[31] ? 6'h1f : _write_idx2_T_95; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_97 = _write_idx2_T[30] ? 6'h1e : _write_idx2_T_96; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_98 = _write_idx2_T[29] ? 6'h1d : _write_idx2_T_97; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_99 = _write_idx2_T[28] ? 6'h1c : _write_idx2_T_98; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_100 = _write_idx2_T[27] ? 6'h1b : _write_idx2_T_99; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_101 = _write_idx2_T[26] ? 6'h1a : _write_idx2_T_100; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_102 = _write_idx2_T[25] ? 6'h19 : _write_idx2_T_101; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_103 = _write_idx2_T[24] ? 6'h18 : _write_idx2_T_102; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_104 = _write_idx2_T[23] ? 6'h17 : _write_idx2_T_103; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_105 = _write_idx2_T[22] ? 6'h16 : _write_idx2_T_104; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_106 = _write_idx2_T[21] ? 6'h15 : _write_idx2_T_105; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_107 = _write_idx2_T[20] ? 6'h14 : _write_idx2_T_106; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_108 = _write_idx2_T[19] ? 6'h13 : _write_idx2_T_107; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_109 = _write_idx2_T[18] ? 6'h12 : _write_idx2_T_108; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_110 = _write_idx2_T[17] ? 6'h11 : _write_idx2_T_109; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_111 = _write_idx2_T[16] ? 6'h10 : _write_idx2_T_110; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_112 = _write_idx2_T[15] ? 6'hf : _write_idx2_T_111; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_113 = _write_idx2_T[14] ? 6'he : _write_idx2_T_112; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_114 = _write_idx2_T[13] ? 6'hd : _write_idx2_T_113; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_115 = _write_idx2_T[12] ? 6'hc : _write_idx2_T_114; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_116 = _write_idx2_T[11] ? 6'hb : _write_idx2_T_115; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_117 = _write_idx2_T[10] ? 6'ha : _write_idx2_T_116; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_118 = _write_idx2_T[9] ? 6'h9 : _write_idx2_T_117; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_119 = _write_idx2_T[8] ? 6'h8 : _write_idx2_T_118; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_120 = _write_idx2_T[7] ? 6'h7 : _write_idx2_T_119; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_121 = _write_idx2_T[6] ? 6'h6 : _write_idx2_T_120; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_122 = _write_idx2_T[5] ? 6'h5 : _write_idx2_T_121; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_123 = _write_idx2_T[4] ? 6'h4 : _write_idx2_T_122; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_124 = _write_idx2_T[3] ? 6'h3 : _write_idx2_T_123; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_125 = _write_idx2_T[2] ? 6'h2 : _write_idx2_T_124; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_126 = _write_idx2_T[1] ? 6'h1 : _write_idx2_T_125; // @[Mux.scala 47:70]
  wire [5:0] write_idx2 = _write_idx2_T[0] ? 6'h0 : _write_idx2_T_126; // @[Mux.scala 47:70]
  wire  temp2_0 = |io_i_available_funcs_0; // @[reservation_station.scala 118:44]
  wire  temp2_1 = |io_i_available_funcs_1; // @[reservation_station.scala 118:44]
  wire  temp2_2 = |io_i_available_funcs_2; // @[reservation_station.scala 118:44]
  wire  temp2_3 = |io_i_available_funcs_3; // @[reservation_station.scala 118:44]
  wire  temp2_4 = |io_i_available_funcs_4; // @[reservation_station.scala 118:44]
  wire  temp2_5 = |io_i_available_funcs_5; // @[reservation_station.scala 118:44]
  wire [6:0] available_funcs = {1'h0,temp2_5,temp2_4,temp2_3,temp2_2,temp2_1,temp2_0}; // @[reservation_station.scala 120:37]
  wire [7:0] _age_considering_issue_T_1 = reservation_station_0_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_2 = ~_age_considering_issue_T_1; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_3 = reservation_station_0_io_o_age | _age_considering_issue_T_2; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_4 = reservation_station_0_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_5 = |_age_considering_issue_T_4; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_7 = _age_considering_issue_T_5 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_8 = ~_age_considering_issue_T_7; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__0 = _age_considering_issue_T_3 | _age_considering_issue_T_8; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_11 = reservation_station_1_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_12 = ~_age_considering_issue_T_11; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_13 = reservation_station_1_io_o_age | _age_considering_issue_T_12; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_14 = reservation_station_1_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_15 = |_age_considering_issue_T_14; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_17 = _age_considering_issue_T_15 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_18 = ~_age_considering_issue_T_17; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__1 = _age_considering_issue_T_13 | _age_considering_issue_T_18; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_21 = reservation_station_2_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_22 = ~_age_considering_issue_T_21; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_23 = reservation_station_2_io_o_age | _age_considering_issue_T_22; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_24 = reservation_station_2_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_25 = |_age_considering_issue_T_24; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_27 = _age_considering_issue_T_25 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_28 = ~_age_considering_issue_T_27; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__2 = _age_considering_issue_T_23 | _age_considering_issue_T_28; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_31 = reservation_station_3_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_32 = ~_age_considering_issue_T_31; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_33 = reservation_station_3_io_o_age | _age_considering_issue_T_32; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_34 = reservation_station_3_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_35 = |_age_considering_issue_T_34; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_37 = _age_considering_issue_T_35 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_38 = ~_age_considering_issue_T_37; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__3 = _age_considering_issue_T_33 | _age_considering_issue_T_38; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_41 = reservation_station_4_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_42 = ~_age_considering_issue_T_41; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_43 = reservation_station_4_io_o_age | _age_considering_issue_T_42; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_44 = reservation_station_4_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_45 = |_age_considering_issue_T_44; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_47 = _age_considering_issue_T_45 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_48 = ~_age_considering_issue_T_47; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__4 = _age_considering_issue_T_43 | _age_considering_issue_T_48; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_51 = reservation_station_5_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_52 = ~_age_considering_issue_T_51; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_53 = reservation_station_5_io_o_age | _age_considering_issue_T_52; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_54 = reservation_station_5_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_55 = |_age_considering_issue_T_54; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_57 = _age_considering_issue_T_55 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_58 = ~_age_considering_issue_T_57; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__5 = _age_considering_issue_T_53 | _age_considering_issue_T_58; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_61 = reservation_station_6_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_62 = ~_age_considering_issue_T_61; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_63 = reservation_station_6_io_o_age | _age_considering_issue_T_62; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_64 = reservation_station_6_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_65 = |_age_considering_issue_T_64; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_67 = _age_considering_issue_T_65 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_68 = ~_age_considering_issue_T_67; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__6 = _age_considering_issue_T_63 | _age_considering_issue_T_68; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_71 = reservation_station_7_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_72 = ~_age_considering_issue_T_71; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_73 = reservation_station_7_io_o_age | _age_considering_issue_T_72; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_74 = reservation_station_7_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_75 = |_age_considering_issue_T_74; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_77 = _age_considering_issue_T_75 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_78 = ~_age_considering_issue_T_77; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__7 = _age_considering_issue_T_73 | _age_considering_issue_T_78; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_81 = reservation_station_8_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_82 = ~_age_considering_issue_T_81; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_83 = reservation_station_8_io_o_age | _age_considering_issue_T_82; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_84 = reservation_station_8_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_85 = |_age_considering_issue_T_84; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_87 = _age_considering_issue_T_85 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_88 = ~_age_considering_issue_T_87; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__8 = _age_considering_issue_T_83 | _age_considering_issue_T_88; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_91 = reservation_station_9_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_92 = ~_age_considering_issue_T_91; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_93 = reservation_station_9_io_o_age | _age_considering_issue_T_92; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_94 = reservation_station_9_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_95 = |_age_considering_issue_T_94; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_97 = _age_considering_issue_T_95 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_98 = ~_age_considering_issue_T_97; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__9 = _age_considering_issue_T_93 | _age_considering_issue_T_98; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_101 = reservation_station_10_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_102 = ~_age_considering_issue_T_101; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_103 = reservation_station_10_io_o_age | _age_considering_issue_T_102; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_104 = reservation_station_10_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_105 = |_age_considering_issue_T_104; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_107 = _age_considering_issue_T_105 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_108 = ~_age_considering_issue_T_107; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__10 = _age_considering_issue_T_103 | _age_considering_issue_T_108; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_111 = reservation_station_11_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_112 = ~_age_considering_issue_T_111; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_113 = reservation_station_11_io_o_age | _age_considering_issue_T_112; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_114 = reservation_station_11_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_115 = |_age_considering_issue_T_114; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_117 = _age_considering_issue_T_115 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_118 = ~_age_considering_issue_T_117; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__11 = _age_considering_issue_T_113 | _age_considering_issue_T_118; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_121 = reservation_station_12_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_122 = ~_age_considering_issue_T_121; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_123 = reservation_station_12_io_o_age | _age_considering_issue_T_122; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_124 = reservation_station_12_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_125 = |_age_considering_issue_T_124; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_127 = _age_considering_issue_T_125 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_128 = ~_age_considering_issue_T_127; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__12 = _age_considering_issue_T_123 | _age_considering_issue_T_128; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_131 = reservation_station_13_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_132 = ~_age_considering_issue_T_131; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_133 = reservation_station_13_io_o_age | _age_considering_issue_T_132; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_134 = reservation_station_13_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_135 = |_age_considering_issue_T_134; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_137 = _age_considering_issue_T_135 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_138 = ~_age_considering_issue_T_137; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__13 = _age_considering_issue_T_133 | _age_considering_issue_T_138; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_141 = reservation_station_14_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_142 = ~_age_considering_issue_T_141; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_143 = reservation_station_14_io_o_age | _age_considering_issue_T_142; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_144 = reservation_station_14_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_145 = |_age_considering_issue_T_144; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_147 = _age_considering_issue_T_145 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_148 = ~_age_considering_issue_T_147; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__14 = _age_considering_issue_T_143 | _age_considering_issue_T_148; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_151 = reservation_station_15_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_152 = ~_age_considering_issue_T_151; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_153 = reservation_station_15_io_o_age | _age_considering_issue_T_152; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_154 = reservation_station_15_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_155 = |_age_considering_issue_T_154; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_157 = _age_considering_issue_T_155 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_158 = ~_age_considering_issue_T_157; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__15 = _age_considering_issue_T_153 | _age_considering_issue_T_158; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_161 = reservation_station_16_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_162 = ~_age_considering_issue_T_161; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_163 = reservation_station_16_io_o_age | _age_considering_issue_T_162; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_164 = reservation_station_16_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_165 = |_age_considering_issue_T_164; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_167 = _age_considering_issue_T_165 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_168 = ~_age_considering_issue_T_167; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__16 = _age_considering_issue_T_163 | _age_considering_issue_T_168; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_171 = reservation_station_17_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_172 = ~_age_considering_issue_T_171; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_173 = reservation_station_17_io_o_age | _age_considering_issue_T_172; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_174 = reservation_station_17_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_175 = |_age_considering_issue_T_174; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_177 = _age_considering_issue_T_175 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_178 = ~_age_considering_issue_T_177; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__17 = _age_considering_issue_T_173 | _age_considering_issue_T_178; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_181 = reservation_station_18_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_182 = ~_age_considering_issue_T_181; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_183 = reservation_station_18_io_o_age | _age_considering_issue_T_182; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_184 = reservation_station_18_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_185 = |_age_considering_issue_T_184; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_187 = _age_considering_issue_T_185 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_188 = ~_age_considering_issue_T_187; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__18 = _age_considering_issue_T_183 | _age_considering_issue_T_188; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_191 = reservation_station_19_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_192 = ~_age_considering_issue_T_191; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_193 = reservation_station_19_io_o_age | _age_considering_issue_T_192; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_194 = reservation_station_19_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_195 = |_age_considering_issue_T_194; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_197 = _age_considering_issue_T_195 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_198 = ~_age_considering_issue_T_197; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__19 = _age_considering_issue_T_193 | _age_considering_issue_T_198; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_201 = reservation_station_20_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_202 = ~_age_considering_issue_T_201; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_203 = reservation_station_20_io_o_age | _age_considering_issue_T_202; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_204 = reservation_station_20_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_205 = |_age_considering_issue_T_204; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_207 = _age_considering_issue_T_205 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_208 = ~_age_considering_issue_T_207; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__20 = _age_considering_issue_T_203 | _age_considering_issue_T_208; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_211 = reservation_station_21_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_212 = ~_age_considering_issue_T_211; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_213 = reservation_station_21_io_o_age | _age_considering_issue_T_212; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_214 = reservation_station_21_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_215 = |_age_considering_issue_T_214; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_217 = _age_considering_issue_T_215 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_218 = ~_age_considering_issue_T_217; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__21 = _age_considering_issue_T_213 | _age_considering_issue_T_218; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_221 = reservation_station_22_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_222 = ~_age_considering_issue_T_221; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_223 = reservation_station_22_io_o_age | _age_considering_issue_T_222; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_224 = reservation_station_22_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_225 = |_age_considering_issue_T_224; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_227 = _age_considering_issue_T_225 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_228 = ~_age_considering_issue_T_227; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__22 = _age_considering_issue_T_223 | _age_considering_issue_T_228; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_231 = reservation_station_23_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_232 = ~_age_considering_issue_T_231; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_233 = reservation_station_23_io_o_age | _age_considering_issue_T_232; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_234 = reservation_station_23_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_235 = |_age_considering_issue_T_234; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_237 = _age_considering_issue_T_235 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_238 = ~_age_considering_issue_T_237; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__23 = _age_considering_issue_T_233 | _age_considering_issue_T_238; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_241 = reservation_station_24_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_242 = ~_age_considering_issue_T_241; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_243 = reservation_station_24_io_o_age | _age_considering_issue_T_242; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_244 = reservation_station_24_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_245 = |_age_considering_issue_T_244; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_247 = _age_considering_issue_T_245 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_248 = ~_age_considering_issue_T_247; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__24 = _age_considering_issue_T_243 | _age_considering_issue_T_248; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_251 = reservation_station_25_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_252 = ~_age_considering_issue_T_251; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_253 = reservation_station_25_io_o_age | _age_considering_issue_T_252; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_254 = reservation_station_25_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_255 = |_age_considering_issue_T_254; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_257 = _age_considering_issue_T_255 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_258 = ~_age_considering_issue_T_257; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__25 = _age_considering_issue_T_253 | _age_considering_issue_T_258; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_261 = reservation_station_26_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_262 = ~_age_considering_issue_T_261; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_263 = reservation_station_26_io_o_age | _age_considering_issue_T_262; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_264 = reservation_station_26_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_265 = |_age_considering_issue_T_264; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_267 = _age_considering_issue_T_265 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_268 = ~_age_considering_issue_T_267; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__26 = _age_considering_issue_T_263 | _age_considering_issue_T_268; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_271 = reservation_station_27_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_272 = ~_age_considering_issue_T_271; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_273 = reservation_station_27_io_o_age | _age_considering_issue_T_272; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_274 = reservation_station_27_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_275 = |_age_considering_issue_T_274; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_277 = _age_considering_issue_T_275 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_278 = ~_age_considering_issue_T_277; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__27 = _age_considering_issue_T_273 | _age_considering_issue_T_278; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_281 = reservation_station_28_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_282 = ~_age_considering_issue_T_281; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_283 = reservation_station_28_io_o_age | _age_considering_issue_T_282; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_284 = reservation_station_28_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_285 = |_age_considering_issue_T_284; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_287 = _age_considering_issue_T_285 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_288 = ~_age_considering_issue_T_287; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__28 = _age_considering_issue_T_283 | _age_considering_issue_T_288; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_291 = reservation_station_29_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_292 = ~_age_considering_issue_T_291; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_293 = reservation_station_29_io_o_age | _age_considering_issue_T_292; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_294 = reservation_station_29_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_295 = |_age_considering_issue_T_294; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_297 = _age_considering_issue_T_295 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_298 = ~_age_considering_issue_T_297; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__29 = _age_considering_issue_T_293 | _age_considering_issue_T_298; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_301 = reservation_station_30_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_302 = ~_age_considering_issue_T_301; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_303 = reservation_station_30_io_o_age | _age_considering_issue_T_302; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_304 = reservation_station_30_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_305 = |_age_considering_issue_T_304; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_307 = _age_considering_issue_T_305 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_308 = ~_age_considering_issue_T_307; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__30 = _age_considering_issue_T_303 | _age_considering_issue_T_308; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_311 = reservation_station_31_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_312 = ~_age_considering_issue_T_311; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_313 = reservation_station_31_io_o_age | _age_considering_issue_T_312; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_314 = reservation_station_31_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_315 = |_age_considering_issue_T_314; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_317 = _age_considering_issue_T_315 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_318 = ~_age_considering_issue_T_317; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__31 = _age_considering_issue_T_313 | _age_considering_issue_T_318; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_321 = reservation_station_32_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_322 = ~_age_considering_issue_T_321; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_323 = reservation_station_32_io_o_age | _age_considering_issue_T_322; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_324 = reservation_station_32_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_325 = |_age_considering_issue_T_324; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_327 = _age_considering_issue_T_325 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_328 = ~_age_considering_issue_T_327; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__32 = _age_considering_issue_T_323 | _age_considering_issue_T_328; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_331 = reservation_station_33_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_332 = ~_age_considering_issue_T_331; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_333 = reservation_station_33_io_o_age | _age_considering_issue_T_332; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_334 = reservation_station_33_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_335 = |_age_considering_issue_T_334; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_337 = _age_considering_issue_T_335 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_338 = ~_age_considering_issue_T_337; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__33 = _age_considering_issue_T_333 | _age_considering_issue_T_338; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_341 = reservation_station_34_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_342 = ~_age_considering_issue_T_341; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_343 = reservation_station_34_io_o_age | _age_considering_issue_T_342; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_344 = reservation_station_34_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_345 = |_age_considering_issue_T_344; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_347 = _age_considering_issue_T_345 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_348 = ~_age_considering_issue_T_347; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__34 = _age_considering_issue_T_343 | _age_considering_issue_T_348; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_351 = reservation_station_35_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_352 = ~_age_considering_issue_T_351; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_353 = reservation_station_35_io_o_age | _age_considering_issue_T_352; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_354 = reservation_station_35_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_355 = |_age_considering_issue_T_354; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_357 = _age_considering_issue_T_355 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_358 = ~_age_considering_issue_T_357; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__35 = _age_considering_issue_T_353 | _age_considering_issue_T_358; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_361 = reservation_station_36_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_362 = ~_age_considering_issue_T_361; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_363 = reservation_station_36_io_o_age | _age_considering_issue_T_362; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_364 = reservation_station_36_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_365 = |_age_considering_issue_T_364; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_367 = _age_considering_issue_T_365 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_368 = ~_age_considering_issue_T_367; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__36 = _age_considering_issue_T_363 | _age_considering_issue_T_368; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_371 = reservation_station_37_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_372 = ~_age_considering_issue_T_371; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_373 = reservation_station_37_io_o_age | _age_considering_issue_T_372; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_374 = reservation_station_37_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_375 = |_age_considering_issue_T_374; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_377 = _age_considering_issue_T_375 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_378 = ~_age_considering_issue_T_377; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__37 = _age_considering_issue_T_373 | _age_considering_issue_T_378; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_381 = reservation_station_38_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_382 = ~_age_considering_issue_T_381; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_383 = reservation_station_38_io_o_age | _age_considering_issue_T_382; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_384 = reservation_station_38_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_385 = |_age_considering_issue_T_384; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_387 = _age_considering_issue_T_385 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_388 = ~_age_considering_issue_T_387; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__38 = _age_considering_issue_T_383 | _age_considering_issue_T_388; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_391 = reservation_station_39_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_392 = ~_age_considering_issue_T_391; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_393 = reservation_station_39_io_o_age | _age_considering_issue_T_392; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_394 = reservation_station_39_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_395 = |_age_considering_issue_T_394; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_397 = _age_considering_issue_T_395 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_398 = ~_age_considering_issue_T_397; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__39 = _age_considering_issue_T_393 | _age_considering_issue_T_398; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_401 = reservation_station_40_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_402 = ~_age_considering_issue_T_401; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_403 = reservation_station_40_io_o_age | _age_considering_issue_T_402; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_404 = reservation_station_40_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_405 = |_age_considering_issue_T_404; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_407 = _age_considering_issue_T_405 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_408 = ~_age_considering_issue_T_407; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__40 = _age_considering_issue_T_403 | _age_considering_issue_T_408; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_411 = reservation_station_41_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_412 = ~_age_considering_issue_T_411; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_413 = reservation_station_41_io_o_age | _age_considering_issue_T_412; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_414 = reservation_station_41_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_415 = |_age_considering_issue_T_414; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_417 = _age_considering_issue_T_415 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_418 = ~_age_considering_issue_T_417; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__41 = _age_considering_issue_T_413 | _age_considering_issue_T_418; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_421 = reservation_station_42_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_422 = ~_age_considering_issue_T_421; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_423 = reservation_station_42_io_o_age | _age_considering_issue_T_422; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_424 = reservation_station_42_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_425 = |_age_considering_issue_T_424; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_427 = _age_considering_issue_T_425 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_428 = ~_age_considering_issue_T_427; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__42 = _age_considering_issue_T_423 | _age_considering_issue_T_428; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_431 = reservation_station_43_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_432 = ~_age_considering_issue_T_431; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_433 = reservation_station_43_io_o_age | _age_considering_issue_T_432; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_434 = reservation_station_43_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_435 = |_age_considering_issue_T_434; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_437 = _age_considering_issue_T_435 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_438 = ~_age_considering_issue_T_437; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__43 = _age_considering_issue_T_433 | _age_considering_issue_T_438; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_441 = reservation_station_44_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_442 = ~_age_considering_issue_T_441; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_443 = reservation_station_44_io_o_age | _age_considering_issue_T_442; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_444 = reservation_station_44_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_445 = |_age_considering_issue_T_444; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_447 = _age_considering_issue_T_445 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_448 = ~_age_considering_issue_T_447; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__44 = _age_considering_issue_T_443 | _age_considering_issue_T_448; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_451 = reservation_station_45_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_452 = ~_age_considering_issue_T_451; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_453 = reservation_station_45_io_o_age | _age_considering_issue_T_452; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_454 = reservation_station_45_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_455 = |_age_considering_issue_T_454; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_457 = _age_considering_issue_T_455 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_458 = ~_age_considering_issue_T_457; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__45 = _age_considering_issue_T_453 | _age_considering_issue_T_458; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_461 = reservation_station_46_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_462 = ~_age_considering_issue_T_461; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_463 = reservation_station_46_io_o_age | _age_considering_issue_T_462; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_464 = reservation_station_46_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_465 = |_age_considering_issue_T_464; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_467 = _age_considering_issue_T_465 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_468 = ~_age_considering_issue_T_467; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__46 = _age_considering_issue_T_463 | _age_considering_issue_T_468; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_471 = reservation_station_47_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_472 = ~_age_considering_issue_T_471; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_473 = reservation_station_47_io_o_age | _age_considering_issue_T_472; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_474 = reservation_station_47_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_475 = |_age_considering_issue_T_474; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_477 = _age_considering_issue_T_475 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_478 = ~_age_considering_issue_T_477; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__47 = _age_considering_issue_T_473 | _age_considering_issue_T_478; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_481 = reservation_station_48_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_482 = ~_age_considering_issue_T_481; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_483 = reservation_station_48_io_o_age | _age_considering_issue_T_482; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_484 = reservation_station_48_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_485 = |_age_considering_issue_T_484; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_487 = _age_considering_issue_T_485 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_488 = ~_age_considering_issue_T_487; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__48 = _age_considering_issue_T_483 | _age_considering_issue_T_488; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_491 = reservation_station_49_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_492 = ~_age_considering_issue_T_491; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_493 = reservation_station_49_io_o_age | _age_considering_issue_T_492; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_494 = reservation_station_49_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_495 = |_age_considering_issue_T_494; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_497 = _age_considering_issue_T_495 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_498 = ~_age_considering_issue_T_497; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__49 = _age_considering_issue_T_493 | _age_considering_issue_T_498; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_501 = reservation_station_50_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_502 = ~_age_considering_issue_T_501; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_503 = reservation_station_50_io_o_age | _age_considering_issue_T_502; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_504 = reservation_station_50_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_505 = |_age_considering_issue_T_504; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_507 = _age_considering_issue_T_505 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_508 = ~_age_considering_issue_T_507; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__50 = _age_considering_issue_T_503 | _age_considering_issue_T_508; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_511 = reservation_station_51_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_512 = ~_age_considering_issue_T_511; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_513 = reservation_station_51_io_o_age | _age_considering_issue_T_512; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_514 = reservation_station_51_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_515 = |_age_considering_issue_T_514; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_517 = _age_considering_issue_T_515 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_518 = ~_age_considering_issue_T_517; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__51 = _age_considering_issue_T_513 | _age_considering_issue_T_518; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_521 = reservation_station_52_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_522 = ~_age_considering_issue_T_521; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_523 = reservation_station_52_io_o_age | _age_considering_issue_T_522; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_524 = reservation_station_52_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_525 = |_age_considering_issue_T_524; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_527 = _age_considering_issue_T_525 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_528 = ~_age_considering_issue_T_527; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__52 = _age_considering_issue_T_523 | _age_considering_issue_T_528; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_531 = reservation_station_53_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_532 = ~_age_considering_issue_T_531; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_533 = reservation_station_53_io_o_age | _age_considering_issue_T_532; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_534 = reservation_station_53_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_535 = |_age_considering_issue_T_534; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_537 = _age_considering_issue_T_535 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_538 = ~_age_considering_issue_T_537; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__53 = _age_considering_issue_T_533 | _age_considering_issue_T_538; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_541 = reservation_station_54_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_542 = ~_age_considering_issue_T_541; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_543 = reservation_station_54_io_o_age | _age_considering_issue_T_542; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_544 = reservation_station_54_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_545 = |_age_considering_issue_T_544; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_547 = _age_considering_issue_T_545 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_548 = ~_age_considering_issue_T_547; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__54 = _age_considering_issue_T_543 | _age_considering_issue_T_548; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_551 = reservation_station_55_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_552 = ~_age_considering_issue_T_551; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_553 = reservation_station_55_io_o_age | _age_considering_issue_T_552; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_554 = reservation_station_55_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_555 = |_age_considering_issue_T_554; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_557 = _age_considering_issue_T_555 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_558 = ~_age_considering_issue_T_557; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__55 = _age_considering_issue_T_553 | _age_considering_issue_T_558; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_561 = reservation_station_56_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_562 = ~_age_considering_issue_T_561; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_563 = reservation_station_56_io_o_age | _age_considering_issue_T_562; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_564 = reservation_station_56_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_565 = |_age_considering_issue_T_564; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_567 = _age_considering_issue_T_565 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_568 = ~_age_considering_issue_T_567; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__56 = _age_considering_issue_T_563 | _age_considering_issue_T_568; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_571 = reservation_station_57_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_572 = ~_age_considering_issue_T_571; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_573 = reservation_station_57_io_o_age | _age_considering_issue_T_572; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_574 = reservation_station_57_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_575 = |_age_considering_issue_T_574; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_577 = _age_considering_issue_T_575 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_578 = ~_age_considering_issue_T_577; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__57 = _age_considering_issue_T_573 | _age_considering_issue_T_578; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_581 = reservation_station_58_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_582 = ~_age_considering_issue_T_581; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_583 = reservation_station_58_io_o_age | _age_considering_issue_T_582; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_584 = reservation_station_58_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_585 = |_age_considering_issue_T_584; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_587 = _age_considering_issue_T_585 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_588 = ~_age_considering_issue_T_587; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__58 = _age_considering_issue_T_583 | _age_considering_issue_T_588; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_591 = reservation_station_59_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_592 = ~_age_considering_issue_T_591; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_593 = reservation_station_59_io_o_age | _age_considering_issue_T_592; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_594 = reservation_station_59_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_595 = |_age_considering_issue_T_594; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_597 = _age_considering_issue_T_595 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_598 = ~_age_considering_issue_T_597; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__59 = _age_considering_issue_T_593 | _age_considering_issue_T_598; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_601 = reservation_station_60_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_602 = ~_age_considering_issue_T_601; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_603 = reservation_station_60_io_o_age | _age_considering_issue_T_602; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_604 = reservation_station_60_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_605 = |_age_considering_issue_T_604; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_607 = _age_considering_issue_T_605 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_608 = ~_age_considering_issue_T_607; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__60 = _age_considering_issue_T_603 | _age_considering_issue_T_608; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_611 = reservation_station_61_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_612 = ~_age_considering_issue_T_611; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_613 = reservation_station_61_io_o_age | _age_considering_issue_T_612; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_614 = reservation_station_61_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_615 = |_age_considering_issue_T_614; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_617 = _age_considering_issue_T_615 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_618 = ~_age_considering_issue_T_617; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__61 = _age_considering_issue_T_613 | _age_considering_issue_T_618; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_621 = reservation_station_62_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_622 = ~_age_considering_issue_T_621; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_623 = reservation_station_62_io_o_age | _age_considering_issue_T_622; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_624 = reservation_station_62_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_625 = |_age_considering_issue_T_624; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_627 = _age_considering_issue_T_625 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_628 = ~_age_considering_issue_T_627; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__62 = _age_considering_issue_T_623 | _age_considering_issue_T_628; // @[reservation_station.scala 123:9]
  wire [7:0] _age_considering_issue_T_631 = reservation_station_63_io_o_ready_to_issue ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_632 = ~_age_considering_issue_T_631; // @[reservation_station.scala 122:96]
  wire [7:0] _age_considering_issue_T_633 = reservation_station_63_io_o_age | _age_considering_issue_T_632; // @[reservation_station.scala 122:93]
  wire [6:0] _age_considering_issue_T_634 = reservation_station_63_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 123:63]
  wire  _age_considering_issue_T_635 = |_age_considering_issue_T_634; // @[reservation_station.scala 123:82]
  wire [7:0] _age_considering_issue_T_637 = _age_considering_issue_T_635 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_T_638 = ~_age_considering_issue_T_637; // @[reservation_station.scala 123:11]
  wire [7:0] age_considering_issue__63 = _age_considering_issue_T_633 | _age_considering_issue_T_638; // @[reservation_station.scala 123:9]
  wire [5:0] _issue1_idx_T_1 = age_considering_issue__0 < age_considering_issue__1 ? 6'h0 : 6'h1; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_3 = age_considering_issue__0 < age_considering_issue__1 ? age_considering_issue__0 :
    age_considering_issue__1; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_5 = _issue1_idx_T_3 < age_considering_issue__2 ? _issue1_idx_T_1 : 6'h2; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_7 = _issue1_idx_T_3 < age_considering_issue__2 ? _issue1_idx_T_3 : age_considering_issue__2; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_9 = _issue1_idx_T_7 < age_considering_issue__3 ? _issue1_idx_T_5 : 6'h3; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_11 = _issue1_idx_T_7 < age_considering_issue__3 ? _issue1_idx_T_7 : age_considering_issue__3; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_13 = _issue1_idx_T_11 < age_considering_issue__4 ? _issue1_idx_T_9 : 6'h4; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_15 = _issue1_idx_T_11 < age_considering_issue__4 ? _issue1_idx_T_11 :
    age_considering_issue__4; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_17 = _issue1_idx_T_15 < age_considering_issue__5 ? _issue1_idx_T_13 : 6'h5; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_19 = _issue1_idx_T_15 < age_considering_issue__5 ? _issue1_idx_T_15 :
    age_considering_issue__5; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_21 = _issue1_idx_T_19 < age_considering_issue__6 ? _issue1_idx_T_17 : 6'h6; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_23 = _issue1_idx_T_19 < age_considering_issue__6 ? _issue1_idx_T_19 :
    age_considering_issue__6; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_25 = _issue1_idx_T_23 < age_considering_issue__7 ? _issue1_idx_T_21 : 6'h7; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_27 = _issue1_idx_T_23 < age_considering_issue__7 ? _issue1_idx_T_23 :
    age_considering_issue__7; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_29 = _issue1_idx_T_27 < age_considering_issue__8 ? _issue1_idx_T_25 : 6'h8; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_31 = _issue1_idx_T_27 < age_considering_issue__8 ? _issue1_idx_T_27 :
    age_considering_issue__8; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_33 = _issue1_idx_T_31 < age_considering_issue__9 ? _issue1_idx_T_29 : 6'h9; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_35 = _issue1_idx_T_31 < age_considering_issue__9 ? _issue1_idx_T_31 :
    age_considering_issue__9; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_37 = _issue1_idx_T_35 < age_considering_issue__10 ? _issue1_idx_T_33 : 6'ha; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_39 = _issue1_idx_T_35 < age_considering_issue__10 ? _issue1_idx_T_35 :
    age_considering_issue__10; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_41 = _issue1_idx_T_39 < age_considering_issue__11 ? _issue1_idx_T_37 : 6'hb; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_43 = _issue1_idx_T_39 < age_considering_issue__11 ? _issue1_idx_T_39 :
    age_considering_issue__11; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_45 = _issue1_idx_T_43 < age_considering_issue__12 ? _issue1_idx_T_41 : 6'hc; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_47 = _issue1_idx_T_43 < age_considering_issue__12 ? _issue1_idx_T_43 :
    age_considering_issue__12; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_49 = _issue1_idx_T_47 < age_considering_issue__13 ? _issue1_idx_T_45 : 6'hd; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_51 = _issue1_idx_T_47 < age_considering_issue__13 ? _issue1_idx_T_47 :
    age_considering_issue__13; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_53 = _issue1_idx_T_51 < age_considering_issue__14 ? _issue1_idx_T_49 : 6'he; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_55 = _issue1_idx_T_51 < age_considering_issue__14 ? _issue1_idx_T_51 :
    age_considering_issue__14; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_57 = _issue1_idx_T_55 < age_considering_issue__15 ? _issue1_idx_T_53 : 6'hf; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_59 = _issue1_idx_T_55 < age_considering_issue__15 ? _issue1_idx_T_55 :
    age_considering_issue__15; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_61 = _issue1_idx_T_59 < age_considering_issue__16 ? _issue1_idx_T_57 : 6'h10; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_63 = _issue1_idx_T_59 < age_considering_issue__16 ? _issue1_idx_T_59 :
    age_considering_issue__16; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_65 = _issue1_idx_T_63 < age_considering_issue__17 ? _issue1_idx_T_61 : 6'h11; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_67 = _issue1_idx_T_63 < age_considering_issue__17 ? _issue1_idx_T_63 :
    age_considering_issue__17; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_69 = _issue1_idx_T_67 < age_considering_issue__18 ? _issue1_idx_T_65 : 6'h12; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_71 = _issue1_idx_T_67 < age_considering_issue__18 ? _issue1_idx_T_67 :
    age_considering_issue__18; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_73 = _issue1_idx_T_71 < age_considering_issue__19 ? _issue1_idx_T_69 : 6'h13; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_75 = _issue1_idx_T_71 < age_considering_issue__19 ? _issue1_idx_T_71 :
    age_considering_issue__19; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_77 = _issue1_idx_T_75 < age_considering_issue__20 ? _issue1_idx_T_73 : 6'h14; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_79 = _issue1_idx_T_75 < age_considering_issue__20 ? _issue1_idx_T_75 :
    age_considering_issue__20; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_81 = _issue1_idx_T_79 < age_considering_issue__21 ? _issue1_idx_T_77 : 6'h15; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_83 = _issue1_idx_T_79 < age_considering_issue__21 ? _issue1_idx_T_79 :
    age_considering_issue__21; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_85 = _issue1_idx_T_83 < age_considering_issue__22 ? _issue1_idx_T_81 : 6'h16; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_87 = _issue1_idx_T_83 < age_considering_issue__22 ? _issue1_idx_T_83 :
    age_considering_issue__22; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_89 = _issue1_idx_T_87 < age_considering_issue__23 ? _issue1_idx_T_85 : 6'h17; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_91 = _issue1_idx_T_87 < age_considering_issue__23 ? _issue1_idx_T_87 :
    age_considering_issue__23; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_93 = _issue1_idx_T_91 < age_considering_issue__24 ? _issue1_idx_T_89 : 6'h18; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_95 = _issue1_idx_T_91 < age_considering_issue__24 ? _issue1_idx_T_91 :
    age_considering_issue__24; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_97 = _issue1_idx_T_95 < age_considering_issue__25 ? _issue1_idx_T_93 : 6'h19; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_99 = _issue1_idx_T_95 < age_considering_issue__25 ? _issue1_idx_T_95 :
    age_considering_issue__25; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_101 = _issue1_idx_T_99 < age_considering_issue__26 ? _issue1_idx_T_97 : 6'h1a; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_103 = _issue1_idx_T_99 < age_considering_issue__26 ? _issue1_idx_T_99 :
    age_considering_issue__26; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_105 = _issue1_idx_T_103 < age_considering_issue__27 ? _issue1_idx_T_101 : 6'h1b; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_107 = _issue1_idx_T_103 < age_considering_issue__27 ? _issue1_idx_T_103 :
    age_considering_issue__27; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_109 = _issue1_idx_T_107 < age_considering_issue__28 ? _issue1_idx_T_105 : 6'h1c; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_111 = _issue1_idx_T_107 < age_considering_issue__28 ? _issue1_idx_T_107 :
    age_considering_issue__28; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_113 = _issue1_idx_T_111 < age_considering_issue__29 ? _issue1_idx_T_109 : 6'h1d; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_115 = _issue1_idx_T_111 < age_considering_issue__29 ? _issue1_idx_T_111 :
    age_considering_issue__29; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_117 = _issue1_idx_T_115 < age_considering_issue__30 ? _issue1_idx_T_113 : 6'h1e; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_119 = _issue1_idx_T_115 < age_considering_issue__30 ? _issue1_idx_T_115 :
    age_considering_issue__30; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_121 = _issue1_idx_T_119 < age_considering_issue__31 ? _issue1_idx_T_117 : 6'h1f; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_123 = _issue1_idx_T_119 < age_considering_issue__31 ? _issue1_idx_T_119 :
    age_considering_issue__31; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_125 = _issue1_idx_T_123 < age_considering_issue__32 ? _issue1_idx_T_121 : 6'h20; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_127 = _issue1_idx_T_123 < age_considering_issue__32 ? _issue1_idx_T_123 :
    age_considering_issue__32; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_129 = _issue1_idx_T_127 < age_considering_issue__33 ? _issue1_idx_T_125 : 6'h21; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_131 = _issue1_idx_T_127 < age_considering_issue__33 ? _issue1_idx_T_127 :
    age_considering_issue__33; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_133 = _issue1_idx_T_131 < age_considering_issue__34 ? _issue1_idx_T_129 : 6'h22; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_135 = _issue1_idx_T_131 < age_considering_issue__34 ? _issue1_idx_T_131 :
    age_considering_issue__34; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_137 = _issue1_idx_T_135 < age_considering_issue__35 ? _issue1_idx_T_133 : 6'h23; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_139 = _issue1_idx_T_135 < age_considering_issue__35 ? _issue1_idx_T_135 :
    age_considering_issue__35; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_141 = _issue1_idx_T_139 < age_considering_issue__36 ? _issue1_idx_T_137 : 6'h24; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_143 = _issue1_idx_T_139 < age_considering_issue__36 ? _issue1_idx_T_139 :
    age_considering_issue__36; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_145 = _issue1_idx_T_143 < age_considering_issue__37 ? _issue1_idx_T_141 : 6'h25; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_147 = _issue1_idx_T_143 < age_considering_issue__37 ? _issue1_idx_T_143 :
    age_considering_issue__37; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_149 = _issue1_idx_T_147 < age_considering_issue__38 ? _issue1_idx_T_145 : 6'h26; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_151 = _issue1_idx_T_147 < age_considering_issue__38 ? _issue1_idx_T_147 :
    age_considering_issue__38; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_153 = _issue1_idx_T_151 < age_considering_issue__39 ? _issue1_idx_T_149 : 6'h27; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_155 = _issue1_idx_T_151 < age_considering_issue__39 ? _issue1_idx_T_151 :
    age_considering_issue__39; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_157 = _issue1_idx_T_155 < age_considering_issue__40 ? _issue1_idx_T_153 : 6'h28; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_159 = _issue1_idx_T_155 < age_considering_issue__40 ? _issue1_idx_T_155 :
    age_considering_issue__40; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_161 = _issue1_idx_T_159 < age_considering_issue__41 ? _issue1_idx_T_157 : 6'h29; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_163 = _issue1_idx_T_159 < age_considering_issue__41 ? _issue1_idx_T_159 :
    age_considering_issue__41; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_165 = _issue1_idx_T_163 < age_considering_issue__42 ? _issue1_idx_T_161 : 6'h2a; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_167 = _issue1_idx_T_163 < age_considering_issue__42 ? _issue1_idx_T_163 :
    age_considering_issue__42; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_169 = _issue1_idx_T_167 < age_considering_issue__43 ? _issue1_idx_T_165 : 6'h2b; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_171 = _issue1_idx_T_167 < age_considering_issue__43 ? _issue1_idx_T_167 :
    age_considering_issue__43; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_173 = _issue1_idx_T_171 < age_considering_issue__44 ? _issue1_idx_T_169 : 6'h2c; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_175 = _issue1_idx_T_171 < age_considering_issue__44 ? _issue1_idx_T_171 :
    age_considering_issue__44; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_177 = _issue1_idx_T_175 < age_considering_issue__45 ? _issue1_idx_T_173 : 6'h2d; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_179 = _issue1_idx_T_175 < age_considering_issue__45 ? _issue1_idx_T_175 :
    age_considering_issue__45; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_181 = _issue1_idx_T_179 < age_considering_issue__46 ? _issue1_idx_T_177 : 6'h2e; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_183 = _issue1_idx_T_179 < age_considering_issue__46 ? _issue1_idx_T_179 :
    age_considering_issue__46; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_185 = _issue1_idx_T_183 < age_considering_issue__47 ? _issue1_idx_T_181 : 6'h2f; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_187 = _issue1_idx_T_183 < age_considering_issue__47 ? _issue1_idx_T_183 :
    age_considering_issue__47; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_189 = _issue1_idx_T_187 < age_considering_issue__48 ? _issue1_idx_T_185 : 6'h30; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_191 = _issue1_idx_T_187 < age_considering_issue__48 ? _issue1_idx_T_187 :
    age_considering_issue__48; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_193 = _issue1_idx_T_191 < age_considering_issue__49 ? _issue1_idx_T_189 : 6'h31; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_195 = _issue1_idx_T_191 < age_considering_issue__49 ? _issue1_idx_T_191 :
    age_considering_issue__49; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_197 = _issue1_idx_T_195 < age_considering_issue__50 ? _issue1_idx_T_193 : 6'h32; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_199 = _issue1_idx_T_195 < age_considering_issue__50 ? _issue1_idx_T_195 :
    age_considering_issue__50; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_201 = _issue1_idx_T_199 < age_considering_issue__51 ? _issue1_idx_T_197 : 6'h33; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_203 = _issue1_idx_T_199 < age_considering_issue__51 ? _issue1_idx_T_199 :
    age_considering_issue__51; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_205 = _issue1_idx_T_203 < age_considering_issue__52 ? _issue1_idx_T_201 : 6'h34; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_207 = _issue1_idx_T_203 < age_considering_issue__52 ? _issue1_idx_T_203 :
    age_considering_issue__52; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_209 = _issue1_idx_T_207 < age_considering_issue__53 ? _issue1_idx_T_205 : 6'h35; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_211 = _issue1_idx_T_207 < age_considering_issue__53 ? _issue1_idx_T_207 :
    age_considering_issue__53; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_213 = _issue1_idx_T_211 < age_considering_issue__54 ? _issue1_idx_T_209 : 6'h36; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_215 = _issue1_idx_T_211 < age_considering_issue__54 ? _issue1_idx_T_211 :
    age_considering_issue__54; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_217 = _issue1_idx_T_215 < age_considering_issue__55 ? _issue1_idx_T_213 : 6'h37; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_219 = _issue1_idx_T_215 < age_considering_issue__55 ? _issue1_idx_T_215 :
    age_considering_issue__55; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_221 = _issue1_idx_T_219 < age_considering_issue__56 ? _issue1_idx_T_217 : 6'h38; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_223 = _issue1_idx_T_219 < age_considering_issue__56 ? _issue1_idx_T_219 :
    age_considering_issue__56; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_225 = _issue1_idx_T_223 < age_considering_issue__57 ? _issue1_idx_T_221 : 6'h39; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_227 = _issue1_idx_T_223 < age_considering_issue__57 ? _issue1_idx_T_223 :
    age_considering_issue__57; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_229 = _issue1_idx_T_227 < age_considering_issue__58 ? _issue1_idx_T_225 : 6'h3a; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_231 = _issue1_idx_T_227 < age_considering_issue__58 ? _issue1_idx_T_227 :
    age_considering_issue__58; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_233 = _issue1_idx_T_231 < age_considering_issue__59 ? _issue1_idx_T_229 : 6'h3b; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_235 = _issue1_idx_T_231 < age_considering_issue__59 ? _issue1_idx_T_231 :
    age_considering_issue__59; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_237 = _issue1_idx_T_235 < age_considering_issue__60 ? _issue1_idx_T_233 : 6'h3c; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_239 = _issue1_idx_T_235 < age_considering_issue__60 ? _issue1_idx_T_235 :
    age_considering_issue__60; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_241 = _issue1_idx_T_239 < age_considering_issue__61 ? _issue1_idx_T_237 : 6'h3d; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_243 = _issue1_idx_T_239 < age_considering_issue__61 ? _issue1_idx_T_239 :
    age_considering_issue__61; // @[reservation_station.scala 127:82]
  wire [5:0] _issue1_idx_T_245 = _issue1_idx_T_243 < age_considering_issue__62 ? _issue1_idx_T_241 : 6'h3e; // @[reservation_station.scala 127:57]
  wire [7:0] _issue1_idx_T_247 = _issue1_idx_T_243 < age_considering_issue__62 ? _issue1_idx_T_243 :
    age_considering_issue__62; // @[reservation_station.scala 127:82]
  wire [5:0] issue1_idx = _issue1_idx_T_247 < age_considering_issue__63 ? _issue1_idx_T_245 : 6'h3f; // @[reservation_station.scala 127:57]
  wire  _issue1_func_code_T = 6'h0 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_1 = 6'h1 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_2 = 6'h2 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_3 = 6'h3 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_4 = 6'h4 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_5 = 6'h5 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_6 = 6'h6 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_7 = 6'h7 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_8 = 6'h8 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_9 = 6'h9 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_10 = 6'ha == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_11 = 6'hb == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_12 = 6'hc == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_13 = 6'hd == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_14 = 6'he == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_15 = 6'hf == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_16 = 6'h10 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_17 = 6'h11 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_18 = 6'h12 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_19 = 6'h13 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_20 = 6'h14 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_21 = 6'h15 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_22 = 6'h16 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_23 = 6'h17 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_24 = 6'h18 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_25 = 6'h19 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_26 = 6'h1a == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_27 = 6'h1b == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_28 = 6'h1c == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_29 = 6'h1d == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_30 = 6'h1e == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_31 = 6'h1f == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_32 = 6'h20 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_33 = 6'h21 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_34 = 6'h22 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_35 = 6'h23 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_36 = 6'h24 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_37 = 6'h25 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_38 = 6'h26 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_39 = 6'h27 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_40 = 6'h28 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_41 = 6'h29 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_42 = 6'h2a == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_43 = 6'h2b == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_44 = 6'h2c == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_45 = 6'h2d == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_46 = 6'h2e == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_47 = 6'h2f == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_48 = 6'h30 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_49 = 6'h31 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_50 = 6'h32 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_51 = 6'h33 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_52 = 6'h34 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_53 = 6'h35 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_54 = 6'h36 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_55 = 6'h37 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_56 = 6'h38 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_57 = 6'h39 == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_58 = 6'h3a == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_59 = 6'h3b == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_60 = 6'h3c == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_61 = 6'h3d == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_62 = 6'h3e == issue1_idx; // @[reservation_station.scala 130:80]
  wire  _issue1_func_code_T_63 = 6'h3f == issue1_idx; // @[reservation_station.scala 130:80]
  wire [6:0] _issue1_func_code_T_64 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_func_code : 7'h40; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_65 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_func_code :
    _issue1_func_code_T_64; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_66 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_func_code :
    _issue1_func_code_T_65; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_67 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_func_code :
    _issue1_func_code_T_66; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_68 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_func_code :
    _issue1_func_code_T_67; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_69 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_func_code :
    _issue1_func_code_T_68; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_70 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_func_code :
    _issue1_func_code_T_69; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_71 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_func_code :
    _issue1_func_code_T_70; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_72 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_func_code :
    _issue1_func_code_T_71; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_73 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_func_code :
    _issue1_func_code_T_72; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_74 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_func_code :
    _issue1_func_code_T_73; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_75 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_func_code :
    _issue1_func_code_T_74; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_76 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_func_code :
    _issue1_func_code_T_75; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_77 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_func_code :
    _issue1_func_code_T_76; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_78 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_func_code :
    _issue1_func_code_T_77; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_79 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_func_code :
    _issue1_func_code_T_78; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_80 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_func_code :
    _issue1_func_code_T_79; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_81 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_func_code :
    _issue1_func_code_T_80; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_82 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_func_code :
    _issue1_func_code_T_81; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_83 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_func_code :
    _issue1_func_code_T_82; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_84 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_func_code :
    _issue1_func_code_T_83; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_85 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_func_code :
    _issue1_func_code_T_84; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_86 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_func_code :
    _issue1_func_code_T_85; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_87 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_func_code :
    _issue1_func_code_T_86; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_88 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_func_code :
    _issue1_func_code_T_87; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_89 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_func_code :
    _issue1_func_code_T_88; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_90 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_func_code :
    _issue1_func_code_T_89; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_91 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_func_code :
    _issue1_func_code_T_90; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_92 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_func_code :
    _issue1_func_code_T_91; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_93 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_func_code :
    _issue1_func_code_T_92; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_94 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_func_code :
    _issue1_func_code_T_93; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_95 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_func_code :
    _issue1_func_code_T_94; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_96 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_func_code :
    _issue1_func_code_T_95; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_97 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_func_code :
    _issue1_func_code_T_96; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_98 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_func_code :
    _issue1_func_code_T_97; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_99 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_func_code :
    _issue1_func_code_T_98; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_100 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_func_code :
    _issue1_func_code_T_99; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_101 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_func_code :
    _issue1_func_code_T_100; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_102 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_func_code :
    _issue1_func_code_T_101; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_103 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_func_code :
    _issue1_func_code_T_102; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_104 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_func_code :
    _issue1_func_code_T_103; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_105 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_func_code :
    _issue1_func_code_T_104; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_106 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_func_code :
    _issue1_func_code_T_105; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_107 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_func_code :
    _issue1_func_code_T_106; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_108 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_func_code :
    _issue1_func_code_T_107; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_109 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_func_code :
    _issue1_func_code_T_108; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_110 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_func_code :
    _issue1_func_code_T_109; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_111 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_func_code :
    _issue1_func_code_T_110; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_112 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_func_code :
    _issue1_func_code_T_111; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_113 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_func_code :
    _issue1_func_code_T_112; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_114 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_func_code :
    _issue1_func_code_T_113; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_115 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_func_code :
    _issue1_func_code_T_114; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_116 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_func_code :
    _issue1_func_code_T_115; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_117 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_func_code :
    _issue1_func_code_T_116; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_118 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_func_code :
    _issue1_func_code_T_117; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_119 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_func_code :
    _issue1_func_code_T_118; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_120 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_func_code :
    _issue1_func_code_T_119; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_121 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_func_code :
    _issue1_func_code_T_120; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_122 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_func_code :
    _issue1_func_code_T_121; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_123 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_func_code :
    _issue1_func_code_T_122; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_124 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_func_code :
    _issue1_func_code_T_123; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_125 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_func_code :
    _issue1_func_code_T_124; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_126 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_func_code :
    _issue1_func_code_T_125; // @[Mux.scala 101:16]
  wire [6:0] issue1_func_code = _issue1_func_code_T ? reservation_station_0_io_o_uop_func_code : _issue1_func_code_T_126
    ; // @[Mux.scala 101:16]
  wire [2:0] hi = issue1_func_code[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] lo = issue1_func_code[3:0]; // @[OneHot.scala 31:18]
  wire  _T = |hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_19 = {{1'd0}, hi}; // @[OneHot.scala 32:28]
  wire [3:0] _T_1 = _GEN_19 | lo; // @[OneHot.scala 32:28]
  wire [1:0] hi_1 = _T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_1 = _T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _T_2 = |hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _T_3 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  wire [2:0] _T_6 = {_T,_T_2,_T_3[1]}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_1 = 3'h1 == _T_6 ? io_i_available_funcs_1 : io_i_available_funcs_0; // @[reservation_station.scala 151:{109,109}]
  wire [1:0] _GEN_2 = 3'h2 == _T_6 ? io_i_available_funcs_2 : _GEN_1; // @[reservation_station.scala 151:{109,109}]
  wire [1:0] _GEN_3 = 3'h3 == _T_6 ? io_i_available_funcs_3 : _GEN_2; // @[reservation_station.scala 151:{109,109}]
  wire [1:0] _GEN_4 = 3'h4 == _T_6 ? io_i_available_funcs_4 : _GEN_3; // @[reservation_station.scala 151:{109,109}]
  wire [1:0] _GEN_5 = 3'h5 == _T_6 ? io_i_available_funcs_5 : _GEN_4; // @[reservation_station.scala 151:{109,109}]
  wire [1:0] _GEN_6 = 3'h6 == _T_6 ? 2'h0 : _GEN_5; // @[reservation_station.scala 151:{109,109}]
  wire [1:0] _available_funcs_with_mask_T_8 = _GEN_6 - 2'h1; // @[reservation_station.scala 151:109]
  wire [1:0] available_funcs_with_mask_0 = 3'h0 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_0; // @[reservation_station.scala 133:31 151:{59,59}]
  wire [1:0] available_funcs_with_mask_1 = 3'h1 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_1; // @[reservation_station.scala 133:31 151:{59,59}]
  wire [1:0] available_funcs_with_mask_2 = 3'h2 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_2; // @[reservation_station.scala 133:31 151:{59,59}]
  wire [1:0] available_funcs_with_mask_3 = 3'h3 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_3; // @[reservation_station.scala 133:31 151:{59,59}]
  wire [1:0] available_funcs_with_mask_4 = 3'h4 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_4; // @[reservation_station.scala 133:31 151:{59,59}]
  wire [1:0] available_funcs_with_mask_5 = 3'h5 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_5; // @[reservation_station.scala 133:31 151:{59,59}]
  wire [1:0] available_funcs_with_mask_6 = 3'h6 == _T_6 ? _available_funcs_with_mask_T_8 : 2'h0; // @[reservation_station.scala 133:31 151:{59,59}]
  wire  temp3_0 = |available_funcs_with_mask_0; // @[reservation_station.scala 155:49]
  wire  temp3_1 = |available_funcs_with_mask_1; // @[reservation_station.scala 155:49]
  wire  temp3_2 = |available_funcs_with_mask_2; // @[reservation_station.scala 155:49]
  wire  temp3_3 = |available_funcs_with_mask_3; // @[reservation_station.scala 155:49]
  wire  temp3_4 = |available_funcs_with_mask_4; // @[reservation_station.scala 155:49]
  wire  temp3_5 = |available_funcs_with_mask_5; // @[reservation_station.scala 155:49]
  wire  temp3_6 = |available_funcs_with_mask_6; // @[reservation_station.scala 155:49]
  wire [6:0] available_funcs2_bits = {temp3_6,temp3_5,temp3_4,temp3_3,temp3_2,temp3_1,temp3_0}; // @[reservation_station.scala 157:46]
  wire [7:0] _age_considering_issue_2_T_2 = _issue1_func_code_T ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_3 = age_considering_issue__0 | _age_considering_issue_2_T_2; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_4 = reservation_station_0_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_5 = |_age_considering_issue_2_T_4; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_7 = _age_considering_issue_2_T_5 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_8 = ~_age_considering_issue_2_T_7; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_0 = _age_considering_issue_2_T_3 | _age_considering_issue_2_T_8; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_12 = _issue1_func_code_T_1 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_13 = age_considering_issue__1 | _age_considering_issue_2_T_12; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_14 = reservation_station_1_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_15 = |_age_considering_issue_2_T_14; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_17 = _age_considering_issue_2_T_15 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_18 = ~_age_considering_issue_2_T_17; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_1 = _age_considering_issue_2_T_13 | _age_considering_issue_2_T_18; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_22 = _issue1_func_code_T_2 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_23 = age_considering_issue__2 | _age_considering_issue_2_T_22; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_24 = reservation_station_2_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_25 = |_age_considering_issue_2_T_24; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_27 = _age_considering_issue_2_T_25 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_28 = ~_age_considering_issue_2_T_27; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_2 = _age_considering_issue_2_T_23 | _age_considering_issue_2_T_28; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_32 = _issue1_func_code_T_3 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_33 = age_considering_issue__3 | _age_considering_issue_2_T_32; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_34 = reservation_station_3_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_35 = |_age_considering_issue_2_T_34; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_37 = _age_considering_issue_2_T_35 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_38 = ~_age_considering_issue_2_T_37; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_3 = _age_considering_issue_2_T_33 | _age_considering_issue_2_T_38; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_42 = _issue1_func_code_T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_43 = age_considering_issue__4 | _age_considering_issue_2_T_42; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_44 = reservation_station_4_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_45 = |_age_considering_issue_2_T_44; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_47 = _age_considering_issue_2_T_45 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_48 = ~_age_considering_issue_2_T_47; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_4 = _age_considering_issue_2_T_43 | _age_considering_issue_2_T_48; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_52 = _issue1_func_code_T_5 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_53 = age_considering_issue__5 | _age_considering_issue_2_T_52; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_54 = reservation_station_5_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_55 = |_age_considering_issue_2_T_54; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_57 = _age_considering_issue_2_T_55 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_58 = ~_age_considering_issue_2_T_57; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_5 = _age_considering_issue_2_T_53 | _age_considering_issue_2_T_58; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_62 = _issue1_func_code_T_6 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_63 = age_considering_issue__6 | _age_considering_issue_2_T_62; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_64 = reservation_station_6_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_65 = |_age_considering_issue_2_T_64; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_67 = _age_considering_issue_2_T_65 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_68 = ~_age_considering_issue_2_T_67; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_6 = _age_considering_issue_2_T_63 | _age_considering_issue_2_T_68; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_72 = _issue1_func_code_T_7 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_73 = age_considering_issue__7 | _age_considering_issue_2_T_72; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_74 = reservation_station_7_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_75 = |_age_considering_issue_2_T_74; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_77 = _age_considering_issue_2_T_75 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_78 = ~_age_considering_issue_2_T_77; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_7 = _age_considering_issue_2_T_73 | _age_considering_issue_2_T_78; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_82 = _issue1_func_code_T_8 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_83 = age_considering_issue__8 | _age_considering_issue_2_T_82; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_84 = reservation_station_8_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_85 = |_age_considering_issue_2_T_84; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_87 = _age_considering_issue_2_T_85 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_88 = ~_age_considering_issue_2_T_87; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_8 = _age_considering_issue_2_T_83 | _age_considering_issue_2_T_88; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_92 = _issue1_func_code_T_9 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_93 = age_considering_issue__9 | _age_considering_issue_2_T_92; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_94 = reservation_station_9_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_95 = |_age_considering_issue_2_T_94; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_97 = _age_considering_issue_2_T_95 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_98 = ~_age_considering_issue_2_T_97; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_9 = _age_considering_issue_2_T_93 | _age_considering_issue_2_T_98; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_102 = _issue1_func_code_T_10 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_103 = age_considering_issue__10 | _age_considering_issue_2_T_102; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_104 = reservation_station_10_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_105 = |_age_considering_issue_2_T_104; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_107 = _age_considering_issue_2_T_105 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_108 = ~_age_considering_issue_2_T_107; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_10 = _age_considering_issue_2_T_103 | _age_considering_issue_2_T_108; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_112 = _issue1_func_code_T_11 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_113 = age_considering_issue__11 | _age_considering_issue_2_T_112; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_114 = reservation_station_11_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_115 = |_age_considering_issue_2_T_114; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_117 = _age_considering_issue_2_T_115 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_118 = ~_age_considering_issue_2_T_117; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_11 = _age_considering_issue_2_T_113 | _age_considering_issue_2_T_118; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_122 = _issue1_func_code_T_12 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_123 = age_considering_issue__12 | _age_considering_issue_2_T_122; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_124 = reservation_station_12_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_125 = |_age_considering_issue_2_T_124; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_127 = _age_considering_issue_2_T_125 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_128 = ~_age_considering_issue_2_T_127; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_12 = _age_considering_issue_2_T_123 | _age_considering_issue_2_T_128; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_132 = _issue1_func_code_T_13 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_133 = age_considering_issue__13 | _age_considering_issue_2_T_132; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_134 = reservation_station_13_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_135 = |_age_considering_issue_2_T_134; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_137 = _age_considering_issue_2_T_135 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_138 = ~_age_considering_issue_2_T_137; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_13 = _age_considering_issue_2_T_133 | _age_considering_issue_2_T_138; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_142 = _issue1_func_code_T_14 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_143 = age_considering_issue__14 | _age_considering_issue_2_T_142; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_144 = reservation_station_14_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_145 = |_age_considering_issue_2_T_144; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_147 = _age_considering_issue_2_T_145 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_148 = ~_age_considering_issue_2_T_147; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_14 = _age_considering_issue_2_T_143 | _age_considering_issue_2_T_148; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_152 = _issue1_func_code_T_15 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_153 = age_considering_issue__15 | _age_considering_issue_2_T_152; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_154 = reservation_station_15_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_155 = |_age_considering_issue_2_T_154; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_157 = _age_considering_issue_2_T_155 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_158 = ~_age_considering_issue_2_T_157; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_15 = _age_considering_issue_2_T_153 | _age_considering_issue_2_T_158; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_162 = _issue1_func_code_T_16 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_163 = age_considering_issue__16 | _age_considering_issue_2_T_162; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_164 = reservation_station_16_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_165 = |_age_considering_issue_2_T_164; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_167 = _age_considering_issue_2_T_165 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_168 = ~_age_considering_issue_2_T_167; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_16 = _age_considering_issue_2_T_163 | _age_considering_issue_2_T_168; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_172 = _issue1_func_code_T_17 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_173 = age_considering_issue__17 | _age_considering_issue_2_T_172; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_174 = reservation_station_17_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_175 = |_age_considering_issue_2_T_174; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_177 = _age_considering_issue_2_T_175 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_178 = ~_age_considering_issue_2_T_177; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_17 = _age_considering_issue_2_T_173 | _age_considering_issue_2_T_178; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_182 = _issue1_func_code_T_18 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_183 = age_considering_issue__18 | _age_considering_issue_2_T_182; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_184 = reservation_station_18_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_185 = |_age_considering_issue_2_T_184; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_187 = _age_considering_issue_2_T_185 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_188 = ~_age_considering_issue_2_T_187; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_18 = _age_considering_issue_2_T_183 | _age_considering_issue_2_T_188; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_192 = _issue1_func_code_T_19 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_193 = age_considering_issue__19 | _age_considering_issue_2_T_192; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_194 = reservation_station_19_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_195 = |_age_considering_issue_2_T_194; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_197 = _age_considering_issue_2_T_195 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_198 = ~_age_considering_issue_2_T_197; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_19 = _age_considering_issue_2_T_193 | _age_considering_issue_2_T_198; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_202 = _issue1_func_code_T_20 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_203 = age_considering_issue__20 | _age_considering_issue_2_T_202; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_204 = reservation_station_20_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_205 = |_age_considering_issue_2_T_204; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_207 = _age_considering_issue_2_T_205 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_208 = ~_age_considering_issue_2_T_207; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_20 = _age_considering_issue_2_T_203 | _age_considering_issue_2_T_208; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_212 = _issue1_func_code_T_21 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_213 = age_considering_issue__21 | _age_considering_issue_2_T_212; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_214 = reservation_station_21_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_215 = |_age_considering_issue_2_T_214; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_217 = _age_considering_issue_2_T_215 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_218 = ~_age_considering_issue_2_T_217; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_21 = _age_considering_issue_2_T_213 | _age_considering_issue_2_T_218; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_222 = _issue1_func_code_T_22 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_223 = age_considering_issue__22 | _age_considering_issue_2_T_222; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_224 = reservation_station_22_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_225 = |_age_considering_issue_2_T_224; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_227 = _age_considering_issue_2_T_225 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_228 = ~_age_considering_issue_2_T_227; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_22 = _age_considering_issue_2_T_223 | _age_considering_issue_2_T_228; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_232 = _issue1_func_code_T_23 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_233 = age_considering_issue__23 | _age_considering_issue_2_T_232; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_234 = reservation_station_23_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_235 = |_age_considering_issue_2_T_234; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_237 = _age_considering_issue_2_T_235 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_238 = ~_age_considering_issue_2_T_237; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_23 = _age_considering_issue_2_T_233 | _age_considering_issue_2_T_238; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_242 = _issue1_func_code_T_24 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_243 = age_considering_issue__24 | _age_considering_issue_2_T_242; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_244 = reservation_station_24_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_245 = |_age_considering_issue_2_T_244; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_247 = _age_considering_issue_2_T_245 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_248 = ~_age_considering_issue_2_T_247; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_24 = _age_considering_issue_2_T_243 | _age_considering_issue_2_T_248; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_252 = _issue1_func_code_T_25 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_253 = age_considering_issue__25 | _age_considering_issue_2_T_252; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_254 = reservation_station_25_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_255 = |_age_considering_issue_2_T_254; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_257 = _age_considering_issue_2_T_255 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_258 = ~_age_considering_issue_2_T_257; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_25 = _age_considering_issue_2_T_253 | _age_considering_issue_2_T_258; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_262 = _issue1_func_code_T_26 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_263 = age_considering_issue__26 | _age_considering_issue_2_T_262; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_264 = reservation_station_26_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_265 = |_age_considering_issue_2_T_264; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_267 = _age_considering_issue_2_T_265 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_268 = ~_age_considering_issue_2_T_267; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_26 = _age_considering_issue_2_T_263 | _age_considering_issue_2_T_268; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_272 = _issue1_func_code_T_27 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_273 = age_considering_issue__27 | _age_considering_issue_2_T_272; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_274 = reservation_station_27_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_275 = |_age_considering_issue_2_T_274; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_277 = _age_considering_issue_2_T_275 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_278 = ~_age_considering_issue_2_T_277; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_27 = _age_considering_issue_2_T_273 | _age_considering_issue_2_T_278; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_282 = _issue1_func_code_T_28 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_283 = age_considering_issue__28 | _age_considering_issue_2_T_282; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_284 = reservation_station_28_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_285 = |_age_considering_issue_2_T_284; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_287 = _age_considering_issue_2_T_285 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_288 = ~_age_considering_issue_2_T_287; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_28 = _age_considering_issue_2_T_283 | _age_considering_issue_2_T_288; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_292 = _issue1_func_code_T_29 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_293 = age_considering_issue__29 | _age_considering_issue_2_T_292; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_294 = reservation_station_29_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_295 = |_age_considering_issue_2_T_294; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_297 = _age_considering_issue_2_T_295 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_298 = ~_age_considering_issue_2_T_297; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_29 = _age_considering_issue_2_T_293 | _age_considering_issue_2_T_298; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_302 = _issue1_func_code_T_30 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_303 = age_considering_issue__30 | _age_considering_issue_2_T_302; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_304 = reservation_station_30_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_305 = |_age_considering_issue_2_T_304; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_307 = _age_considering_issue_2_T_305 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_308 = ~_age_considering_issue_2_T_307; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_30 = _age_considering_issue_2_T_303 | _age_considering_issue_2_T_308; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_312 = _issue1_func_code_T_31 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_313 = age_considering_issue__31 | _age_considering_issue_2_T_312; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_314 = reservation_station_31_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_315 = |_age_considering_issue_2_T_314; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_317 = _age_considering_issue_2_T_315 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_318 = ~_age_considering_issue_2_T_317; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_31 = _age_considering_issue_2_T_313 | _age_considering_issue_2_T_318; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_322 = _issue1_func_code_T_32 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_323 = age_considering_issue__32 | _age_considering_issue_2_T_322; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_324 = reservation_station_32_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_325 = |_age_considering_issue_2_T_324; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_327 = _age_considering_issue_2_T_325 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_328 = ~_age_considering_issue_2_T_327; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_32 = _age_considering_issue_2_T_323 | _age_considering_issue_2_T_328; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_332 = _issue1_func_code_T_33 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_333 = age_considering_issue__33 | _age_considering_issue_2_T_332; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_334 = reservation_station_33_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_335 = |_age_considering_issue_2_T_334; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_337 = _age_considering_issue_2_T_335 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_338 = ~_age_considering_issue_2_T_337; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_33 = _age_considering_issue_2_T_333 | _age_considering_issue_2_T_338; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_342 = _issue1_func_code_T_34 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_343 = age_considering_issue__34 | _age_considering_issue_2_T_342; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_344 = reservation_station_34_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_345 = |_age_considering_issue_2_T_344; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_347 = _age_considering_issue_2_T_345 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_348 = ~_age_considering_issue_2_T_347; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_34 = _age_considering_issue_2_T_343 | _age_considering_issue_2_T_348; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_352 = _issue1_func_code_T_35 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_353 = age_considering_issue__35 | _age_considering_issue_2_T_352; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_354 = reservation_station_35_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_355 = |_age_considering_issue_2_T_354; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_357 = _age_considering_issue_2_T_355 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_358 = ~_age_considering_issue_2_T_357; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_35 = _age_considering_issue_2_T_353 | _age_considering_issue_2_T_358; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_362 = _issue1_func_code_T_36 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_363 = age_considering_issue__36 | _age_considering_issue_2_T_362; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_364 = reservation_station_36_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_365 = |_age_considering_issue_2_T_364; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_367 = _age_considering_issue_2_T_365 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_368 = ~_age_considering_issue_2_T_367; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_36 = _age_considering_issue_2_T_363 | _age_considering_issue_2_T_368; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_372 = _issue1_func_code_T_37 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_373 = age_considering_issue__37 | _age_considering_issue_2_T_372; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_374 = reservation_station_37_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_375 = |_age_considering_issue_2_T_374; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_377 = _age_considering_issue_2_T_375 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_378 = ~_age_considering_issue_2_T_377; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_37 = _age_considering_issue_2_T_373 | _age_considering_issue_2_T_378; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_382 = _issue1_func_code_T_38 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_383 = age_considering_issue__38 | _age_considering_issue_2_T_382; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_384 = reservation_station_38_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_385 = |_age_considering_issue_2_T_384; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_387 = _age_considering_issue_2_T_385 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_388 = ~_age_considering_issue_2_T_387; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_38 = _age_considering_issue_2_T_383 | _age_considering_issue_2_T_388; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_392 = _issue1_func_code_T_39 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_393 = age_considering_issue__39 | _age_considering_issue_2_T_392; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_394 = reservation_station_39_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_395 = |_age_considering_issue_2_T_394; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_397 = _age_considering_issue_2_T_395 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_398 = ~_age_considering_issue_2_T_397; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_39 = _age_considering_issue_2_T_393 | _age_considering_issue_2_T_398; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_402 = _issue1_func_code_T_40 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_403 = age_considering_issue__40 | _age_considering_issue_2_T_402; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_404 = reservation_station_40_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_405 = |_age_considering_issue_2_T_404; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_407 = _age_considering_issue_2_T_405 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_408 = ~_age_considering_issue_2_T_407; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_40 = _age_considering_issue_2_T_403 | _age_considering_issue_2_T_408; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_412 = _issue1_func_code_T_41 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_413 = age_considering_issue__41 | _age_considering_issue_2_T_412; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_414 = reservation_station_41_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_415 = |_age_considering_issue_2_T_414; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_417 = _age_considering_issue_2_T_415 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_418 = ~_age_considering_issue_2_T_417; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_41 = _age_considering_issue_2_T_413 | _age_considering_issue_2_T_418; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_422 = _issue1_func_code_T_42 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_423 = age_considering_issue__42 | _age_considering_issue_2_T_422; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_424 = reservation_station_42_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_425 = |_age_considering_issue_2_T_424; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_427 = _age_considering_issue_2_T_425 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_428 = ~_age_considering_issue_2_T_427; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_42 = _age_considering_issue_2_T_423 | _age_considering_issue_2_T_428; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_432 = _issue1_func_code_T_43 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_433 = age_considering_issue__43 | _age_considering_issue_2_T_432; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_434 = reservation_station_43_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_435 = |_age_considering_issue_2_T_434; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_437 = _age_considering_issue_2_T_435 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_438 = ~_age_considering_issue_2_T_437; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_43 = _age_considering_issue_2_T_433 | _age_considering_issue_2_T_438; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_442 = _issue1_func_code_T_44 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_443 = age_considering_issue__44 | _age_considering_issue_2_T_442; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_444 = reservation_station_44_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_445 = |_age_considering_issue_2_T_444; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_447 = _age_considering_issue_2_T_445 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_448 = ~_age_considering_issue_2_T_447; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_44 = _age_considering_issue_2_T_443 | _age_considering_issue_2_T_448; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_452 = _issue1_func_code_T_45 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_453 = age_considering_issue__45 | _age_considering_issue_2_T_452; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_454 = reservation_station_45_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_455 = |_age_considering_issue_2_T_454; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_457 = _age_considering_issue_2_T_455 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_458 = ~_age_considering_issue_2_T_457; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_45 = _age_considering_issue_2_T_453 | _age_considering_issue_2_T_458; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_462 = _issue1_func_code_T_46 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_463 = age_considering_issue__46 | _age_considering_issue_2_T_462; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_464 = reservation_station_46_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_465 = |_age_considering_issue_2_T_464; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_467 = _age_considering_issue_2_T_465 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_468 = ~_age_considering_issue_2_T_467; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_46 = _age_considering_issue_2_T_463 | _age_considering_issue_2_T_468; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_472 = _issue1_func_code_T_47 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_473 = age_considering_issue__47 | _age_considering_issue_2_T_472; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_474 = reservation_station_47_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_475 = |_age_considering_issue_2_T_474; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_477 = _age_considering_issue_2_T_475 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_478 = ~_age_considering_issue_2_T_477; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_47 = _age_considering_issue_2_T_473 | _age_considering_issue_2_T_478; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_482 = _issue1_func_code_T_48 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_483 = age_considering_issue__48 | _age_considering_issue_2_T_482; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_484 = reservation_station_48_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_485 = |_age_considering_issue_2_T_484; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_487 = _age_considering_issue_2_T_485 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_488 = ~_age_considering_issue_2_T_487; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_48 = _age_considering_issue_2_T_483 | _age_considering_issue_2_T_488; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_492 = _issue1_func_code_T_49 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_493 = age_considering_issue__49 | _age_considering_issue_2_T_492; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_494 = reservation_station_49_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_495 = |_age_considering_issue_2_T_494; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_497 = _age_considering_issue_2_T_495 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_498 = ~_age_considering_issue_2_T_497; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_49 = _age_considering_issue_2_T_493 | _age_considering_issue_2_T_498; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_502 = _issue1_func_code_T_50 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_503 = age_considering_issue__50 | _age_considering_issue_2_T_502; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_504 = reservation_station_50_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_505 = |_age_considering_issue_2_T_504; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_507 = _age_considering_issue_2_T_505 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_508 = ~_age_considering_issue_2_T_507; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_50 = _age_considering_issue_2_T_503 | _age_considering_issue_2_T_508; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_512 = _issue1_func_code_T_51 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_513 = age_considering_issue__51 | _age_considering_issue_2_T_512; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_514 = reservation_station_51_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_515 = |_age_considering_issue_2_T_514; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_517 = _age_considering_issue_2_T_515 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_518 = ~_age_considering_issue_2_T_517; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_51 = _age_considering_issue_2_T_513 | _age_considering_issue_2_T_518; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_522 = _issue1_func_code_T_52 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_523 = age_considering_issue__52 | _age_considering_issue_2_T_522; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_524 = reservation_station_52_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_525 = |_age_considering_issue_2_T_524; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_527 = _age_considering_issue_2_T_525 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_528 = ~_age_considering_issue_2_T_527; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_52 = _age_considering_issue_2_T_523 | _age_considering_issue_2_T_528; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_532 = _issue1_func_code_T_53 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_533 = age_considering_issue__53 | _age_considering_issue_2_T_532; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_534 = reservation_station_53_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_535 = |_age_considering_issue_2_T_534; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_537 = _age_considering_issue_2_T_535 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_538 = ~_age_considering_issue_2_T_537; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_53 = _age_considering_issue_2_T_533 | _age_considering_issue_2_T_538; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_542 = _issue1_func_code_T_54 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_543 = age_considering_issue__54 | _age_considering_issue_2_T_542; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_544 = reservation_station_54_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_545 = |_age_considering_issue_2_T_544; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_547 = _age_considering_issue_2_T_545 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_548 = ~_age_considering_issue_2_T_547; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_54 = _age_considering_issue_2_T_543 | _age_considering_issue_2_T_548; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_552 = _issue1_func_code_T_55 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_553 = age_considering_issue__55 | _age_considering_issue_2_T_552; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_554 = reservation_station_55_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_555 = |_age_considering_issue_2_T_554; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_557 = _age_considering_issue_2_T_555 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_558 = ~_age_considering_issue_2_T_557; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_55 = _age_considering_issue_2_T_553 | _age_considering_issue_2_T_558; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_562 = _issue1_func_code_T_56 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_563 = age_considering_issue__56 | _age_considering_issue_2_T_562; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_564 = reservation_station_56_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_565 = |_age_considering_issue_2_T_564; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_567 = _age_considering_issue_2_T_565 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_568 = ~_age_considering_issue_2_T_567; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_56 = _age_considering_issue_2_T_563 | _age_considering_issue_2_T_568; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_572 = _issue1_func_code_T_57 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_573 = age_considering_issue__57 | _age_considering_issue_2_T_572; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_574 = reservation_station_57_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_575 = |_age_considering_issue_2_T_574; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_577 = _age_considering_issue_2_T_575 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_578 = ~_age_considering_issue_2_T_577; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_57 = _age_considering_issue_2_T_573 | _age_considering_issue_2_T_578; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_582 = _issue1_func_code_T_58 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_583 = age_considering_issue__58 | _age_considering_issue_2_T_582; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_584 = reservation_station_58_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_585 = |_age_considering_issue_2_T_584; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_587 = _age_considering_issue_2_T_585 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_588 = ~_age_considering_issue_2_T_587; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_58 = _age_considering_issue_2_T_583 | _age_considering_issue_2_T_588; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_592 = _issue1_func_code_T_59 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_593 = age_considering_issue__59 | _age_considering_issue_2_T_592; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_594 = reservation_station_59_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_595 = |_age_considering_issue_2_T_594; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_597 = _age_considering_issue_2_T_595 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_598 = ~_age_considering_issue_2_T_597; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_59 = _age_considering_issue_2_T_593 | _age_considering_issue_2_T_598; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_602 = _issue1_func_code_T_60 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_603 = age_considering_issue__60 | _age_considering_issue_2_T_602; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_604 = reservation_station_60_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_605 = |_age_considering_issue_2_T_604; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_607 = _age_considering_issue_2_T_605 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_608 = ~_age_considering_issue_2_T_607; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_60 = _age_considering_issue_2_T_603 | _age_considering_issue_2_T_608; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_612 = _issue1_func_code_T_61 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_613 = age_considering_issue__61 | _age_considering_issue_2_T_612; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_614 = reservation_station_61_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_615 = |_age_considering_issue_2_T_614; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_617 = _age_considering_issue_2_T_615 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_618 = ~_age_considering_issue_2_T_617; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_61 = _age_considering_issue_2_T_613 | _age_considering_issue_2_T_618; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_622 = _issue1_func_code_T_62 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_623 = age_considering_issue__62 | _age_considering_issue_2_T_622; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_624 = reservation_station_62_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_625 = |_age_considering_issue_2_T_624; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_627 = _age_considering_issue_2_T_625 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_628 = ~_age_considering_issue_2_T_627; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_62 = _age_considering_issue_2_T_623 | _age_considering_issue_2_T_628; // @[reservation_station.scala 159:8]
  wire [7:0] _age_considering_issue_2_T_632 = _issue1_func_code_T_63 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_633 = age_considering_issue__63 | _age_considering_issue_2_T_632; // @[reservation_station.scala 158:86]
  wire [6:0] _age_considering_issue_2_T_634 = reservation_station_63_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 159:61]
  wire  _age_considering_issue_2_T_635 = |_age_considering_issue_2_T_634; // @[reservation_station.scala 159:86]
  wire [7:0] _age_considering_issue_2_T_637 = _age_considering_issue_2_T_635 ? 8'hff : 8'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _age_considering_issue_2_T_638 = ~_age_considering_issue_2_T_637; // @[reservation_station.scala 159:10]
  wire [7:0] age_considering_issue_2_63 = _age_considering_issue_2_T_633 | _age_considering_issue_2_T_638; // @[reservation_station.scala 159:8]
  wire [5:0] _issue2_idx_T_1 = age_considering_issue_2_62 < age_considering_issue_2_63 ? 6'h3e : 6'h3f; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_3 = age_considering_issue_2_62 < age_considering_issue_2_63 ? age_considering_issue_2_62 :
    age_considering_issue_2_63; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_5 = age_considering_issue_2_61 < _issue2_idx_T_3 ? 6'h3d : _issue2_idx_T_1; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_7 = age_considering_issue_2_61 < _issue2_idx_T_3 ? age_considering_issue_2_61 :
    _issue2_idx_T_3; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_9 = age_considering_issue_2_60 < _issue2_idx_T_7 ? 6'h3c : _issue2_idx_T_5; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_11 = age_considering_issue_2_60 < _issue2_idx_T_7 ? age_considering_issue_2_60 :
    _issue2_idx_T_7; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_13 = age_considering_issue_2_59 < _issue2_idx_T_11 ? 6'h3b : _issue2_idx_T_9; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_15 = age_considering_issue_2_59 < _issue2_idx_T_11 ? age_considering_issue_2_59 :
    _issue2_idx_T_11; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_17 = age_considering_issue_2_58 < _issue2_idx_T_15 ? 6'h3a : _issue2_idx_T_13; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_19 = age_considering_issue_2_58 < _issue2_idx_T_15 ? age_considering_issue_2_58 :
    _issue2_idx_T_15; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_21 = age_considering_issue_2_57 < _issue2_idx_T_19 ? 6'h39 : _issue2_idx_T_17; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_23 = age_considering_issue_2_57 < _issue2_idx_T_19 ? age_considering_issue_2_57 :
    _issue2_idx_T_19; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_25 = age_considering_issue_2_56 < _issue2_idx_T_23 ? 6'h38 : _issue2_idx_T_21; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_27 = age_considering_issue_2_56 < _issue2_idx_T_23 ? age_considering_issue_2_56 :
    _issue2_idx_T_23; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_29 = age_considering_issue_2_55 < _issue2_idx_T_27 ? 6'h37 : _issue2_idx_T_25; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_31 = age_considering_issue_2_55 < _issue2_idx_T_27 ? age_considering_issue_2_55 :
    _issue2_idx_T_27; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_33 = age_considering_issue_2_54 < _issue2_idx_T_31 ? 6'h36 : _issue2_idx_T_29; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_35 = age_considering_issue_2_54 < _issue2_idx_T_31 ? age_considering_issue_2_54 :
    _issue2_idx_T_31; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_37 = age_considering_issue_2_53 < _issue2_idx_T_35 ? 6'h35 : _issue2_idx_T_33; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_39 = age_considering_issue_2_53 < _issue2_idx_T_35 ? age_considering_issue_2_53 :
    _issue2_idx_T_35; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_41 = age_considering_issue_2_52 < _issue2_idx_T_39 ? 6'h34 : _issue2_idx_T_37; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_43 = age_considering_issue_2_52 < _issue2_idx_T_39 ? age_considering_issue_2_52 :
    _issue2_idx_T_39; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_45 = age_considering_issue_2_51 < _issue2_idx_T_43 ? 6'h33 : _issue2_idx_T_41; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_47 = age_considering_issue_2_51 < _issue2_idx_T_43 ? age_considering_issue_2_51 :
    _issue2_idx_T_43; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_49 = age_considering_issue_2_50 < _issue2_idx_T_47 ? 6'h32 : _issue2_idx_T_45; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_51 = age_considering_issue_2_50 < _issue2_idx_T_47 ? age_considering_issue_2_50 :
    _issue2_idx_T_47; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_53 = age_considering_issue_2_49 < _issue2_idx_T_51 ? 6'h31 : _issue2_idx_T_49; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_55 = age_considering_issue_2_49 < _issue2_idx_T_51 ? age_considering_issue_2_49 :
    _issue2_idx_T_51; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_57 = age_considering_issue_2_48 < _issue2_idx_T_55 ? 6'h30 : _issue2_idx_T_53; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_59 = age_considering_issue_2_48 < _issue2_idx_T_55 ? age_considering_issue_2_48 :
    _issue2_idx_T_55; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_61 = age_considering_issue_2_47 < _issue2_idx_T_59 ? 6'h2f : _issue2_idx_T_57; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_63 = age_considering_issue_2_47 < _issue2_idx_T_59 ? age_considering_issue_2_47 :
    _issue2_idx_T_59; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_65 = age_considering_issue_2_46 < _issue2_idx_T_63 ? 6'h2e : _issue2_idx_T_61; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_67 = age_considering_issue_2_46 < _issue2_idx_T_63 ? age_considering_issue_2_46 :
    _issue2_idx_T_63; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_69 = age_considering_issue_2_45 < _issue2_idx_T_67 ? 6'h2d : _issue2_idx_T_65; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_71 = age_considering_issue_2_45 < _issue2_idx_T_67 ? age_considering_issue_2_45 :
    _issue2_idx_T_67; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_73 = age_considering_issue_2_44 < _issue2_idx_T_71 ? 6'h2c : _issue2_idx_T_69; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_75 = age_considering_issue_2_44 < _issue2_idx_T_71 ? age_considering_issue_2_44 :
    _issue2_idx_T_71; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_77 = age_considering_issue_2_43 < _issue2_idx_T_75 ? 6'h2b : _issue2_idx_T_73; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_79 = age_considering_issue_2_43 < _issue2_idx_T_75 ? age_considering_issue_2_43 :
    _issue2_idx_T_75; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_81 = age_considering_issue_2_42 < _issue2_idx_T_79 ? 6'h2a : _issue2_idx_T_77; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_83 = age_considering_issue_2_42 < _issue2_idx_T_79 ? age_considering_issue_2_42 :
    _issue2_idx_T_79; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_85 = age_considering_issue_2_41 < _issue2_idx_T_83 ? 6'h29 : _issue2_idx_T_81; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_87 = age_considering_issue_2_41 < _issue2_idx_T_83 ? age_considering_issue_2_41 :
    _issue2_idx_T_83; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_89 = age_considering_issue_2_40 < _issue2_idx_T_87 ? 6'h28 : _issue2_idx_T_85; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_91 = age_considering_issue_2_40 < _issue2_idx_T_87 ? age_considering_issue_2_40 :
    _issue2_idx_T_87; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_93 = age_considering_issue_2_39 < _issue2_idx_T_91 ? 6'h27 : _issue2_idx_T_89; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_95 = age_considering_issue_2_39 < _issue2_idx_T_91 ? age_considering_issue_2_39 :
    _issue2_idx_T_91; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_97 = age_considering_issue_2_38 < _issue2_idx_T_95 ? 6'h26 : _issue2_idx_T_93; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_99 = age_considering_issue_2_38 < _issue2_idx_T_95 ? age_considering_issue_2_38 :
    _issue2_idx_T_95; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_101 = age_considering_issue_2_37 < _issue2_idx_T_99 ? 6'h25 : _issue2_idx_T_97; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_103 = age_considering_issue_2_37 < _issue2_idx_T_99 ? age_considering_issue_2_37 :
    _issue2_idx_T_99; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_105 = age_considering_issue_2_36 < _issue2_idx_T_103 ? 6'h24 : _issue2_idx_T_101; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_107 = age_considering_issue_2_36 < _issue2_idx_T_103 ? age_considering_issue_2_36 :
    _issue2_idx_T_103; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_109 = age_considering_issue_2_35 < _issue2_idx_T_107 ? 6'h23 : _issue2_idx_T_105; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_111 = age_considering_issue_2_35 < _issue2_idx_T_107 ? age_considering_issue_2_35 :
    _issue2_idx_T_107; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_113 = age_considering_issue_2_34 < _issue2_idx_T_111 ? 6'h22 : _issue2_idx_T_109; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_115 = age_considering_issue_2_34 < _issue2_idx_T_111 ? age_considering_issue_2_34 :
    _issue2_idx_T_111; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_117 = age_considering_issue_2_33 < _issue2_idx_T_115 ? 6'h21 : _issue2_idx_T_113; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_119 = age_considering_issue_2_33 < _issue2_idx_T_115 ? age_considering_issue_2_33 :
    _issue2_idx_T_115; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_121 = age_considering_issue_2_32 < _issue2_idx_T_119 ? 6'h20 : _issue2_idx_T_117; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_123 = age_considering_issue_2_32 < _issue2_idx_T_119 ? age_considering_issue_2_32 :
    _issue2_idx_T_119; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_125 = age_considering_issue_2_31 < _issue2_idx_T_123 ? 6'h1f : _issue2_idx_T_121; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_127 = age_considering_issue_2_31 < _issue2_idx_T_123 ? age_considering_issue_2_31 :
    _issue2_idx_T_123; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_129 = age_considering_issue_2_30 < _issue2_idx_T_127 ? 6'h1e : _issue2_idx_T_125; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_131 = age_considering_issue_2_30 < _issue2_idx_T_127 ? age_considering_issue_2_30 :
    _issue2_idx_T_127; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_133 = age_considering_issue_2_29 < _issue2_idx_T_131 ? 6'h1d : _issue2_idx_T_129; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_135 = age_considering_issue_2_29 < _issue2_idx_T_131 ? age_considering_issue_2_29 :
    _issue2_idx_T_131; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_137 = age_considering_issue_2_28 < _issue2_idx_T_135 ? 6'h1c : _issue2_idx_T_133; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_139 = age_considering_issue_2_28 < _issue2_idx_T_135 ? age_considering_issue_2_28 :
    _issue2_idx_T_135; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_141 = age_considering_issue_2_27 < _issue2_idx_T_139 ? 6'h1b : _issue2_idx_T_137; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_143 = age_considering_issue_2_27 < _issue2_idx_T_139 ? age_considering_issue_2_27 :
    _issue2_idx_T_139; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_145 = age_considering_issue_2_26 < _issue2_idx_T_143 ? 6'h1a : _issue2_idx_T_141; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_147 = age_considering_issue_2_26 < _issue2_idx_T_143 ? age_considering_issue_2_26 :
    _issue2_idx_T_143; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_149 = age_considering_issue_2_25 < _issue2_idx_T_147 ? 6'h19 : _issue2_idx_T_145; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_151 = age_considering_issue_2_25 < _issue2_idx_T_147 ? age_considering_issue_2_25 :
    _issue2_idx_T_147; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_153 = age_considering_issue_2_24 < _issue2_idx_T_151 ? 6'h18 : _issue2_idx_T_149; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_155 = age_considering_issue_2_24 < _issue2_idx_T_151 ? age_considering_issue_2_24 :
    _issue2_idx_T_151; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_157 = age_considering_issue_2_23 < _issue2_idx_T_155 ? 6'h17 : _issue2_idx_T_153; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_159 = age_considering_issue_2_23 < _issue2_idx_T_155 ? age_considering_issue_2_23 :
    _issue2_idx_T_155; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_161 = age_considering_issue_2_22 < _issue2_idx_T_159 ? 6'h16 : _issue2_idx_T_157; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_163 = age_considering_issue_2_22 < _issue2_idx_T_159 ? age_considering_issue_2_22 :
    _issue2_idx_T_159; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_165 = age_considering_issue_2_21 < _issue2_idx_T_163 ? 6'h15 : _issue2_idx_T_161; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_167 = age_considering_issue_2_21 < _issue2_idx_T_163 ? age_considering_issue_2_21 :
    _issue2_idx_T_163; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_169 = age_considering_issue_2_20 < _issue2_idx_T_167 ? 6'h14 : _issue2_idx_T_165; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_171 = age_considering_issue_2_20 < _issue2_idx_T_167 ? age_considering_issue_2_20 :
    _issue2_idx_T_167; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_173 = age_considering_issue_2_19 < _issue2_idx_T_171 ? 6'h13 : _issue2_idx_T_169; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_175 = age_considering_issue_2_19 < _issue2_idx_T_171 ? age_considering_issue_2_19 :
    _issue2_idx_T_171; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_177 = age_considering_issue_2_18 < _issue2_idx_T_175 ? 6'h12 : _issue2_idx_T_173; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_179 = age_considering_issue_2_18 < _issue2_idx_T_175 ? age_considering_issue_2_18 :
    _issue2_idx_T_175; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_181 = age_considering_issue_2_17 < _issue2_idx_T_179 ? 6'h11 : _issue2_idx_T_177; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_183 = age_considering_issue_2_17 < _issue2_idx_T_179 ? age_considering_issue_2_17 :
    _issue2_idx_T_179; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_185 = age_considering_issue_2_16 < _issue2_idx_T_183 ? 6'h10 : _issue2_idx_T_181; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_187 = age_considering_issue_2_16 < _issue2_idx_T_183 ? age_considering_issue_2_16 :
    _issue2_idx_T_183; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_189 = age_considering_issue_2_15 < _issue2_idx_T_187 ? 6'hf : _issue2_idx_T_185; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_191 = age_considering_issue_2_15 < _issue2_idx_T_187 ? age_considering_issue_2_15 :
    _issue2_idx_T_187; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_193 = age_considering_issue_2_14 < _issue2_idx_T_191 ? 6'he : _issue2_idx_T_189; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_195 = age_considering_issue_2_14 < _issue2_idx_T_191 ? age_considering_issue_2_14 :
    _issue2_idx_T_191; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_197 = age_considering_issue_2_13 < _issue2_idx_T_195 ? 6'hd : _issue2_idx_T_193; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_199 = age_considering_issue_2_13 < _issue2_idx_T_195 ? age_considering_issue_2_13 :
    _issue2_idx_T_195; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_201 = age_considering_issue_2_12 < _issue2_idx_T_199 ? 6'hc : _issue2_idx_T_197; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_203 = age_considering_issue_2_12 < _issue2_idx_T_199 ? age_considering_issue_2_12 :
    _issue2_idx_T_199; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_205 = age_considering_issue_2_11 < _issue2_idx_T_203 ? 6'hb : _issue2_idx_T_201; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_207 = age_considering_issue_2_11 < _issue2_idx_T_203 ? age_considering_issue_2_11 :
    _issue2_idx_T_203; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_209 = age_considering_issue_2_10 < _issue2_idx_T_207 ? 6'ha : _issue2_idx_T_205; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_211 = age_considering_issue_2_10 < _issue2_idx_T_207 ? age_considering_issue_2_10 :
    _issue2_idx_T_207; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_213 = age_considering_issue_2_9 < _issue2_idx_T_211 ? 6'h9 : _issue2_idx_T_209; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_215 = age_considering_issue_2_9 < _issue2_idx_T_211 ? age_considering_issue_2_9 :
    _issue2_idx_T_211; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_217 = age_considering_issue_2_8 < _issue2_idx_T_215 ? 6'h8 : _issue2_idx_T_213; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_219 = age_considering_issue_2_8 < _issue2_idx_T_215 ? age_considering_issue_2_8 :
    _issue2_idx_T_215; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_221 = age_considering_issue_2_7 < _issue2_idx_T_219 ? 6'h7 : _issue2_idx_T_217; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_223 = age_considering_issue_2_7 < _issue2_idx_T_219 ? age_considering_issue_2_7 :
    _issue2_idx_T_219; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_225 = age_considering_issue_2_6 < _issue2_idx_T_223 ? 6'h6 : _issue2_idx_T_221; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_227 = age_considering_issue_2_6 < _issue2_idx_T_223 ? age_considering_issue_2_6 :
    _issue2_idx_T_223; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_229 = age_considering_issue_2_5 < _issue2_idx_T_227 ? 6'h5 : _issue2_idx_T_225; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_231 = age_considering_issue_2_5 < _issue2_idx_T_227 ? age_considering_issue_2_5 :
    _issue2_idx_T_227; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_233 = age_considering_issue_2_4 < _issue2_idx_T_231 ? 6'h4 : _issue2_idx_T_229; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_235 = age_considering_issue_2_4 < _issue2_idx_T_231 ? age_considering_issue_2_4 :
    _issue2_idx_T_231; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_237 = age_considering_issue_2_3 < _issue2_idx_T_235 ? 6'h3 : _issue2_idx_T_233; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_239 = age_considering_issue_2_3 < _issue2_idx_T_235 ? age_considering_issue_2_3 :
    _issue2_idx_T_235; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_241 = age_considering_issue_2_2 < _issue2_idx_T_239 ? 6'h2 : _issue2_idx_T_237; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_243 = age_considering_issue_2_2 < _issue2_idx_T_239 ? age_considering_issue_2_2 :
    _issue2_idx_T_239; // @[reservation_station.scala 164:85]
  wire [5:0] _issue2_idx_T_245 = age_considering_issue_2_1 < _issue2_idx_T_243 ? 6'h1 : _issue2_idx_T_241; // @[reservation_station.scala 164:60]
  wire [7:0] _issue2_idx_T_247 = age_considering_issue_2_1 < _issue2_idx_T_243 ? age_considering_issue_2_1 :
    _issue2_idx_T_243; // @[reservation_station.scala 164:85]
  wire [5:0] issue2_idx = age_considering_issue_2_0 < _issue2_idx_T_247 ? 6'h0 : _issue2_idx_T_245; // @[reservation_station.scala 164:60]
  wire  _issue_num_T = issue1_idx == 6'h3f; // @[reservation_station.scala 168:21]
  wire  _issue_num_T_1 = issue2_idx == 6'h3f; // @[reservation_station.scala 168:42]
  wire  _issue_num_T_2 = issue1_idx == 6'h3f & issue2_idx == 6'h3f; // @[reservation_station.scala 168:29]
  wire  _issue_num_T_4 = issue2_idx != 6'h3f; // @[reservation_station.scala 169:43]
  wire  _issue_num_T_6 = issue1_idx != 6'h3f; // @[reservation_station.scala 169:66]
  wire  _issue_num_T_9 = _issue_num_T & issue2_idx != 6'h3f | issue1_idx != 6'h3f & _issue_num_T_1; // @[reservation_station.scala 169:52]
  wire  _issue_num_T_12 = _issue_num_T_6 & _issue_num_T_4; // @[reservation_station.scala 170:29]
  wire [1:0] _issue_num_T_13 = _issue_num_T_12 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _issue_num_T_14 = _issue_num_T_9 ? 2'h1 : _issue_num_T_13; // @[Mux.scala 101:16]
  wire [1:0] issue_num = _issue_num_T_2 ? 2'h0 : _issue_num_T_14; // @[Mux.scala 101:16]
  reg  issued_age_pack_issue_valid_0; // @[reservation_station.scala 173:35]
  reg  issued_age_pack_issue_valid_1; // @[reservation_station.scala 173:35]
  reg [7:0] issued_age_pack_max_age; // @[reservation_station.scala 173:35]
  reg [7:0] issued_age_pack_issued_ages_0; // @[reservation_station.scala 173:35]
  reg [7:0] issued_age_pack_issued_ages_1; // @[reservation_station.scala 173:35]
  wire  _issue0_valid_T_1 = issue_num == 2'h2; // @[reservation_station.scala 177:51]
  wire  issue0_valid = issue_num == 2'h1 | issue_num == 2'h2; // @[reservation_station.scala 177:38]
  wire  _write_num_T_2 = write_idx1 == 6'h3f | write_idx2 == 6'h3f; // @[reservation_station.scala 182:29]
  wire  _write_num_T_6 = ~_write_num_T_2; // @[reservation_station.scala 183:11]
  wire  _write_num_T_8 = ~_write_num_T_2 & (io_i_dispatch_packs_0_valid & io_i_dispatch_packs_1_valid); // @[reservation_station.scala 183:53]
  wire  _write_num_T_18 = _write_num_T_6 & (io_i_dispatch_packs_0_valid & ~io_i_dispatch_packs_1_valid | ~
    io_i_dispatch_packs_0_valid & io_i_dispatch_packs_1_valid); // @[reservation_station.scala 184:53]
  wire [1:0] _write_num_T_20 = _write_num_T_8 ? 2'h2 : {{1'd0}, _write_num_T_18}; // @[Mux.scala 101:16]
  wire [1:0] write_num = _write_num_T_2 ? 2'h0 : _write_num_T_20; // @[Mux.scala 101:16]
  wire [7:0] _GEN_21 = {{6'd0}, issue_num}; // @[reservation_station.scala 220:46]
  wire [7:0] _max_age_temp_T_1 = issued_age_pack_max_age - _GEN_21; // @[reservation_station.scala 220:46]
  wire [7:0] _GEN_22 = {{6'd0}, write_num}; // @[reservation_station.scala 220:58]
  wire [7:0] max_age_temp = _max_age_temp_T_1 + _GEN_22; // @[reservation_station.scala 220:58]
  wire [7:0] _issued_age_pack_issued_ages_0_T_64 = _issue1_func_code_T_63 ? reservation_station_63_io_o_age : 8'h3f; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_65 = _issue1_func_code_T_62 ? reservation_station_62_io_o_age :
    _issued_age_pack_issued_ages_0_T_64; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_66 = _issue1_func_code_T_61 ? reservation_station_61_io_o_age :
    _issued_age_pack_issued_ages_0_T_65; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_67 = _issue1_func_code_T_60 ? reservation_station_60_io_o_age :
    _issued_age_pack_issued_ages_0_T_66; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_68 = _issue1_func_code_T_59 ? reservation_station_59_io_o_age :
    _issued_age_pack_issued_ages_0_T_67; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_69 = _issue1_func_code_T_58 ? reservation_station_58_io_o_age :
    _issued_age_pack_issued_ages_0_T_68; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_70 = _issue1_func_code_T_57 ? reservation_station_57_io_o_age :
    _issued_age_pack_issued_ages_0_T_69; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_71 = _issue1_func_code_T_56 ? reservation_station_56_io_o_age :
    _issued_age_pack_issued_ages_0_T_70; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_72 = _issue1_func_code_T_55 ? reservation_station_55_io_o_age :
    _issued_age_pack_issued_ages_0_T_71; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_73 = _issue1_func_code_T_54 ? reservation_station_54_io_o_age :
    _issued_age_pack_issued_ages_0_T_72; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_74 = _issue1_func_code_T_53 ? reservation_station_53_io_o_age :
    _issued_age_pack_issued_ages_0_T_73; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_75 = _issue1_func_code_T_52 ? reservation_station_52_io_o_age :
    _issued_age_pack_issued_ages_0_T_74; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_76 = _issue1_func_code_T_51 ? reservation_station_51_io_o_age :
    _issued_age_pack_issued_ages_0_T_75; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_77 = _issue1_func_code_T_50 ? reservation_station_50_io_o_age :
    _issued_age_pack_issued_ages_0_T_76; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_78 = _issue1_func_code_T_49 ? reservation_station_49_io_o_age :
    _issued_age_pack_issued_ages_0_T_77; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_79 = _issue1_func_code_T_48 ? reservation_station_48_io_o_age :
    _issued_age_pack_issued_ages_0_T_78; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_80 = _issue1_func_code_T_47 ? reservation_station_47_io_o_age :
    _issued_age_pack_issued_ages_0_T_79; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_81 = _issue1_func_code_T_46 ? reservation_station_46_io_o_age :
    _issued_age_pack_issued_ages_0_T_80; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_82 = _issue1_func_code_T_45 ? reservation_station_45_io_o_age :
    _issued_age_pack_issued_ages_0_T_81; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_83 = _issue1_func_code_T_44 ? reservation_station_44_io_o_age :
    _issued_age_pack_issued_ages_0_T_82; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_84 = _issue1_func_code_T_43 ? reservation_station_43_io_o_age :
    _issued_age_pack_issued_ages_0_T_83; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_85 = _issue1_func_code_T_42 ? reservation_station_42_io_o_age :
    _issued_age_pack_issued_ages_0_T_84; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_86 = _issue1_func_code_T_41 ? reservation_station_41_io_o_age :
    _issued_age_pack_issued_ages_0_T_85; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_87 = _issue1_func_code_T_40 ? reservation_station_40_io_o_age :
    _issued_age_pack_issued_ages_0_T_86; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_88 = _issue1_func_code_T_39 ? reservation_station_39_io_o_age :
    _issued_age_pack_issued_ages_0_T_87; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_89 = _issue1_func_code_T_38 ? reservation_station_38_io_o_age :
    _issued_age_pack_issued_ages_0_T_88; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_90 = _issue1_func_code_T_37 ? reservation_station_37_io_o_age :
    _issued_age_pack_issued_ages_0_T_89; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_91 = _issue1_func_code_T_36 ? reservation_station_36_io_o_age :
    _issued_age_pack_issued_ages_0_T_90; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_92 = _issue1_func_code_T_35 ? reservation_station_35_io_o_age :
    _issued_age_pack_issued_ages_0_T_91; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_93 = _issue1_func_code_T_34 ? reservation_station_34_io_o_age :
    _issued_age_pack_issued_ages_0_T_92; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_94 = _issue1_func_code_T_33 ? reservation_station_33_io_o_age :
    _issued_age_pack_issued_ages_0_T_93; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_95 = _issue1_func_code_T_32 ? reservation_station_32_io_o_age :
    _issued_age_pack_issued_ages_0_T_94; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_96 = _issue1_func_code_T_31 ? reservation_station_31_io_o_age :
    _issued_age_pack_issued_ages_0_T_95; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_97 = _issue1_func_code_T_30 ? reservation_station_30_io_o_age :
    _issued_age_pack_issued_ages_0_T_96; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_98 = _issue1_func_code_T_29 ? reservation_station_29_io_o_age :
    _issued_age_pack_issued_ages_0_T_97; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_99 = _issue1_func_code_T_28 ? reservation_station_28_io_o_age :
    _issued_age_pack_issued_ages_0_T_98; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_100 = _issue1_func_code_T_27 ? reservation_station_27_io_o_age :
    _issued_age_pack_issued_ages_0_T_99; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_101 = _issue1_func_code_T_26 ? reservation_station_26_io_o_age :
    _issued_age_pack_issued_ages_0_T_100; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_102 = _issue1_func_code_T_25 ? reservation_station_25_io_o_age :
    _issued_age_pack_issued_ages_0_T_101; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_103 = _issue1_func_code_T_24 ? reservation_station_24_io_o_age :
    _issued_age_pack_issued_ages_0_T_102; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_104 = _issue1_func_code_T_23 ? reservation_station_23_io_o_age :
    _issued_age_pack_issued_ages_0_T_103; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_105 = _issue1_func_code_T_22 ? reservation_station_22_io_o_age :
    _issued_age_pack_issued_ages_0_T_104; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_106 = _issue1_func_code_T_21 ? reservation_station_21_io_o_age :
    _issued_age_pack_issued_ages_0_T_105; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_107 = _issue1_func_code_T_20 ? reservation_station_20_io_o_age :
    _issued_age_pack_issued_ages_0_T_106; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_108 = _issue1_func_code_T_19 ? reservation_station_19_io_o_age :
    _issued_age_pack_issued_ages_0_T_107; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_109 = _issue1_func_code_T_18 ? reservation_station_18_io_o_age :
    _issued_age_pack_issued_ages_0_T_108; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_110 = _issue1_func_code_T_17 ? reservation_station_17_io_o_age :
    _issued_age_pack_issued_ages_0_T_109; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_111 = _issue1_func_code_T_16 ? reservation_station_16_io_o_age :
    _issued_age_pack_issued_ages_0_T_110; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_112 = _issue1_func_code_T_15 ? reservation_station_15_io_o_age :
    _issued_age_pack_issued_ages_0_T_111; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_113 = _issue1_func_code_T_14 ? reservation_station_14_io_o_age :
    _issued_age_pack_issued_ages_0_T_112; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_114 = _issue1_func_code_T_13 ? reservation_station_13_io_o_age :
    _issued_age_pack_issued_ages_0_T_113; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_115 = _issue1_func_code_T_12 ? reservation_station_12_io_o_age :
    _issued_age_pack_issued_ages_0_T_114; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_116 = _issue1_func_code_T_11 ? reservation_station_11_io_o_age :
    _issued_age_pack_issued_ages_0_T_115; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_117 = _issue1_func_code_T_10 ? reservation_station_10_io_o_age :
    _issued_age_pack_issued_ages_0_T_116; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_118 = _issue1_func_code_T_9 ? reservation_station_9_io_o_age :
    _issued_age_pack_issued_ages_0_T_117; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_119 = _issue1_func_code_T_8 ? reservation_station_8_io_o_age :
    _issued_age_pack_issued_ages_0_T_118; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_120 = _issue1_func_code_T_7 ? reservation_station_7_io_o_age :
    _issued_age_pack_issued_ages_0_T_119; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_121 = _issue1_func_code_T_6 ? reservation_station_6_io_o_age :
    _issued_age_pack_issued_ages_0_T_120; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_122 = _issue1_func_code_T_5 ? reservation_station_5_io_o_age :
    _issued_age_pack_issued_ages_0_T_121; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_123 = _issue1_func_code_T_4 ? reservation_station_4_io_o_age :
    _issued_age_pack_issued_ages_0_T_122; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_124 = _issue1_func_code_T_3 ? reservation_station_3_io_o_age :
    _issued_age_pack_issued_ages_0_T_123; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_0_T_125 = _issue1_func_code_T_2 ? reservation_station_2_io_o_age :
    _issued_age_pack_issued_ages_0_T_124; // @[Mux.scala 101:16]
  wire  _issued_age_pack_issued_ages_1_T = 6'h0 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_1 = 6'h1 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_2 = 6'h2 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_3 = 6'h3 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_4 = 6'h4 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_5 = 6'h5 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_6 = 6'h6 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_7 = 6'h7 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_8 = 6'h8 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_9 = 6'h9 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_10 = 6'ha == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_11 = 6'hb == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_12 = 6'hc == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_13 = 6'hd == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_14 = 6'he == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_15 = 6'hf == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_16 = 6'h10 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_17 = 6'h11 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_18 = 6'h12 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_19 = 6'h13 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_20 = 6'h14 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_21 = 6'h15 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_22 = 6'h16 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_23 = 6'h17 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_24 = 6'h18 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_25 = 6'h19 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_26 = 6'h1a == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_27 = 6'h1b == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_28 = 6'h1c == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_29 = 6'h1d == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_30 = 6'h1e == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_31 = 6'h1f == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_32 = 6'h20 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_33 = 6'h21 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_34 = 6'h22 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_35 = 6'h23 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_36 = 6'h24 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_37 = 6'h25 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_38 = 6'h26 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_39 = 6'h27 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_40 = 6'h28 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_41 = 6'h29 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_42 = 6'h2a == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_43 = 6'h2b == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_44 = 6'h2c == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_45 = 6'h2d == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_46 = 6'h2e == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_47 = 6'h2f == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_48 = 6'h30 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_49 = 6'h31 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_50 = 6'h32 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_51 = 6'h33 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_52 = 6'h34 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_53 = 6'h35 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_54 = 6'h36 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_55 = 6'h37 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_56 = 6'h38 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_57 = 6'h39 == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_58 = 6'h3a == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_59 = 6'h3b == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_60 = 6'h3c == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_61 = 6'h3d == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_62 = 6'h3e == issue2_idx; // @[reservation_station.scala 228:80]
  wire  _issued_age_pack_issued_ages_1_T_63 = 6'h3f == issue2_idx; // @[reservation_station.scala 228:80]
  wire [7:0] _issued_age_pack_issued_ages_1_T_64 = _issued_age_pack_issued_ages_1_T_63 ? reservation_station_63_io_o_age
     : 8'h3f; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_65 = _issued_age_pack_issued_ages_1_T_62 ? reservation_station_62_io_o_age
     : _issued_age_pack_issued_ages_1_T_64; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_66 = _issued_age_pack_issued_ages_1_T_61 ? reservation_station_61_io_o_age
     : _issued_age_pack_issued_ages_1_T_65; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_67 = _issued_age_pack_issued_ages_1_T_60 ? reservation_station_60_io_o_age
     : _issued_age_pack_issued_ages_1_T_66; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_68 = _issued_age_pack_issued_ages_1_T_59 ? reservation_station_59_io_o_age
     : _issued_age_pack_issued_ages_1_T_67; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_69 = _issued_age_pack_issued_ages_1_T_58 ? reservation_station_58_io_o_age
     : _issued_age_pack_issued_ages_1_T_68; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_70 = _issued_age_pack_issued_ages_1_T_57 ? reservation_station_57_io_o_age
     : _issued_age_pack_issued_ages_1_T_69; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_71 = _issued_age_pack_issued_ages_1_T_56 ? reservation_station_56_io_o_age
     : _issued_age_pack_issued_ages_1_T_70; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_72 = _issued_age_pack_issued_ages_1_T_55 ? reservation_station_55_io_o_age
     : _issued_age_pack_issued_ages_1_T_71; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_73 = _issued_age_pack_issued_ages_1_T_54 ? reservation_station_54_io_o_age
     : _issued_age_pack_issued_ages_1_T_72; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_74 = _issued_age_pack_issued_ages_1_T_53 ? reservation_station_53_io_o_age
     : _issued_age_pack_issued_ages_1_T_73; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_75 = _issued_age_pack_issued_ages_1_T_52 ? reservation_station_52_io_o_age
     : _issued_age_pack_issued_ages_1_T_74; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_76 = _issued_age_pack_issued_ages_1_T_51 ? reservation_station_51_io_o_age
     : _issued_age_pack_issued_ages_1_T_75; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_77 = _issued_age_pack_issued_ages_1_T_50 ? reservation_station_50_io_o_age
     : _issued_age_pack_issued_ages_1_T_76; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_78 = _issued_age_pack_issued_ages_1_T_49 ? reservation_station_49_io_o_age
     : _issued_age_pack_issued_ages_1_T_77; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_79 = _issued_age_pack_issued_ages_1_T_48 ? reservation_station_48_io_o_age
     : _issued_age_pack_issued_ages_1_T_78; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_80 = _issued_age_pack_issued_ages_1_T_47 ? reservation_station_47_io_o_age
     : _issued_age_pack_issued_ages_1_T_79; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_81 = _issued_age_pack_issued_ages_1_T_46 ? reservation_station_46_io_o_age
     : _issued_age_pack_issued_ages_1_T_80; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_82 = _issued_age_pack_issued_ages_1_T_45 ? reservation_station_45_io_o_age
     : _issued_age_pack_issued_ages_1_T_81; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_83 = _issued_age_pack_issued_ages_1_T_44 ? reservation_station_44_io_o_age
     : _issued_age_pack_issued_ages_1_T_82; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_84 = _issued_age_pack_issued_ages_1_T_43 ? reservation_station_43_io_o_age
     : _issued_age_pack_issued_ages_1_T_83; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_85 = _issued_age_pack_issued_ages_1_T_42 ? reservation_station_42_io_o_age
     : _issued_age_pack_issued_ages_1_T_84; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_86 = _issued_age_pack_issued_ages_1_T_41 ? reservation_station_41_io_o_age
     : _issued_age_pack_issued_ages_1_T_85; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_87 = _issued_age_pack_issued_ages_1_T_40 ? reservation_station_40_io_o_age
     : _issued_age_pack_issued_ages_1_T_86; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_88 = _issued_age_pack_issued_ages_1_T_39 ? reservation_station_39_io_o_age
     : _issued_age_pack_issued_ages_1_T_87; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_89 = _issued_age_pack_issued_ages_1_T_38 ? reservation_station_38_io_o_age
     : _issued_age_pack_issued_ages_1_T_88; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_90 = _issued_age_pack_issued_ages_1_T_37 ? reservation_station_37_io_o_age
     : _issued_age_pack_issued_ages_1_T_89; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_91 = _issued_age_pack_issued_ages_1_T_36 ? reservation_station_36_io_o_age
     : _issued_age_pack_issued_ages_1_T_90; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_92 = _issued_age_pack_issued_ages_1_T_35 ? reservation_station_35_io_o_age
     : _issued_age_pack_issued_ages_1_T_91; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_93 = _issued_age_pack_issued_ages_1_T_34 ? reservation_station_34_io_o_age
     : _issued_age_pack_issued_ages_1_T_92; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_94 = _issued_age_pack_issued_ages_1_T_33 ? reservation_station_33_io_o_age
     : _issued_age_pack_issued_ages_1_T_93; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_95 = _issued_age_pack_issued_ages_1_T_32 ? reservation_station_32_io_o_age
     : _issued_age_pack_issued_ages_1_T_94; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_96 = _issued_age_pack_issued_ages_1_T_31 ? reservation_station_31_io_o_age
     : _issued_age_pack_issued_ages_1_T_95; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_97 = _issued_age_pack_issued_ages_1_T_30 ? reservation_station_30_io_o_age
     : _issued_age_pack_issued_ages_1_T_96; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_98 = _issued_age_pack_issued_ages_1_T_29 ? reservation_station_29_io_o_age
     : _issued_age_pack_issued_ages_1_T_97; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_99 = _issued_age_pack_issued_ages_1_T_28 ? reservation_station_28_io_o_age
     : _issued_age_pack_issued_ages_1_T_98; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_100 = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_age : _issued_age_pack_issued_ages_1_T_99; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_101 = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_age : _issued_age_pack_issued_ages_1_T_100; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_102 = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_age : _issued_age_pack_issued_ages_1_T_101; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_103 = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_age : _issued_age_pack_issued_ages_1_T_102; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_104 = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_age : _issued_age_pack_issued_ages_1_T_103; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_105 = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_age : _issued_age_pack_issued_ages_1_T_104; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_106 = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_age : _issued_age_pack_issued_ages_1_T_105; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_107 = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_age : _issued_age_pack_issued_ages_1_T_106; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_108 = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_age : _issued_age_pack_issued_ages_1_T_107; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_109 = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_age : _issued_age_pack_issued_ages_1_T_108; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_110 = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_age : _issued_age_pack_issued_ages_1_T_109; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_111 = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_age : _issued_age_pack_issued_ages_1_T_110; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_112 = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_age : _issued_age_pack_issued_ages_1_T_111; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_113 = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_age : _issued_age_pack_issued_ages_1_T_112; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_114 = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_age : _issued_age_pack_issued_ages_1_T_113; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_115 = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_age : _issued_age_pack_issued_ages_1_T_114; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_116 = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_age : _issued_age_pack_issued_ages_1_T_115; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_117 = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_age : _issued_age_pack_issued_ages_1_T_116; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_118 = _issued_age_pack_issued_ages_1_T_9 ? reservation_station_9_io_o_age
     : _issued_age_pack_issued_ages_1_T_117; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_119 = _issued_age_pack_issued_ages_1_T_8 ? reservation_station_8_io_o_age
     : _issued_age_pack_issued_ages_1_T_118; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_120 = _issued_age_pack_issued_ages_1_T_7 ? reservation_station_7_io_o_age
     : _issued_age_pack_issued_ages_1_T_119; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_121 = _issued_age_pack_issued_ages_1_T_6 ? reservation_station_6_io_o_age
     : _issued_age_pack_issued_ages_1_T_120; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_122 = _issued_age_pack_issued_ages_1_T_5 ? reservation_station_5_io_o_age
     : _issued_age_pack_issued_ages_1_T_121; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_123 = _issued_age_pack_issued_ages_1_T_4 ? reservation_station_4_io_o_age
     : _issued_age_pack_issued_ages_1_T_122; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_124 = _issued_age_pack_issued_ages_1_T_3 ? reservation_station_3_io_o_age
     : _issued_age_pack_issued_ages_1_T_123; // @[Mux.scala 101:16]
  wire [7:0] _issued_age_pack_issued_ages_1_T_125 = _issued_age_pack_issued_ages_1_T_2 ? reservation_station_2_io_o_age
     : _issued_age_pack_issued_ages_1_T_124; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_64_pc = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_pc :
    reservation_station_0_io_o_uop_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_64_inst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_inst :
    reservation_station_0_io_o_uop_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_func_code = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_func_code :
    reservation_station_0_io_o_uop_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_branch_predict_pack_valid = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_valid : reservation_station_0_io_o_uop_branch_predict_pack_valid
    ; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_branch_predict_pack_target = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_target :
    reservation_station_0_io_o_uop_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_64_branch_predict_pack_branch_type = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_branch_type :
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_branch_predict_pack_select = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_select :
    reservation_station_0_io_o_uop_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_branch_predict_pack_taken = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_taken : reservation_station_0_io_o_uop_branch_predict_pack_taken
    ; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_phy_dst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_phy_dst :
    reservation_station_0_io_o_uop_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_stale_dst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_stale_dst :
    reservation_station_0_io_o_uop_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_arch_dst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_arch_dst :
    reservation_station_0_io_o_uop_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_64_inst_type = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_inst_type :
    reservation_station_0_io_o_uop_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_regWen = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_regWen :
    reservation_station_0_io_o_uop_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_src1_valid = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src1_valid :
    reservation_station_0_io_o_uop_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_phy_rs1 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_phy_rs1 :
    reservation_station_0_io_o_uop_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_arch_rs1 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_arch_rs1 :
    reservation_station_0_io_o_uop_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_src2_valid = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src2_valid :
    reservation_station_0_io_o_uop_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_phy_rs2 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_phy_rs2 :
    reservation_station_0_io_o_uop_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_arch_rs2 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_arch_rs2 :
    reservation_station_0_io_o_uop_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_rob_idx = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_rob_idx :
    reservation_station_0_io_o_uop_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_imm = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_imm :
    reservation_station_0_io_o_uop_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_src1_value = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src1_value
     : reservation_station_0_io_o_uop_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_src2_value = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src2_value
     : reservation_station_0_io_o_uop_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_64_op1_sel = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_op1_sel :
    reservation_station_0_io_o_uop_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_64_op2_sel = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_op2_sel :
    reservation_station_0_io_o_uop_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_alu_sel = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_alu_sel :
    reservation_station_0_io_o_uop_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_64_branch_type = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_branch_type
     : reservation_station_0_io_o_uop_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_64_mem_type = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_mem_type :
    reservation_station_0_io_o_uop_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_65_pc = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_pc :
    _io_o_issue_packs_0_T_64_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_65_inst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_inst :
    _io_o_issue_packs_0_T_64_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_func_code = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_func_code :
    _io_o_issue_packs_0_T_64_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_branch_predict_pack_valid = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_64_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_branch_predict_pack_target = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_64_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_65_branch_predict_pack_branch_type = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_64_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_branch_predict_pack_select = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_64_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_branch_predict_pack_taken = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_64_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_phy_dst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_64_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_stale_dst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_64_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_arch_dst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_64_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_65_inst_type = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_64_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_regWen = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_regWen :
    _io_o_issue_packs_0_T_64_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_src1_valid = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_64_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_phy_rs1 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_64_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_arch_rs1 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_64_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_src2_valid = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_64_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_phy_rs2 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_64_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_arch_rs2 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_64_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_rob_idx = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_64_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_imm = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_imm :
    _io_o_issue_packs_0_T_64_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_src1_value = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_64_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_src2_value = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_64_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_65_op1_sel = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_64_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_65_op2_sel = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_64_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_alu_sel = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_64_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_65_branch_type = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_64_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_65_mem_type = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_64_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_66_pc = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_pc :
    _io_o_issue_packs_0_T_65_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_66_inst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_inst :
    _io_o_issue_packs_0_T_65_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_func_code = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_func_code :
    _io_o_issue_packs_0_T_65_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_branch_predict_pack_valid = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_65_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_branch_predict_pack_target = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_65_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_66_branch_predict_pack_branch_type = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_65_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_branch_predict_pack_select = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_65_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_branch_predict_pack_taken = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_65_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_phy_dst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_65_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_stale_dst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_65_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_arch_dst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_65_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_66_inst_type = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_65_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_regWen = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_regWen :
    _io_o_issue_packs_0_T_65_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_src1_valid = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_65_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_phy_rs1 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_65_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_arch_rs1 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_65_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_src2_valid = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_65_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_phy_rs2 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_65_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_arch_rs2 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_65_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_rob_idx = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_65_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_imm = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_imm :
    _io_o_issue_packs_0_T_65_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_src1_value = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_65_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_src2_value = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_65_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_66_op1_sel = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_65_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_66_op2_sel = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_65_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_alu_sel = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_65_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_66_branch_type = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_65_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_66_mem_type = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_65_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_67_pc = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_pc :
    _io_o_issue_packs_0_T_66_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_67_inst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_inst :
    _io_o_issue_packs_0_T_66_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_func_code = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_func_code :
    _io_o_issue_packs_0_T_66_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_branch_predict_pack_valid = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_66_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_branch_predict_pack_target = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_66_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_67_branch_predict_pack_branch_type = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_66_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_branch_predict_pack_select = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_66_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_branch_predict_pack_taken = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_66_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_phy_dst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_66_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_stale_dst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_66_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_arch_dst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_66_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_67_inst_type = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_66_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_regWen = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_regWen :
    _io_o_issue_packs_0_T_66_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_src1_valid = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_66_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_phy_rs1 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_66_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_arch_rs1 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_66_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_src2_valid = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_66_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_phy_rs2 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_66_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_arch_rs2 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_66_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_rob_idx = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_66_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_imm = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_imm :
    _io_o_issue_packs_0_T_66_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_src1_value = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_66_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_src2_value = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_66_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_67_op1_sel = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_66_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_67_op2_sel = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_66_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_alu_sel = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_66_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_67_branch_type = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_66_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_67_mem_type = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_66_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_68_pc = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_pc :
    _io_o_issue_packs_0_T_67_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_68_inst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_inst :
    _io_o_issue_packs_0_T_67_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_func_code = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_func_code :
    _io_o_issue_packs_0_T_67_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_branch_predict_pack_valid = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_67_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_branch_predict_pack_target = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_67_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_68_branch_predict_pack_branch_type = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_67_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_branch_predict_pack_select = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_67_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_branch_predict_pack_taken = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_67_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_phy_dst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_67_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_stale_dst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_67_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_arch_dst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_67_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_68_inst_type = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_67_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_regWen = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_regWen :
    _io_o_issue_packs_0_T_67_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_src1_valid = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_67_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_phy_rs1 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_67_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_arch_rs1 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_67_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_src2_valid = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_67_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_phy_rs2 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_67_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_arch_rs2 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_67_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_rob_idx = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_67_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_imm = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_imm :
    _io_o_issue_packs_0_T_67_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_src1_value = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_67_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_src2_value = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_67_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_68_op1_sel = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_67_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_68_op2_sel = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_67_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_alu_sel = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_67_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_68_branch_type = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_67_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_68_mem_type = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_67_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_69_pc = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_pc :
    _io_o_issue_packs_0_T_68_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_69_inst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_inst :
    _io_o_issue_packs_0_T_68_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_func_code = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_func_code :
    _io_o_issue_packs_0_T_68_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_branch_predict_pack_valid = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_68_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_branch_predict_pack_target = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_68_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_69_branch_predict_pack_branch_type = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_68_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_branch_predict_pack_select = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_68_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_branch_predict_pack_taken = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_68_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_phy_dst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_68_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_stale_dst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_68_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_arch_dst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_68_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_69_inst_type = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_68_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_regWen = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_regWen :
    _io_o_issue_packs_0_T_68_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_src1_valid = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_68_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_phy_rs1 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_68_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_arch_rs1 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_68_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_src2_valid = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_68_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_phy_rs2 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_68_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_arch_rs2 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_68_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_rob_idx = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_68_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_imm = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_imm :
    _io_o_issue_packs_0_T_68_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_src1_value = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_68_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_src2_value = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_68_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_69_op1_sel = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_68_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_69_op2_sel = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_68_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_alu_sel = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_68_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_69_branch_type = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_68_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_69_mem_type = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_68_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_70_pc = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_pc :
    _io_o_issue_packs_0_T_69_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_70_inst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_inst :
    _io_o_issue_packs_0_T_69_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_func_code = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_func_code :
    _io_o_issue_packs_0_T_69_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_branch_predict_pack_valid = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_69_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_branch_predict_pack_target = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_69_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_70_branch_predict_pack_branch_type = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_69_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_branch_predict_pack_select = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_69_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_branch_predict_pack_taken = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_69_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_phy_dst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_69_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_stale_dst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_69_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_arch_dst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_69_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_70_inst_type = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_69_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_regWen = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_regWen :
    _io_o_issue_packs_0_T_69_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_src1_valid = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_69_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_phy_rs1 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_69_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_arch_rs1 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_69_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_src2_valid = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_69_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_phy_rs2 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_69_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_arch_rs2 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_69_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_rob_idx = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_69_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_imm = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_imm :
    _io_o_issue_packs_0_T_69_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_src1_value = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_69_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_src2_value = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_69_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_70_op1_sel = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_69_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_70_op2_sel = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_69_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_alu_sel = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_69_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_70_branch_type = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_69_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_70_mem_type = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_69_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_71_pc = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_pc :
    _io_o_issue_packs_0_T_70_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_71_inst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_inst :
    _io_o_issue_packs_0_T_70_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_func_code = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_func_code :
    _io_o_issue_packs_0_T_70_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_branch_predict_pack_valid = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_70_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_branch_predict_pack_target = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_70_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_71_branch_predict_pack_branch_type = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_70_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_branch_predict_pack_select = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_70_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_branch_predict_pack_taken = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_70_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_phy_dst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_70_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_stale_dst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_70_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_arch_dst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_70_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_71_inst_type = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_70_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_regWen = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_regWen :
    _io_o_issue_packs_0_T_70_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_src1_valid = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_70_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_phy_rs1 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_70_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_arch_rs1 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_70_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_src2_valid = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_70_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_phy_rs2 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_70_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_arch_rs2 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_70_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_rob_idx = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_70_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_imm = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_imm :
    _io_o_issue_packs_0_T_70_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_src1_value = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_70_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_src2_value = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_70_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_71_op1_sel = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_70_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_71_op2_sel = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_70_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_alu_sel = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_70_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_71_branch_type = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_70_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_71_mem_type = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_70_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_72_pc = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_pc :
    _io_o_issue_packs_0_T_71_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_72_inst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_inst :
    _io_o_issue_packs_0_T_71_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_func_code = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_func_code :
    _io_o_issue_packs_0_T_71_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_branch_predict_pack_valid = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_71_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_branch_predict_pack_target = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_71_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_72_branch_predict_pack_branch_type = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_71_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_branch_predict_pack_select = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_71_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_branch_predict_pack_taken = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_71_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_phy_dst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_71_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_stale_dst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_71_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_arch_dst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_71_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_72_inst_type = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_71_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_regWen = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_regWen :
    _io_o_issue_packs_0_T_71_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_src1_valid = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_71_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_phy_rs1 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_71_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_arch_rs1 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_71_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_src2_valid = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_71_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_phy_rs2 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_71_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_arch_rs2 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_71_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_rob_idx = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_71_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_imm = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_imm :
    _io_o_issue_packs_0_T_71_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_src1_value = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_71_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_src2_value = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_71_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_72_op1_sel = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_71_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_72_op2_sel = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_71_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_alu_sel = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_71_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_72_branch_type = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_71_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_72_mem_type = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_71_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_73_pc = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_pc :
    _io_o_issue_packs_0_T_72_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_73_inst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_inst :
    _io_o_issue_packs_0_T_72_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_func_code = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_func_code :
    _io_o_issue_packs_0_T_72_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_branch_predict_pack_valid = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_72_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_branch_predict_pack_target = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_72_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_73_branch_predict_pack_branch_type = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_72_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_branch_predict_pack_select = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_72_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_branch_predict_pack_taken = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_72_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_phy_dst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_72_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_stale_dst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_72_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_arch_dst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_72_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_73_inst_type = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_72_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_regWen = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_regWen :
    _io_o_issue_packs_0_T_72_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_src1_valid = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_72_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_phy_rs1 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_72_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_arch_rs1 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_72_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_src2_valid = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_72_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_phy_rs2 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_72_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_arch_rs2 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_72_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_rob_idx = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_72_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_imm = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_imm :
    _io_o_issue_packs_0_T_72_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_src1_value = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_72_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_src2_value = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_72_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_73_op1_sel = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_72_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_73_op2_sel = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_72_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_alu_sel = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_72_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_73_branch_type = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_72_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_73_mem_type = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_72_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_74_pc = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_pc :
    _io_o_issue_packs_0_T_73_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_74_inst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_inst :
    _io_o_issue_packs_0_T_73_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_func_code = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_func_code :
    _io_o_issue_packs_0_T_73_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_branch_predict_pack_valid = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_73_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_branch_predict_pack_target = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_73_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_74_branch_predict_pack_branch_type = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_73_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_branch_predict_pack_select = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_73_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_branch_predict_pack_taken = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_73_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_phy_dst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_73_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_stale_dst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_73_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_arch_dst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_73_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_74_inst_type = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_73_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_regWen = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_regWen :
    _io_o_issue_packs_0_T_73_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_src1_valid = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_73_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_phy_rs1 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_73_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_arch_rs1 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_73_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_src2_valid = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_73_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_phy_rs2 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_73_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_arch_rs2 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_73_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_rob_idx = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_73_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_imm = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_imm :
    _io_o_issue_packs_0_T_73_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_src1_value = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_73_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_src2_value = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_73_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_74_op1_sel = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_73_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_74_op2_sel = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_73_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_alu_sel = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_73_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_74_branch_type = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_73_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_74_mem_type = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_73_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_75_pc = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_pc :
    _io_o_issue_packs_0_T_74_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_75_inst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_inst :
    _io_o_issue_packs_0_T_74_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_func_code = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_func_code :
    _io_o_issue_packs_0_T_74_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_branch_predict_pack_valid = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_74_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_branch_predict_pack_target = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_74_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_75_branch_predict_pack_branch_type = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_74_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_branch_predict_pack_select = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_74_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_branch_predict_pack_taken = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_74_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_phy_dst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_74_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_stale_dst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_74_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_arch_dst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_74_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_75_inst_type = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_74_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_regWen = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_regWen :
    _io_o_issue_packs_0_T_74_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_src1_valid = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_74_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_phy_rs1 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_74_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_arch_rs1 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_74_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_src2_valid = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_74_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_phy_rs2 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_74_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_arch_rs2 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_74_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_rob_idx = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_74_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_imm = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_imm :
    _io_o_issue_packs_0_T_74_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_src1_value = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_74_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_src2_value = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_74_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_75_op1_sel = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_74_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_75_op2_sel = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_74_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_alu_sel = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_74_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_75_branch_type = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_74_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_75_mem_type = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_74_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_76_pc = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_pc :
    _io_o_issue_packs_0_T_75_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_76_inst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_inst :
    _io_o_issue_packs_0_T_75_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_func_code = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_func_code :
    _io_o_issue_packs_0_T_75_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_branch_predict_pack_valid = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_75_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_branch_predict_pack_target = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_75_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_76_branch_predict_pack_branch_type = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_75_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_branch_predict_pack_select = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_75_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_branch_predict_pack_taken = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_75_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_phy_dst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_75_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_stale_dst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_75_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_arch_dst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_75_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_76_inst_type = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_75_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_regWen = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_regWen :
    _io_o_issue_packs_0_T_75_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_src1_valid = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_75_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_phy_rs1 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_75_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_arch_rs1 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_75_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_src2_valid = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_75_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_phy_rs2 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_75_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_arch_rs2 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_75_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_rob_idx = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_75_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_imm = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_imm :
    _io_o_issue_packs_0_T_75_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_src1_value = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_75_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_src2_value = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_75_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_76_op1_sel = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_75_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_76_op2_sel = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_75_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_alu_sel = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_75_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_76_branch_type = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_75_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_76_mem_type = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_75_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_77_pc = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_pc :
    _io_o_issue_packs_0_T_76_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_77_inst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_inst :
    _io_o_issue_packs_0_T_76_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_func_code = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_func_code :
    _io_o_issue_packs_0_T_76_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_branch_predict_pack_valid = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_76_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_branch_predict_pack_target = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_76_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_77_branch_predict_pack_branch_type = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_76_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_branch_predict_pack_select = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_76_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_branch_predict_pack_taken = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_76_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_phy_dst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_76_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_stale_dst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_76_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_arch_dst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_76_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_77_inst_type = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_76_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_regWen = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_regWen :
    _io_o_issue_packs_0_T_76_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_src1_valid = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_76_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_phy_rs1 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_76_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_arch_rs1 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_76_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_src2_valid = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_76_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_phy_rs2 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_76_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_arch_rs2 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_76_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_rob_idx = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_76_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_imm = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_imm :
    _io_o_issue_packs_0_T_76_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_src1_value = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_76_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_src2_value = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_76_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_77_op1_sel = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_76_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_77_op2_sel = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_76_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_alu_sel = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_76_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_77_branch_type = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_76_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_77_mem_type = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_76_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_78_pc = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_pc :
    _io_o_issue_packs_0_T_77_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_78_inst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_inst :
    _io_o_issue_packs_0_T_77_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_func_code = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_func_code :
    _io_o_issue_packs_0_T_77_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_branch_predict_pack_valid = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_77_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_branch_predict_pack_target = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_77_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_78_branch_predict_pack_branch_type = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_77_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_branch_predict_pack_select = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_77_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_branch_predict_pack_taken = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_77_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_phy_dst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_77_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_stale_dst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_77_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_arch_dst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_77_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_78_inst_type = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_77_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_regWen = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_regWen :
    _io_o_issue_packs_0_T_77_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_src1_valid = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_77_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_phy_rs1 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_77_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_arch_rs1 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_77_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_src2_valid = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_77_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_phy_rs2 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_77_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_arch_rs2 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_77_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_rob_idx = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_77_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_imm = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_imm :
    _io_o_issue_packs_0_T_77_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_src1_value = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_77_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_src2_value = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_77_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_78_op1_sel = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_77_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_78_op2_sel = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_77_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_alu_sel = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_77_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_78_branch_type = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_77_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_78_mem_type = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_77_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_79_pc = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_pc :
    _io_o_issue_packs_0_T_78_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_79_inst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_inst :
    _io_o_issue_packs_0_T_78_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_func_code = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_func_code :
    _io_o_issue_packs_0_T_78_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_branch_predict_pack_valid = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_78_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_branch_predict_pack_target = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_78_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_79_branch_predict_pack_branch_type = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_78_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_branch_predict_pack_select = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_78_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_branch_predict_pack_taken = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_78_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_phy_dst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_78_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_stale_dst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_78_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_arch_dst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_78_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_79_inst_type = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_78_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_regWen = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_regWen :
    _io_o_issue_packs_0_T_78_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_src1_valid = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_78_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_phy_rs1 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_78_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_arch_rs1 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_78_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_src2_valid = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_78_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_phy_rs2 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_78_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_arch_rs2 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_78_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_rob_idx = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_78_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_imm = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_imm :
    _io_o_issue_packs_0_T_78_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_src1_value = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_78_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_src2_value = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_78_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_79_op1_sel = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_78_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_79_op2_sel = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_78_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_alu_sel = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_78_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_79_branch_type = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_78_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_79_mem_type = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_78_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_80_pc = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_pc :
    _io_o_issue_packs_0_T_79_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_80_inst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_inst :
    _io_o_issue_packs_0_T_79_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_func_code = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_func_code :
    _io_o_issue_packs_0_T_79_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_branch_predict_pack_valid = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_79_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_branch_predict_pack_target = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_79_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_80_branch_predict_pack_branch_type = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_79_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_branch_predict_pack_select = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_79_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_branch_predict_pack_taken = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_79_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_phy_dst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_79_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_stale_dst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_79_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_arch_dst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_79_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_80_inst_type = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_79_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_regWen = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_regWen :
    _io_o_issue_packs_0_T_79_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_src1_valid = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_79_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_phy_rs1 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_79_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_arch_rs1 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_79_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_src2_valid = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_79_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_phy_rs2 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_79_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_arch_rs2 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_79_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_rob_idx = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_79_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_imm = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_imm :
    _io_o_issue_packs_0_T_79_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_src1_value = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_79_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_src2_value = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_79_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_80_op1_sel = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_79_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_80_op2_sel = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_79_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_alu_sel = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_79_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_80_branch_type = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_79_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_80_mem_type = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_79_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_81_pc = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_pc :
    _io_o_issue_packs_0_T_80_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_81_inst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_inst :
    _io_o_issue_packs_0_T_80_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_func_code = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_func_code :
    _io_o_issue_packs_0_T_80_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_branch_predict_pack_valid = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_80_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_branch_predict_pack_target = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_80_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_81_branch_predict_pack_branch_type = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_80_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_branch_predict_pack_select = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_80_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_branch_predict_pack_taken = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_80_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_phy_dst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_80_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_stale_dst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_80_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_arch_dst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_80_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_81_inst_type = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_80_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_regWen = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_regWen :
    _io_o_issue_packs_0_T_80_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_src1_valid = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_80_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_phy_rs1 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_80_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_arch_rs1 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_80_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_src2_valid = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_80_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_phy_rs2 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_80_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_arch_rs2 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_80_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_rob_idx = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_80_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_imm = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_imm :
    _io_o_issue_packs_0_T_80_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_src1_value = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_80_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_src2_value = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_80_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_81_op1_sel = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_80_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_81_op2_sel = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_80_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_alu_sel = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_80_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_81_branch_type = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_80_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_81_mem_type = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_80_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_82_pc = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_pc :
    _io_o_issue_packs_0_T_81_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_82_inst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_inst :
    _io_o_issue_packs_0_T_81_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_func_code = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_func_code :
    _io_o_issue_packs_0_T_81_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_branch_predict_pack_valid = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_81_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_branch_predict_pack_target = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_81_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_82_branch_predict_pack_branch_type = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_81_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_branch_predict_pack_select = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_81_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_branch_predict_pack_taken = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_81_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_phy_dst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_81_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_stale_dst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_81_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_arch_dst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_81_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_82_inst_type = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_81_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_regWen = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_regWen :
    _io_o_issue_packs_0_T_81_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_src1_valid = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_81_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_phy_rs1 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_81_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_arch_rs1 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_81_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_src2_valid = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_81_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_phy_rs2 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_81_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_arch_rs2 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_81_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_rob_idx = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_81_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_imm = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_imm :
    _io_o_issue_packs_0_T_81_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_src1_value = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_81_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_src2_value = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_81_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_82_op1_sel = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_81_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_82_op2_sel = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_81_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_alu_sel = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_81_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_82_branch_type = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_81_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_82_mem_type = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_81_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_83_pc = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_pc :
    _io_o_issue_packs_0_T_82_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_83_inst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_inst :
    _io_o_issue_packs_0_T_82_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_func_code = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_func_code :
    _io_o_issue_packs_0_T_82_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_branch_predict_pack_valid = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_82_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_branch_predict_pack_target = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_82_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_83_branch_predict_pack_branch_type = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_82_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_branch_predict_pack_select = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_82_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_branch_predict_pack_taken = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_82_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_phy_dst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_82_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_stale_dst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_82_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_arch_dst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_82_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_83_inst_type = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_82_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_regWen = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_regWen :
    _io_o_issue_packs_0_T_82_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_src1_valid = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_82_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_phy_rs1 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_82_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_arch_rs1 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_82_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_src2_valid = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_82_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_phy_rs2 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_82_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_arch_rs2 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_82_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_rob_idx = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_82_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_imm = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_imm :
    _io_o_issue_packs_0_T_82_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_src1_value = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_82_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_src2_value = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_82_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_83_op1_sel = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_82_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_83_op2_sel = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_82_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_alu_sel = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_82_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_83_branch_type = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_82_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_83_mem_type = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_82_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_84_pc = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_pc :
    _io_o_issue_packs_0_T_83_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_84_inst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_inst :
    _io_o_issue_packs_0_T_83_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_func_code = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_func_code :
    _io_o_issue_packs_0_T_83_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_branch_predict_pack_valid = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_83_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_branch_predict_pack_target = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_83_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_84_branch_predict_pack_branch_type = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_83_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_branch_predict_pack_select = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_83_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_branch_predict_pack_taken = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_83_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_phy_dst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_83_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_stale_dst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_83_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_arch_dst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_83_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_84_inst_type = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_83_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_regWen = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_regWen :
    _io_o_issue_packs_0_T_83_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_src1_valid = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_83_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_phy_rs1 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_83_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_arch_rs1 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_83_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_src2_valid = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_83_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_phy_rs2 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_83_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_arch_rs2 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_83_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_rob_idx = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_83_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_imm = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_imm :
    _io_o_issue_packs_0_T_83_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_src1_value = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_83_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_src2_value = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_83_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_84_op1_sel = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_83_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_84_op2_sel = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_83_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_alu_sel = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_83_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_84_branch_type = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_83_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_84_mem_type = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_83_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_85_pc = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_pc :
    _io_o_issue_packs_0_T_84_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_85_inst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_inst :
    _io_o_issue_packs_0_T_84_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_func_code = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_func_code :
    _io_o_issue_packs_0_T_84_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_branch_predict_pack_valid = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_84_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_branch_predict_pack_target = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_84_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_85_branch_predict_pack_branch_type = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_84_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_branch_predict_pack_select = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_84_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_branch_predict_pack_taken = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_84_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_phy_dst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_84_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_stale_dst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_84_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_arch_dst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_84_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_85_inst_type = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_84_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_regWen = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_regWen :
    _io_o_issue_packs_0_T_84_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_src1_valid = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_84_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_phy_rs1 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_84_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_arch_rs1 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_84_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_src2_valid = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_84_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_phy_rs2 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_84_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_arch_rs2 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_84_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_rob_idx = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_84_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_imm = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_imm :
    _io_o_issue_packs_0_T_84_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_src1_value = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_84_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_src2_value = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_84_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_85_op1_sel = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_84_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_85_op2_sel = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_84_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_alu_sel = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_84_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_85_branch_type = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_84_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_85_mem_type = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_84_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_86_pc = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_pc :
    _io_o_issue_packs_0_T_85_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_86_inst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_inst :
    _io_o_issue_packs_0_T_85_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_func_code = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_func_code :
    _io_o_issue_packs_0_T_85_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_branch_predict_pack_valid = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_85_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_branch_predict_pack_target = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_85_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_86_branch_predict_pack_branch_type = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_85_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_branch_predict_pack_select = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_85_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_branch_predict_pack_taken = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_85_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_phy_dst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_85_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_stale_dst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_85_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_arch_dst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_85_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_86_inst_type = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_85_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_regWen = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_regWen :
    _io_o_issue_packs_0_T_85_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_src1_valid = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_85_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_phy_rs1 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_85_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_arch_rs1 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_85_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_src2_valid = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_85_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_phy_rs2 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_85_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_arch_rs2 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_85_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_rob_idx = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_85_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_imm = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_imm :
    _io_o_issue_packs_0_T_85_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_src1_value = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_85_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_src2_value = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_85_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_86_op1_sel = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_85_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_86_op2_sel = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_85_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_alu_sel = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_85_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_86_branch_type = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_85_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_86_mem_type = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_85_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_87_pc = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_pc :
    _io_o_issue_packs_0_T_86_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_87_inst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_inst :
    _io_o_issue_packs_0_T_86_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_func_code = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_func_code :
    _io_o_issue_packs_0_T_86_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_branch_predict_pack_valid = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_86_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_branch_predict_pack_target = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_86_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_87_branch_predict_pack_branch_type = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_86_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_branch_predict_pack_select = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_86_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_branch_predict_pack_taken = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_86_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_phy_dst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_86_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_stale_dst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_86_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_arch_dst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_86_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_87_inst_type = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_86_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_regWen = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_regWen :
    _io_o_issue_packs_0_T_86_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_src1_valid = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_86_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_phy_rs1 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_86_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_arch_rs1 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_86_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_src2_valid = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_86_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_phy_rs2 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_86_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_arch_rs2 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_86_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_rob_idx = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_86_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_imm = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_imm :
    _io_o_issue_packs_0_T_86_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_src1_value = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_86_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_src2_value = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_86_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_87_op1_sel = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_86_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_87_op2_sel = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_86_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_alu_sel = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_86_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_87_branch_type = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_86_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_87_mem_type = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_86_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_88_pc = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_pc :
    _io_o_issue_packs_0_T_87_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_88_inst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_inst :
    _io_o_issue_packs_0_T_87_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_func_code = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_func_code :
    _io_o_issue_packs_0_T_87_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_branch_predict_pack_valid = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_87_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_branch_predict_pack_target = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_87_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_88_branch_predict_pack_branch_type = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_87_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_branch_predict_pack_select = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_87_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_branch_predict_pack_taken = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_87_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_phy_dst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_87_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_stale_dst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_87_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_arch_dst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_87_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_88_inst_type = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_87_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_regWen = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_regWen :
    _io_o_issue_packs_0_T_87_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_src1_valid = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_87_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_phy_rs1 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_87_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_arch_rs1 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_87_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_src2_valid = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_87_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_phy_rs2 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_87_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_arch_rs2 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_87_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_rob_idx = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_87_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_imm = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_imm :
    _io_o_issue_packs_0_T_87_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_src1_value = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_87_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_src2_value = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_87_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_88_op1_sel = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_87_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_88_op2_sel = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_87_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_alu_sel = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_87_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_88_branch_type = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_87_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_88_mem_type = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_87_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_89_pc = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_pc :
    _io_o_issue_packs_0_T_88_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_89_inst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_inst :
    _io_o_issue_packs_0_T_88_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_func_code = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_func_code :
    _io_o_issue_packs_0_T_88_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_branch_predict_pack_valid = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_88_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_branch_predict_pack_target = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_88_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_89_branch_predict_pack_branch_type = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_88_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_branch_predict_pack_select = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_88_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_branch_predict_pack_taken = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_88_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_phy_dst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_88_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_stale_dst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_88_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_arch_dst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_88_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_89_inst_type = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_88_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_regWen = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_regWen :
    _io_o_issue_packs_0_T_88_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_src1_valid = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_88_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_phy_rs1 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_88_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_arch_rs1 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_88_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_src2_valid = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_88_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_phy_rs2 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_88_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_arch_rs2 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_88_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_rob_idx = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_88_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_imm = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_imm :
    _io_o_issue_packs_0_T_88_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_src1_value = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_88_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_src2_value = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_88_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_89_op1_sel = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_88_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_89_op2_sel = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_88_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_alu_sel = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_88_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_89_branch_type = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_88_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_89_mem_type = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_88_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_90_pc = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_pc :
    _io_o_issue_packs_0_T_89_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_90_inst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_inst :
    _io_o_issue_packs_0_T_89_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_func_code = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_func_code :
    _io_o_issue_packs_0_T_89_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_branch_predict_pack_valid = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_89_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_branch_predict_pack_target = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_89_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_90_branch_predict_pack_branch_type = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_89_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_branch_predict_pack_select = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_89_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_branch_predict_pack_taken = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_89_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_phy_dst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_89_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_stale_dst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_89_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_arch_dst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_89_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_90_inst_type = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_89_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_regWen = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_regWen :
    _io_o_issue_packs_0_T_89_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_src1_valid = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_89_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_phy_rs1 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_89_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_arch_rs1 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_89_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_src2_valid = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_89_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_phy_rs2 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_89_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_arch_rs2 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_89_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_rob_idx = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_89_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_imm = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_imm :
    _io_o_issue_packs_0_T_89_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_src1_value = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_89_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_src2_value = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_89_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_90_op1_sel = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_89_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_90_op2_sel = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_89_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_alu_sel = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_89_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_90_branch_type = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_89_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_90_mem_type = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_89_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_91_pc = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_pc :
    _io_o_issue_packs_0_T_90_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_91_inst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_inst :
    _io_o_issue_packs_0_T_90_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_func_code = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_func_code :
    _io_o_issue_packs_0_T_90_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_branch_predict_pack_valid = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_90_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_branch_predict_pack_target = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_90_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_91_branch_predict_pack_branch_type = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_90_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_branch_predict_pack_select = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_90_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_branch_predict_pack_taken = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_90_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_phy_dst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_90_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_stale_dst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_90_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_arch_dst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_90_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_91_inst_type = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_90_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_regWen = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_regWen :
    _io_o_issue_packs_0_T_90_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_src1_valid = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_90_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_phy_rs1 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_90_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_arch_rs1 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_90_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_src2_valid = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_90_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_phy_rs2 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_90_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_arch_rs2 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_90_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_rob_idx = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_90_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_imm = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_imm :
    _io_o_issue_packs_0_T_90_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_src1_value = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_90_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_src2_value = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_90_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_91_op1_sel = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_90_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_91_op2_sel = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_90_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_alu_sel = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_90_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_91_branch_type = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_90_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_91_mem_type = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_90_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_92_pc = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_pc :
    _io_o_issue_packs_0_T_91_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_92_inst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_inst :
    _io_o_issue_packs_0_T_91_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_func_code = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_func_code :
    _io_o_issue_packs_0_T_91_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_branch_predict_pack_valid = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_91_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_branch_predict_pack_target = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_91_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_92_branch_predict_pack_branch_type = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_91_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_branch_predict_pack_select = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_91_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_branch_predict_pack_taken = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_91_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_phy_dst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_91_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_stale_dst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_91_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_arch_dst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_91_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_92_inst_type = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_91_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_regWen = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_regWen :
    _io_o_issue_packs_0_T_91_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_src1_valid = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_91_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_phy_rs1 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_91_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_arch_rs1 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_91_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_src2_valid = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_91_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_phy_rs2 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_91_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_arch_rs2 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_91_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_rob_idx = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_91_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_imm = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_imm :
    _io_o_issue_packs_0_T_91_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_src1_value = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_91_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_src2_value = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_91_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_92_op1_sel = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_91_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_92_op2_sel = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_91_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_alu_sel = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_91_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_92_branch_type = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_91_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_92_mem_type = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_91_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_93_pc = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_pc :
    _io_o_issue_packs_0_T_92_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_93_inst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_inst :
    _io_o_issue_packs_0_T_92_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_func_code = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_func_code :
    _io_o_issue_packs_0_T_92_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_branch_predict_pack_valid = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_92_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_branch_predict_pack_target = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_92_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_93_branch_predict_pack_branch_type = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_92_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_branch_predict_pack_select = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_92_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_branch_predict_pack_taken = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_92_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_phy_dst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_92_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_stale_dst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_92_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_arch_dst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_92_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_93_inst_type = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_92_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_regWen = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_regWen :
    _io_o_issue_packs_0_T_92_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_src1_valid = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_92_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_phy_rs1 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_92_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_arch_rs1 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_92_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_src2_valid = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_92_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_phy_rs2 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_92_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_arch_rs2 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_92_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_rob_idx = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_92_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_imm = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_imm :
    _io_o_issue_packs_0_T_92_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_src1_value = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_92_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_src2_value = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_92_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_93_op1_sel = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_92_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_93_op2_sel = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_92_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_alu_sel = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_92_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_93_branch_type = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_92_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_93_mem_type = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_92_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_94_pc = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_pc :
    _io_o_issue_packs_0_T_93_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_94_inst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_inst :
    _io_o_issue_packs_0_T_93_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_func_code = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_func_code :
    _io_o_issue_packs_0_T_93_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_branch_predict_pack_valid = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_93_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_branch_predict_pack_target = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_93_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_94_branch_predict_pack_branch_type = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_93_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_branch_predict_pack_select = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_93_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_branch_predict_pack_taken = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_93_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_phy_dst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_93_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_stale_dst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_93_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_arch_dst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_93_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_94_inst_type = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_93_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_regWen = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_regWen :
    _io_o_issue_packs_0_T_93_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_src1_valid = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_93_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_phy_rs1 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_93_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_arch_rs1 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_93_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_src2_valid = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_93_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_phy_rs2 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_93_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_arch_rs2 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_93_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_rob_idx = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_93_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_imm = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_imm :
    _io_o_issue_packs_0_T_93_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_src1_value = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_93_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_src2_value = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_93_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_94_op1_sel = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_93_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_94_op2_sel = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_93_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_alu_sel = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_93_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_94_branch_type = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_93_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_94_mem_type = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_93_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_95_pc = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_pc :
    _io_o_issue_packs_0_T_94_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_95_inst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_inst :
    _io_o_issue_packs_0_T_94_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_func_code = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_func_code :
    _io_o_issue_packs_0_T_94_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_branch_predict_pack_valid = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_94_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_branch_predict_pack_target = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_94_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_95_branch_predict_pack_branch_type = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_94_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_branch_predict_pack_select = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_94_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_branch_predict_pack_taken = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_94_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_phy_dst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_94_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_stale_dst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_94_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_arch_dst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_94_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_95_inst_type = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_94_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_regWen = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_regWen :
    _io_o_issue_packs_0_T_94_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_src1_valid = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_94_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_phy_rs1 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_94_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_arch_rs1 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_94_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_src2_valid = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_94_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_phy_rs2 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_94_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_arch_rs2 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_94_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_rob_idx = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_94_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_imm = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_imm :
    _io_o_issue_packs_0_T_94_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_src1_value = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_94_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_src2_value = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_94_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_95_op1_sel = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_94_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_95_op2_sel = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_94_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_alu_sel = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_94_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_95_branch_type = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_94_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_95_mem_type = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_94_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_96_pc = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_pc :
    _io_o_issue_packs_0_T_95_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_96_inst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_inst :
    _io_o_issue_packs_0_T_95_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_func_code = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_func_code :
    _io_o_issue_packs_0_T_95_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_branch_predict_pack_valid = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_95_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_branch_predict_pack_target = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_95_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_96_branch_predict_pack_branch_type = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_95_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_branch_predict_pack_select = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_95_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_branch_predict_pack_taken = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_95_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_phy_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_95_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_stale_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_95_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_arch_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_95_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_96_inst_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_95_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_regWen = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_regWen :
    _io_o_issue_packs_0_T_95_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_src1_valid = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_95_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_phy_rs1 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_95_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_arch_rs1 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_95_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_src2_valid = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_95_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_phy_rs2 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_95_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_arch_rs2 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_95_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_rob_idx = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_95_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_imm = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_imm :
    _io_o_issue_packs_0_T_95_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_src1_value = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_95_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_src2_value = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_95_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_96_op1_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_95_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_96_op2_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_95_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_alu_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_95_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_96_branch_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_95_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_96_mem_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_95_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_97_pc = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_pc :
    _io_o_issue_packs_0_T_96_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_97_inst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_inst :
    _io_o_issue_packs_0_T_96_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_func_code = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_func_code :
    _io_o_issue_packs_0_T_96_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_branch_predict_pack_valid = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_96_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_branch_predict_pack_target = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_96_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_97_branch_predict_pack_branch_type = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_96_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_branch_predict_pack_select = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_96_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_branch_predict_pack_taken = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_96_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_phy_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_96_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_stale_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_96_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_arch_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_96_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_97_inst_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_96_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_regWen = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_regWen :
    _io_o_issue_packs_0_T_96_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_src1_valid = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_96_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_phy_rs1 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_96_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_arch_rs1 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_96_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_src2_valid = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_96_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_phy_rs2 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_96_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_arch_rs2 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_96_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_rob_idx = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_96_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_imm = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_imm :
    _io_o_issue_packs_0_T_96_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_src1_value = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_96_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_src2_value = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_96_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_97_op1_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_96_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_97_op2_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_96_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_alu_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_96_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_97_branch_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_96_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_97_mem_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_96_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_98_pc = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_pc :
    _io_o_issue_packs_0_T_97_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_98_inst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_inst :
    _io_o_issue_packs_0_T_97_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_func_code = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_func_code :
    _io_o_issue_packs_0_T_97_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_branch_predict_pack_valid = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_97_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_branch_predict_pack_target = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_97_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_98_branch_predict_pack_branch_type = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_97_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_branch_predict_pack_select = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_97_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_branch_predict_pack_taken = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_97_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_phy_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_97_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_stale_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_97_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_arch_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_97_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_98_inst_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_97_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_regWen = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_regWen :
    _io_o_issue_packs_0_T_97_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_src1_valid = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_97_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_phy_rs1 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_97_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_arch_rs1 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_97_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_src2_valid = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_97_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_phy_rs2 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_97_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_arch_rs2 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_97_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_rob_idx = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_97_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_imm = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_imm :
    _io_o_issue_packs_0_T_97_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_src1_value = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_97_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_src2_value = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_97_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_98_op1_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_97_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_98_op2_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_97_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_alu_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_97_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_98_branch_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_97_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_98_mem_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_97_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_99_pc = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_pc :
    _io_o_issue_packs_0_T_98_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_99_inst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_inst :
    _io_o_issue_packs_0_T_98_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_func_code = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_func_code :
    _io_o_issue_packs_0_T_98_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_branch_predict_pack_valid = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_98_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_branch_predict_pack_target = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_98_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_99_branch_predict_pack_branch_type = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_98_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_branch_predict_pack_select = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_98_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_branch_predict_pack_taken = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_98_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_phy_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_98_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_stale_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_98_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_arch_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_98_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_99_inst_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_98_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_regWen = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_regWen :
    _io_o_issue_packs_0_T_98_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_src1_valid = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_98_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_phy_rs1 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_98_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_arch_rs1 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_98_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_src2_valid = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_98_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_phy_rs2 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_98_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_arch_rs2 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_98_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_rob_idx = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_98_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_imm = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_imm :
    _io_o_issue_packs_0_T_98_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_src1_value = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_98_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_src2_value = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_98_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_99_op1_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_98_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_99_op2_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_98_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_alu_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_98_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_99_branch_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_98_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_99_mem_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_98_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_100_pc = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_pc :
    _io_o_issue_packs_0_T_99_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_100_inst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_inst :
    _io_o_issue_packs_0_T_99_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_func_code = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_func_code :
    _io_o_issue_packs_0_T_99_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_branch_predict_pack_valid = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_99_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_branch_predict_pack_target = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_99_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_100_branch_predict_pack_branch_type = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_99_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_branch_predict_pack_select = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_99_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_branch_predict_pack_taken = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_99_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_phy_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_99_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_stale_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_99_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_arch_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_99_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_100_inst_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_99_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_regWen = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_regWen :
    _io_o_issue_packs_0_T_99_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_src1_valid = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_99_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_phy_rs1 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_99_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_arch_rs1 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_99_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_src2_valid = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_99_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_phy_rs2 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_99_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_arch_rs2 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_99_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_rob_idx = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_99_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_imm = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_imm :
    _io_o_issue_packs_0_T_99_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_src1_value = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_99_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_src2_value = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_99_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_100_op1_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_99_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_100_op2_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_99_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_alu_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_99_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_100_branch_type = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_type : _io_o_issue_packs_0_T_99_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_100_mem_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_99_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_101_pc = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_pc :
    _io_o_issue_packs_0_T_100_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_101_inst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_inst :
    _io_o_issue_packs_0_T_100_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_func_code = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_func_code :
    _io_o_issue_packs_0_T_100_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_branch_predict_pack_valid = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_100_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_branch_predict_pack_target = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_100_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_101_branch_predict_pack_branch_type = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_100_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_branch_predict_pack_select = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_100_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_branch_predict_pack_taken = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_100_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_phy_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_100_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_stale_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_100_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_arch_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_100_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_101_inst_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_100_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_regWen = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_regWen :
    _io_o_issue_packs_0_T_100_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_src1_valid = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_100_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_phy_rs1 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_100_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_arch_rs1 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_100_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_src2_valid = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_100_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_phy_rs2 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_100_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_arch_rs2 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_100_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_rob_idx = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_100_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_imm = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_imm :
    _io_o_issue_packs_0_T_100_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_src1_value = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_100_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_src2_value = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_100_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_101_op1_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_100_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_101_op2_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_100_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_alu_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_100_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_101_branch_type = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_type : _io_o_issue_packs_0_T_100_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_101_mem_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_100_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_102_pc = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_pc :
    _io_o_issue_packs_0_T_101_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_102_inst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_inst :
    _io_o_issue_packs_0_T_101_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_func_code = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_func_code :
    _io_o_issue_packs_0_T_101_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_branch_predict_pack_valid = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_101_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_branch_predict_pack_target = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_101_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_102_branch_predict_pack_branch_type = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_101_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_branch_predict_pack_select = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_101_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_branch_predict_pack_taken = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_101_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_phy_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_101_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_stale_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_101_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_arch_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_101_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_102_inst_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_101_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_regWen = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_regWen :
    _io_o_issue_packs_0_T_101_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_src1_valid = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_101_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_phy_rs1 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_101_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_arch_rs1 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_101_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_src2_valid = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_101_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_phy_rs2 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_101_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_arch_rs2 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_101_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_rob_idx = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_101_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_imm = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_imm :
    _io_o_issue_packs_0_T_101_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_src1_value = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_101_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_src2_value = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_101_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_102_op1_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_101_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_102_op2_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_101_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_alu_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_101_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_102_branch_type = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_type : _io_o_issue_packs_0_T_101_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_102_mem_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_101_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_103_pc = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_pc :
    _io_o_issue_packs_0_T_102_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_103_inst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_inst :
    _io_o_issue_packs_0_T_102_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_func_code = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_func_code :
    _io_o_issue_packs_0_T_102_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_branch_predict_pack_valid = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_102_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_branch_predict_pack_target = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_102_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_103_branch_predict_pack_branch_type = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_102_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_branch_predict_pack_select = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_102_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_branch_predict_pack_taken = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_102_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_phy_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_102_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_stale_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_102_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_arch_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_102_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_103_inst_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_102_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_regWen = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_regWen :
    _io_o_issue_packs_0_T_102_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_src1_valid = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_102_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_phy_rs1 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_102_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_arch_rs1 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_102_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_src2_valid = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_102_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_phy_rs2 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_102_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_arch_rs2 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_102_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_rob_idx = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_102_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_imm = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_imm :
    _io_o_issue_packs_0_T_102_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_src1_value = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_102_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_src2_value = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_102_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_103_op1_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_102_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_103_op2_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_102_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_alu_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_102_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_103_branch_type = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_type : _io_o_issue_packs_0_T_102_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_103_mem_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_102_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_104_pc = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_pc :
    _io_o_issue_packs_0_T_103_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_104_inst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_inst :
    _io_o_issue_packs_0_T_103_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_func_code = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_func_code :
    _io_o_issue_packs_0_T_103_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_branch_predict_pack_valid = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_103_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_branch_predict_pack_target = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_103_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_104_branch_predict_pack_branch_type = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_103_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_branch_predict_pack_select = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_103_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_branch_predict_pack_taken = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_103_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_phy_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_103_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_stale_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_103_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_arch_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_103_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_104_inst_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_103_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_regWen = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_regWen :
    _io_o_issue_packs_0_T_103_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_src1_valid = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_103_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_phy_rs1 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_103_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_arch_rs1 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_103_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_src2_valid = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_103_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_phy_rs2 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_103_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_arch_rs2 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_103_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_rob_idx = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_103_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_imm = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_imm :
    _io_o_issue_packs_0_T_103_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_src1_value = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_103_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_src2_value = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_103_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_104_op1_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_103_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_104_op2_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_103_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_alu_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_103_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_104_branch_type = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_type : _io_o_issue_packs_0_T_103_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_104_mem_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_103_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_105_pc = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_pc :
    _io_o_issue_packs_0_T_104_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_105_inst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_inst :
    _io_o_issue_packs_0_T_104_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_func_code = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_func_code :
    _io_o_issue_packs_0_T_104_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_branch_predict_pack_valid = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_104_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_branch_predict_pack_target = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_104_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_105_branch_predict_pack_branch_type = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_104_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_branch_predict_pack_select = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_104_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_branch_predict_pack_taken = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_104_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_phy_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_104_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_stale_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_104_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_arch_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_104_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_105_inst_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_104_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_regWen = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_regWen :
    _io_o_issue_packs_0_T_104_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_src1_valid = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_104_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_phy_rs1 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_104_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_arch_rs1 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_104_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_src2_valid = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_104_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_phy_rs2 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_104_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_arch_rs2 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_104_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_rob_idx = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_104_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_imm = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_imm :
    _io_o_issue_packs_0_T_104_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_src1_value = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_104_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_src2_value = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_104_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_105_op1_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_104_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_105_op2_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_104_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_alu_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_104_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_105_branch_type = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_type : _io_o_issue_packs_0_T_104_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_105_mem_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_104_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_106_pc = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_pc :
    _io_o_issue_packs_0_T_105_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_106_inst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_inst :
    _io_o_issue_packs_0_T_105_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_func_code = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_func_code :
    _io_o_issue_packs_0_T_105_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_branch_predict_pack_valid = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_105_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_branch_predict_pack_target = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_105_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_106_branch_predict_pack_branch_type = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_105_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_branch_predict_pack_select = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_105_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_branch_predict_pack_taken = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_105_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_phy_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_105_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_stale_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_105_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_arch_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_105_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_106_inst_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_105_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_regWen = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_regWen :
    _io_o_issue_packs_0_T_105_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_src1_valid = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_105_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_phy_rs1 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_105_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_arch_rs1 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_105_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_src2_valid = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_105_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_phy_rs2 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_105_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_arch_rs2 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_105_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_rob_idx = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_105_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_imm = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_imm :
    _io_o_issue_packs_0_T_105_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_src1_value = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_105_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_src2_value = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_105_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_106_op1_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_105_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_106_op2_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_105_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_alu_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_105_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_106_branch_type = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_type : _io_o_issue_packs_0_T_105_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_106_mem_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_105_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_107_pc = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_pc :
    _io_o_issue_packs_0_T_106_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_107_inst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_inst :
    _io_o_issue_packs_0_T_106_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_func_code = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_func_code :
    _io_o_issue_packs_0_T_106_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_branch_predict_pack_valid = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_106_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_branch_predict_pack_target = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_106_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_107_branch_predict_pack_branch_type = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_106_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_branch_predict_pack_select = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_106_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_branch_predict_pack_taken = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_106_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_phy_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_106_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_stale_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_106_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_arch_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_106_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_107_inst_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_106_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_regWen = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_regWen :
    _io_o_issue_packs_0_T_106_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_src1_valid = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_106_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_phy_rs1 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_106_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_arch_rs1 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_106_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_src2_valid = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_106_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_phy_rs2 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_106_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_arch_rs2 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_106_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_rob_idx = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_106_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_imm = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_imm :
    _io_o_issue_packs_0_T_106_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_src1_value = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_106_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_src2_value = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_106_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_107_op1_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_106_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_107_op2_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_106_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_alu_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_106_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_107_branch_type = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_type : _io_o_issue_packs_0_T_106_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_107_mem_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_106_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_108_pc = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_pc :
    _io_o_issue_packs_0_T_107_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_108_inst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_inst :
    _io_o_issue_packs_0_T_107_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_func_code = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_func_code :
    _io_o_issue_packs_0_T_107_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_branch_predict_pack_valid = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_107_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_branch_predict_pack_target = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_107_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_108_branch_predict_pack_branch_type = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_107_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_branch_predict_pack_select = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_107_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_branch_predict_pack_taken = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_107_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_phy_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_107_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_stale_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_107_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_arch_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_107_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_108_inst_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_107_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_regWen = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_regWen :
    _io_o_issue_packs_0_T_107_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_src1_valid = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_107_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_phy_rs1 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_107_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_arch_rs1 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_107_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_src2_valid = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_107_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_phy_rs2 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_107_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_arch_rs2 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_107_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_rob_idx = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_107_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_imm = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_imm :
    _io_o_issue_packs_0_T_107_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_src1_value = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_107_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_src2_value = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_107_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_108_op1_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_107_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_108_op2_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_107_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_alu_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_107_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_108_branch_type = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_type : _io_o_issue_packs_0_T_107_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_108_mem_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_107_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_109_pc = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_pc :
    _io_o_issue_packs_0_T_108_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_109_inst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_inst :
    _io_o_issue_packs_0_T_108_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_func_code = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_func_code :
    _io_o_issue_packs_0_T_108_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_branch_predict_pack_valid = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_108_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_branch_predict_pack_target = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_108_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_109_branch_predict_pack_branch_type = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_108_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_branch_predict_pack_select = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_108_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_branch_predict_pack_taken = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_108_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_phy_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_108_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_stale_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_108_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_arch_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_108_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_109_inst_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_108_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_regWen = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_regWen :
    _io_o_issue_packs_0_T_108_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_src1_valid = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_108_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_phy_rs1 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_108_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_arch_rs1 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_108_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_src2_valid = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_108_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_phy_rs2 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_108_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_arch_rs2 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_108_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_rob_idx = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_108_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_imm = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_imm :
    _io_o_issue_packs_0_T_108_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_src1_value = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_108_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_src2_value = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_108_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_109_op1_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_108_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_109_op2_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_108_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_alu_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_108_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_109_branch_type = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_type : _io_o_issue_packs_0_T_108_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_109_mem_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_108_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_110_pc = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_pc :
    _io_o_issue_packs_0_T_109_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_110_inst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_inst :
    _io_o_issue_packs_0_T_109_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_func_code = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_func_code :
    _io_o_issue_packs_0_T_109_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_branch_predict_pack_valid = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_109_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_branch_predict_pack_target = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_109_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_110_branch_predict_pack_branch_type = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_109_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_branch_predict_pack_select = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_109_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_branch_predict_pack_taken = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_109_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_phy_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_109_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_stale_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_109_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_arch_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_109_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_110_inst_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_109_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_regWen = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_regWen :
    _io_o_issue_packs_0_T_109_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_src1_valid = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_109_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_phy_rs1 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_109_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_arch_rs1 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_109_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_src2_valid = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_109_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_phy_rs2 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_109_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_arch_rs2 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_109_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_rob_idx = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_109_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_imm = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_imm :
    _io_o_issue_packs_0_T_109_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_src1_value = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_109_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_src2_value = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_109_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_110_op1_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_109_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_110_op2_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_109_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_alu_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_109_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_110_branch_type = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_type : _io_o_issue_packs_0_T_109_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_110_mem_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_109_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_111_pc = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_pc :
    _io_o_issue_packs_0_T_110_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_111_inst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_inst :
    _io_o_issue_packs_0_T_110_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_func_code = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_func_code :
    _io_o_issue_packs_0_T_110_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_branch_predict_pack_valid = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_110_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_branch_predict_pack_target = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_110_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_111_branch_predict_pack_branch_type = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_110_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_branch_predict_pack_select = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_110_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_branch_predict_pack_taken = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_110_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_phy_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_110_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_stale_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_110_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_arch_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_110_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_111_inst_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_110_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_regWen = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_regWen :
    _io_o_issue_packs_0_T_110_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_src1_valid = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_110_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_phy_rs1 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_110_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_arch_rs1 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_110_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_src2_valid = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_110_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_phy_rs2 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_110_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_arch_rs2 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_110_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_rob_idx = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_110_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_imm = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_imm :
    _io_o_issue_packs_0_T_110_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_src1_value = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_110_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_src2_value = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_110_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_111_op1_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_110_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_111_op2_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_110_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_alu_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_110_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_111_branch_type = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_type : _io_o_issue_packs_0_T_110_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_111_mem_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_110_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_112_pc = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_pc :
    _io_o_issue_packs_0_T_111_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_112_inst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_inst :
    _io_o_issue_packs_0_T_111_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_func_code = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_func_code :
    _io_o_issue_packs_0_T_111_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_branch_predict_pack_valid = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_111_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_branch_predict_pack_target = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_111_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_112_branch_predict_pack_branch_type = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_111_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_branch_predict_pack_select = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_111_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_branch_predict_pack_taken = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_111_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_phy_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_111_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_stale_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_111_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_arch_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_111_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_112_inst_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_111_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_regWen = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_regWen :
    _io_o_issue_packs_0_T_111_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_src1_valid = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_111_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_phy_rs1 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_111_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_arch_rs1 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_111_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_src2_valid = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_111_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_phy_rs2 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_111_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_arch_rs2 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_111_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_rob_idx = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_111_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_imm = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_imm :
    _io_o_issue_packs_0_T_111_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_src1_value = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_111_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_src2_value = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_111_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_112_op1_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_111_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_112_op2_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_111_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_alu_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_111_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_112_branch_type = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_type : _io_o_issue_packs_0_T_111_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_112_mem_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_111_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_113_pc = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_pc :
    _io_o_issue_packs_0_T_112_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_113_inst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_inst :
    _io_o_issue_packs_0_T_112_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_func_code = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_func_code :
    _io_o_issue_packs_0_T_112_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_branch_predict_pack_valid = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_112_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_branch_predict_pack_target = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_112_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_113_branch_predict_pack_branch_type = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_112_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_branch_predict_pack_select = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_112_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_branch_predict_pack_taken = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_112_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_phy_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_112_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_stale_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_112_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_arch_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_112_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_113_inst_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_112_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_regWen = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_regWen :
    _io_o_issue_packs_0_T_112_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_src1_valid = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_112_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_phy_rs1 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_112_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_arch_rs1 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_112_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_src2_valid = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_112_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_phy_rs2 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_112_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_arch_rs2 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_112_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_rob_idx = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_112_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_imm = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_imm :
    _io_o_issue_packs_0_T_112_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_src1_value = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_112_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_src2_value = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_112_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_113_op1_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_112_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_113_op2_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_112_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_alu_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_112_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_113_branch_type = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_type : _io_o_issue_packs_0_T_112_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_113_mem_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_112_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_114_pc = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_pc :
    _io_o_issue_packs_0_T_113_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_114_inst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_inst :
    _io_o_issue_packs_0_T_113_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_func_code = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_func_code :
    _io_o_issue_packs_0_T_113_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_branch_predict_pack_valid = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_113_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_branch_predict_pack_target = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_113_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_114_branch_predict_pack_branch_type = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_113_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_branch_predict_pack_select = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_113_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_branch_predict_pack_taken = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_113_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_phy_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_113_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_stale_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_113_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_arch_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_113_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_114_inst_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_113_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_regWen = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_regWen :
    _io_o_issue_packs_0_T_113_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_src1_valid = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_113_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_phy_rs1 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_113_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_arch_rs1 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_113_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_src2_valid = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_113_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_phy_rs2 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_113_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_arch_rs2 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_113_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_rob_idx = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_113_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_imm = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_imm :
    _io_o_issue_packs_0_T_113_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_src1_value = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_113_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_src2_value = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_113_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_114_op1_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_113_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_114_op2_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_113_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_alu_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_113_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_114_branch_type = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_type : _io_o_issue_packs_0_T_113_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_114_mem_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_113_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_115_pc = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_pc :
    _io_o_issue_packs_0_T_114_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_115_inst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_inst :
    _io_o_issue_packs_0_T_114_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_func_code = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_func_code :
    _io_o_issue_packs_0_T_114_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_branch_predict_pack_valid = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_114_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_branch_predict_pack_target = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_114_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_115_branch_predict_pack_branch_type = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_114_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_branch_predict_pack_select = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_114_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_branch_predict_pack_taken = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_114_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_phy_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_114_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_stale_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_114_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_arch_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_114_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_115_inst_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_114_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_regWen = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_regWen :
    _io_o_issue_packs_0_T_114_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_src1_valid = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_114_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_phy_rs1 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_114_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_arch_rs1 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_114_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_src2_valid = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_114_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_phy_rs2 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_114_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_arch_rs2 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_114_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_rob_idx = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_114_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_imm = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_imm :
    _io_o_issue_packs_0_T_114_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_src1_value = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_114_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_src2_value = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_114_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_115_op1_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_114_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_115_op2_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_114_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_alu_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_114_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_115_branch_type = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_type : _io_o_issue_packs_0_T_114_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_115_mem_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_114_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_116_pc = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_pc :
    _io_o_issue_packs_0_T_115_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_116_inst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_inst :
    _io_o_issue_packs_0_T_115_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_func_code = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_func_code :
    _io_o_issue_packs_0_T_115_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_branch_predict_pack_valid = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_115_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_branch_predict_pack_target = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_115_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_116_branch_predict_pack_branch_type = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_115_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_branch_predict_pack_select = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_115_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_branch_predict_pack_taken = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_115_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_phy_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_115_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_stale_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_115_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_arch_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_115_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_116_inst_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_115_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_regWen = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_regWen :
    _io_o_issue_packs_0_T_115_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_src1_valid = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_115_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_phy_rs1 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_115_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_arch_rs1 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_115_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_src2_valid = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_115_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_phy_rs2 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_115_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_arch_rs2 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_115_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_rob_idx = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_115_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_imm = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_imm :
    _io_o_issue_packs_0_T_115_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_src1_value = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_115_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_src2_value = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_115_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_116_op1_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_115_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_116_op2_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_115_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_alu_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_115_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_116_branch_type = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_type : _io_o_issue_packs_0_T_115_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_116_mem_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_115_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_117_pc = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_pc :
    _io_o_issue_packs_0_T_116_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_117_inst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_inst :
    _io_o_issue_packs_0_T_116_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_func_code = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_func_code :
    _io_o_issue_packs_0_T_116_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_branch_predict_pack_valid = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_116_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_branch_predict_pack_target = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_116_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_117_branch_predict_pack_branch_type = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_116_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_branch_predict_pack_select = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_116_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_branch_predict_pack_taken = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_116_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_phy_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_116_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_stale_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_116_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_arch_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_116_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_117_inst_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_116_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_regWen = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_regWen :
    _io_o_issue_packs_0_T_116_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_src1_valid = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_116_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_phy_rs1 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_116_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_arch_rs1 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_116_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_src2_valid = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_116_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_phy_rs2 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_116_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_arch_rs2 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_116_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_rob_idx = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_116_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_imm = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_imm :
    _io_o_issue_packs_0_T_116_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_src1_value = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_116_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_src2_value = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_116_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_117_op1_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_116_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_117_op2_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_116_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_alu_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_116_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_117_branch_type = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_type : _io_o_issue_packs_0_T_116_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_117_mem_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_116_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_118_pc = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_pc :
    _io_o_issue_packs_0_T_117_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_118_inst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_inst :
    _io_o_issue_packs_0_T_117_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_func_code = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_func_code :
    _io_o_issue_packs_0_T_117_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_branch_predict_pack_valid = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_117_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_branch_predict_pack_target = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_117_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_118_branch_predict_pack_branch_type = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_117_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_branch_predict_pack_select = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_117_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_branch_predict_pack_taken = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_117_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_phy_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_117_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_stale_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_117_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_arch_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_117_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_118_inst_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_117_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_regWen = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_regWen :
    _io_o_issue_packs_0_T_117_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_src1_valid = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_117_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_phy_rs1 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_117_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_arch_rs1 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_117_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_src2_valid = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_117_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_phy_rs2 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_117_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_arch_rs2 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_117_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_rob_idx = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_117_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_imm = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_imm :
    _io_o_issue_packs_0_T_117_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_src1_value = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_117_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_src2_value = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_117_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_118_op1_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_117_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_118_op2_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_117_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_alu_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_117_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_118_branch_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_117_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_118_mem_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_117_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_119_pc = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_pc :
    _io_o_issue_packs_0_T_118_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_119_inst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_inst :
    _io_o_issue_packs_0_T_118_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_func_code = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_func_code :
    _io_o_issue_packs_0_T_118_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_branch_predict_pack_valid = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_118_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_branch_predict_pack_target = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_118_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_119_branch_predict_pack_branch_type = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_118_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_branch_predict_pack_select = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_118_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_branch_predict_pack_taken = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_118_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_phy_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_118_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_stale_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_118_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_arch_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_118_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_119_inst_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_118_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_regWen = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_regWen :
    _io_o_issue_packs_0_T_118_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_src1_valid = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_118_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_phy_rs1 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_118_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_arch_rs1 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_118_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_src2_valid = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_118_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_phy_rs2 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_118_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_arch_rs2 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_118_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_rob_idx = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_118_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_imm = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_imm :
    _io_o_issue_packs_0_T_118_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_src1_value = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_118_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_src2_value = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_118_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_119_op1_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_118_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_119_op2_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_118_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_alu_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_118_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_119_branch_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_118_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_119_mem_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_118_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_120_pc = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_pc :
    _io_o_issue_packs_0_T_119_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_120_inst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_inst :
    _io_o_issue_packs_0_T_119_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_func_code = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_func_code :
    _io_o_issue_packs_0_T_119_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_branch_predict_pack_valid = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_119_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_branch_predict_pack_target = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_119_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_120_branch_predict_pack_branch_type = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_119_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_branch_predict_pack_select = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_119_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_branch_predict_pack_taken = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_119_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_phy_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_119_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_stale_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_119_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_arch_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_119_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_120_inst_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_119_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_regWen = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_regWen :
    _io_o_issue_packs_0_T_119_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_src1_valid = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_119_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_phy_rs1 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_119_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_arch_rs1 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_119_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_src2_valid = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_119_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_phy_rs2 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_119_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_arch_rs2 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_119_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_rob_idx = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_119_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_imm = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_imm :
    _io_o_issue_packs_0_T_119_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_src1_value = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_119_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_src2_value = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_119_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_120_op1_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_119_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_120_op2_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_119_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_alu_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_119_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_120_branch_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_119_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_120_mem_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_119_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_121_pc = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_pc :
    _io_o_issue_packs_0_T_120_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_121_inst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_inst :
    _io_o_issue_packs_0_T_120_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_func_code = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_func_code :
    _io_o_issue_packs_0_T_120_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_branch_predict_pack_valid = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_120_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_branch_predict_pack_target = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_120_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_121_branch_predict_pack_branch_type = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_120_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_branch_predict_pack_select = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_120_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_branch_predict_pack_taken = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_120_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_phy_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_120_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_stale_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_120_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_arch_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_120_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_121_inst_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_120_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_regWen = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_regWen :
    _io_o_issue_packs_0_T_120_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_src1_valid = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_120_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_phy_rs1 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_120_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_arch_rs1 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_120_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_src2_valid = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_120_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_phy_rs2 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_120_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_arch_rs2 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_120_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_rob_idx = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_120_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_imm = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_imm :
    _io_o_issue_packs_0_T_120_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_src1_value = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_120_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_src2_value = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_120_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_121_op1_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_120_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_121_op2_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_120_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_alu_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_120_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_121_branch_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_120_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_121_mem_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_120_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_122_pc = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_pc :
    _io_o_issue_packs_0_T_121_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_122_inst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_inst :
    _io_o_issue_packs_0_T_121_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_func_code = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_func_code :
    _io_o_issue_packs_0_T_121_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_branch_predict_pack_valid = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_121_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_branch_predict_pack_target = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_121_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_122_branch_predict_pack_branch_type = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_121_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_branch_predict_pack_select = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_121_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_branch_predict_pack_taken = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_121_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_phy_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_121_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_stale_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_121_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_arch_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_121_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_122_inst_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_121_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_regWen = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_regWen :
    _io_o_issue_packs_0_T_121_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_src1_valid = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_121_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_phy_rs1 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_121_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_arch_rs1 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_121_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_src2_valid = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_121_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_phy_rs2 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_121_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_arch_rs2 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_121_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_rob_idx = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_121_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_imm = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_imm :
    _io_o_issue_packs_0_T_121_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_src1_value = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_121_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_src2_value = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_121_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_122_op1_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_121_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_122_op2_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_121_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_alu_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_121_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_122_branch_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_121_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_122_mem_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_121_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_123_pc = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_pc :
    _io_o_issue_packs_0_T_122_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_123_inst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_inst :
    _io_o_issue_packs_0_T_122_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_func_code = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_func_code :
    _io_o_issue_packs_0_T_122_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_branch_predict_pack_valid = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_122_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_branch_predict_pack_target = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_122_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_123_branch_predict_pack_branch_type = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_122_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_branch_predict_pack_select = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_122_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_branch_predict_pack_taken = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_122_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_phy_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_122_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_stale_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_122_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_arch_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_122_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_123_inst_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_122_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_regWen = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_regWen :
    _io_o_issue_packs_0_T_122_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_src1_valid = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_122_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_phy_rs1 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_122_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_arch_rs1 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_122_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_src2_valid = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_122_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_phy_rs2 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_122_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_arch_rs2 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_122_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_rob_idx = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_122_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_imm = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_imm :
    _io_o_issue_packs_0_T_122_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_src1_value = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_122_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_src2_value = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_122_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_123_op1_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_122_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_123_op2_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_122_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_alu_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_122_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_123_branch_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_122_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_123_mem_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_122_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_124_pc = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_pc :
    _io_o_issue_packs_0_T_123_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_124_inst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_inst :
    _io_o_issue_packs_0_T_123_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_func_code = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_func_code :
    _io_o_issue_packs_0_T_123_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_branch_predict_pack_valid = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_123_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_branch_predict_pack_target = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_123_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_124_branch_predict_pack_branch_type = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_123_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_branch_predict_pack_select = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_123_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_branch_predict_pack_taken = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_123_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_phy_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_123_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_stale_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_123_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_arch_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_123_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_124_inst_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_123_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_regWen = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_regWen :
    _io_o_issue_packs_0_T_123_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_src1_valid = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_123_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_phy_rs1 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_123_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_arch_rs1 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_123_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_src2_valid = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_123_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_phy_rs2 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_123_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_arch_rs2 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_123_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_rob_idx = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_123_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_imm = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_imm :
    _io_o_issue_packs_0_T_123_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_src1_value = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_123_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_src2_value = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_123_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_124_op1_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_123_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_124_op2_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_123_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_alu_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_123_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_124_branch_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_123_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_124_mem_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_123_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_125_pc = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_pc :
    _io_o_issue_packs_0_T_124_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_125_inst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_inst :
    _io_o_issue_packs_0_T_124_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_func_code = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_func_code :
    _io_o_issue_packs_0_T_124_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_branch_predict_pack_valid = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_124_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_branch_predict_pack_target = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_124_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_125_branch_predict_pack_branch_type = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_124_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_branch_predict_pack_select = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_124_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_branch_predict_pack_taken = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_124_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_phy_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_124_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_stale_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_124_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_arch_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_124_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_125_inst_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_124_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_regWen = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_regWen :
    _io_o_issue_packs_0_T_124_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_src1_valid = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_124_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_phy_rs1 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_124_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_arch_rs1 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_124_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_src2_valid = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_124_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_phy_rs2 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_124_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_arch_rs2 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_124_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_rob_idx = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_124_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_imm = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_imm :
    _io_o_issue_packs_0_T_124_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_src1_value = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_124_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_src2_value = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_124_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_125_op1_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_124_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_125_op2_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_124_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_alu_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_124_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_125_branch_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_124_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_125_mem_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_124_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_126_pc = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_pc :
    _io_o_issue_packs_0_T_125_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_126_inst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_inst :
    _io_o_issue_packs_0_T_125_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_func_code = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_func_code :
    _io_o_issue_packs_0_T_125_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_branch_predict_pack_valid = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_125_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_branch_predict_pack_target = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_125_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_126_branch_predict_pack_branch_type = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_125_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_branch_predict_pack_select = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_125_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_branch_predict_pack_taken = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_125_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_phy_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_125_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_stale_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_125_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_arch_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_125_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_126_inst_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_125_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_regWen = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_regWen :
    _io_o_issue_packs_0_T_125_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_src1_valid = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_125_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_phy_rs1 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_125_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_arch_rs1 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_125_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_src2_valid = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_125_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_phy_rs2 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_125_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_arch_rs2 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_125_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_rob_idx = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_125_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_imm = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_imm :
    _io_o_issue_packs_0_T_125_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_src1_value = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_125_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_src2_value = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_125_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_126_op1_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_125_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_126_op2_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_125_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_alu_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_125_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_126_branch_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_125_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_126_mem_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_125_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_64_pc = _issued_age_pack_issued_ages_1_T_63 ? reservation_station_63_io_o_uop_pc :
    reservation_station_0_io_o_uop_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_64_inst = _issued_age_pack_issued_ages_1_T_63 ? reservation_station_63_io_o_uop_inst
     : reservation_station_0_io_o_uop_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_func_code = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_func_code : reservation_station_0_io_o_uop_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_valid : reservation_station_0_io_o_uop_branch_predict_pack_valid
    ; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_target :
    reservation_station_0_io_o_uop_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_64_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_branch_type :
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_select :
    reservation_station_0_io_o_uop_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_taken : reservation_station_0_io_o_uop_branch_predict_pack_taken
    ; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_phy_dst = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_phy_dst : reservation_station_0_io_o_uop_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_stale_dst = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_stale_dst : reservation_station_0_io_o_uop_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_arch_dst = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_arch_dst : reservation_station_0_io_o_uop_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_64_inst_type = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_inst_type : reservation_station_0_io_o_uop_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_regWen = _issued_age_pack_issued_ages_1_T_63 ? reservation_station_63_io_o_uop_regWen
     : reservation_station_0_io_o_uop_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_src1_valid = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_src1_valid : reservation_station_0_io_o_uop_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_phy_rs1 = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_phy_rs1 : reservation_station_0_io_o_uop_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_arch_rs1 = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_arch_rs1 : reservation_station_0_io_o_uop_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_src2_valid = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_src2_valid : reservation_station_0_io_o_uop_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_phy_rs2 = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_phy_rs2 : reservation_station_0_io_o_uop_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_arch_rs2 = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_arch_rs2 : reservation_station_0_io_o_uop_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_rob_idx = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_rob_idx : reservation_station_0_io_o_uop_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_imm = _issued_age_pack_issued_ages_1_T_63 ? reservation_station_63_io_o_uop_imm
     : reservation_station_0_io_o_uop_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_src1_value = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_src1_value : reservation_station_0_io_o_uop_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_src2_value = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_src2_value : reservation_station_0_io_o_uop_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_64_op1_sel = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_op1_sel : reservation_station_0_io_o_uop_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_64_op2_sel = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_op2_sel : reservation_station_0_io_o_uop_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_alu_sel = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_alu_sel : reservation_station_0_io_o_uop_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_64_branch_type = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_branch_type : reservation_station_0_io_o_uop_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_64_mem_type = _issued_age_pack_issued_ages_1_T_63 ?
    reservation_station_63_io_o_uop_mem_type : reservation_station_0_io_o_uop_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_65_pc = _issued_age_pack_issued_ages_1_T_62 ? reservation_station_62_io_o_uop_pc :
    _io_o_issue_packs_1_T_64_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_65_inst = _issued_age_pack_issued_ages_1_T_62 ? reservation_station_62_io_o_uop_inst
     : _io_o_issue_packs_1_T_64_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_func_code = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_func_code : _io_o_issue_packs_1_T_64_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_64_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_64_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_65_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_64_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_64_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_64_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_phy_dst = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_phy_dst : _io_o_issue_packs_1_T_64_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_stale_dst = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_stale_dst : _io_o_issue_packs_1_T_64_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_arch_dst = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_arch_dst : _io_o_issue_packs_1_T_64_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_65_inst_type = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_inst_type : _io_o_issue_packs_1_T_64_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_regWen = _issued_age_pack_issued_ages_1_T_62 ? reservation_station_62_io_o_uop_regWen
     : _io_o_issue_packs_1_T_64_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_src1_valid = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_src1_valid : _io_o_issue_packs_1_T_64_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_phy_rs1 = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_64_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_arch_rs1 = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_64_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_src2_valid = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_src2_valid : _io_o_issue_packs_1_T_64_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_phy_rs2 = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_64_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_arch_rs2 = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_64_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_rob_idx = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_rob_idx : _io_o_issue_packs_1_T_64_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_imm = _issued_age_pack_issued_ages_1_T_62 ? reservation_station_62_io_o_uop_imm
     : _io_o_issue_packs_1_T_64_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_src1_value = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_src1_value : _io_o_issue_packs_1_T_64_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_src2_value = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_src2_value : _io_o_issue_packs_1_T_64_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_65_op1_sel = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_op1_sel : _io_o_issue_packs_1_T_64_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_65_op2_sel = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_op2_sel : _io_o_issue_packs_1_T_64_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_alu_sel = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_alu_sel : _io_o_issue_packs_1_T_64_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_65_branch_type = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_branch_type : _io_o_issue_packs_1_T_64_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_65_mem_type = _issued_age_pack_issued_ages_1_T_62 ?
    reservation_station_62_io_o_uop_mem_type : _io_o_issue_packs_1_T_64_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_66_pc = _issued_age_pack_issued_ages_1_T_61 ? reservation_station_61_io_o_uop_pc :
    _io_o_issue_packs_1_T_65_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_66_inst = _issued_age_pack_issued_ages_1_T_61 ? reservation_station_61_io_o_uop_inst
     : _io_o_issue_packs_1_T_65_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_func_code = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_func_code : _io_o_issue_packs_1_T_65_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_65_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_65_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_66_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_65_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_65_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_65_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_phy_dst = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_phy_dst : _io_o_issue_packs_1_T_65_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_stale_dst = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_stale_dst : _io_o_issue_packs_1_T_65_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_arch_dst = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_arch_dst : _io_o_issue_packs_1_T_65_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_66_inst_type = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_inst_type : _io_o_issue_packs_1_T_65_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_regWen = _issued_age_pack_issued_ages_1_T_61 ? reservation_station_61_io_o_uop_regWen
     : _io_o_issue_packs_1_T_65_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_src1_valid = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_src1_valid : _io_o_issue_packs_1_T_65_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_phy_rs1 = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_65_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_arch_rs1 = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_65_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_src2_valid = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_src2_valid : _io_o_issue_packs_1_T_65_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_phy_rs2 = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_65_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_arch_rs2 = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_65_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_rob_idx = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_rob_idx : _io_o_issue_packs_1_T_65_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_imm = _issued_age_pack_issued_ages_1_T_61 ? reservation_station_61_io_o_uop_imm
     : _io_o_issue_packs_1_T_65_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_src1_value = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_src1_value : _io_o_issue_packs_1_T_65_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_src2_value = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_src2_value : _io_o_issue_packs_1_T_65_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_66_op1_sel = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_op1_sel : _io_o_issue_packs_1_T_65_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_66_op2_sel = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_op2_sel : _io_o_issue_packs_1_T_65_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_alu_sel = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_alu_sel : _io_o_issue_packs_1_T_65_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_66_branch_type = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_branch_type : _io_o_issue_packs_1_T_65_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_66_mem_type = _issued_age_pack_issued_ages_1_T_61 ?
    reservation_station_61_io_o_uop_mem_type : _io_o_issue_packs_1_T_65_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_67_pc = _issued_age_pack_issued_ages_1_T_60 ? reservation_station_60_io_o_uop_pc :
    _io_o_issue_packs_1_T_66_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_67_inst = _issued_age_pack_issued_ages_1_T_60 ? reservation_station_60_io_o_uop_inst
     : _io_o_issue_packs_1_T_66_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_func_code = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_func_code : _io_o_issue_packs_1_T_66_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_66_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_66_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_67_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_66_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_66_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_66_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_phy_dst = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_phy_dst : _io_o_issue_packs_1_T_66_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_stale_dst = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_stale_dst : _io_o_issue_packs_1_T_66_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_arch_dst = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_arch_dst : _io_o_issue_packs_1_T_66_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_67_inst_type = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_inst_type : _io_o_issue_packs_1_T_66_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_regWen = _issued_age_pack_issued_ages_1_T_60 ? reservation_station_60_io_o_uop_regWen
     : _io_o_issue_packs_1_T_66_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_src1_valid = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_src1_valid : _io_o_issue_packs_1_T_66_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_phy_rs1 = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_66_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_arch_rs1 = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_66_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_src2_valid = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_src2_valid : _io_o_issue_packs_1_T_66_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_phy_rs2 = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_66_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_arch_rs2 = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_66_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_rob_idx = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_rob_idx : _io_o_issue_packs_1_T_66_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_imm = _issued_age_pack_issued_ages_1_T_60 ? reservation_station_60_io_o_uop_imm
     : _io_o_issue_packs_1_T_66_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_src1_value = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_src1_value : _io_o_issue_packs_1_T_66_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_src2_value = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_src2_value : _io_o_issue_packs_1_T_66_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_67_op1_sel = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_op1_sel : _io_o_issue_packs_1_T_66_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_67_op2_sel = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_op2_sel : _io_o_issue_packs_1_T_66_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_alu_sel = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_alu_sel : _io_o_issue_packs_1_T_66_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_67_branch_type = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_branch_type : _io_o_issue_packs_1_T_66_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_67_mem_type = _issued_age_pack_issued_ages_1_T_60 ?
    reservation_station_60_io_o_uop_mem_type : _io_o_issue_packs_1_T_66_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_68_pc = _issued_age_pack_issued_ages_1_T_59 ? reservation_station_59_io_o_uop_pc :
    _io_o_issue_packs_1_T_67_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_68_inst = _issued_age_pack_issued_ages_1_T_59 ? reservation_station_59_io_o_uop_inst
     : _io_o_issue_packs_1_T_67_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_func_code = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_func_code : _io_o_issue_packs_1_T_67_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_67_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_67_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_68_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_67_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_67_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_67_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_phy_dst = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_phy_dst : _io_o_issue_packs_1_T_67_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_stale_dst = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_stale_dst : _io_o_issue_packs_1_T_67_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_arch_dst = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_arch_dst : _io_o_issue_packs_1_T_67_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_68_inst_type = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_inst_type : _io_o_issue_packs_1_T_67_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_regWen = _issued_age_pack_issued_ages_1_T_59 ? reservation_station_59_io_o_uop_regWen
     : _io_o_issue_packs_1_T_67_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_src1_valid = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_src1_valid : _io_o_issue_packs_1_T_67_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_phy_rs1 = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_67_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_arch_rs1 = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_67_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_src2_valid = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_src2_valid : _io_o_issue_packs_1_T_67_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_phy_rs2 = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_67_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_arch_rs2 = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_67_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_rob_idx = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_rob_idx : _io_o_issue_packs_1_T_67_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_imm = _issued_age_pack_issued_ages_1_T_59 ? reservation_station_59_io_o_uop_imm
     : _io_o_issue_packs_1_T_67_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_src1_value = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_src1_value : _io_o_issue_packs_1_T_67_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_src2_value = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_src2_value : _io_o_issue_packs_1_T_67_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_68_op1_sel = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_op1_sel : _io_o_issue_packs_1_T_67_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_68_op2_sel = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_op2_sel : _io_o_issue_packs_1_T_67_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_alu_sel = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_alu_sel : _io_o_issue_packs_1_T_67_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_68_branch_type = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_branch_type : _io_o_issue_packs_1_T_67_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_68_mem_type = _issued_age_pack_issued_ages_1_T_59 ?
    reservation_station_59_io_o_uop_mem_type : _io_o_issue_packs_1_T_67_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_69_pc = _issued_age_pack_issued_ages_1_T_58 ? reservation_station_58_io_o_uop_pc :
    _io_o_issue_packs_1_T_68_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_69_inst = _issued_age_pack_issued_ages_1_T_58 ? reservation_station_58_io_o_uop_inst
     : _io_o_issue_packs_1_T_68_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_func_code = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_func_code : _io_o_issue_packs_1_T_68_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_68_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_68_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_69_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_68_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_68_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_68_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_phy_dst = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_phy_dst : _io_o_issue_packs_1_T_68_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_stale_dst = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_stale_dst : _io_o_issue_packs_1_T_68_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_arch_dst = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_arch_dst : _io_o_issue_packs_1_T_68_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_69_inst_type = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_inst_type : _io_o_issue_packs_1_T_68_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_regWen = _issued_age_pack_issued_ages_1_T_58 ? reservation_station_58_io_o_uop_regWen
     : _io_o_issue_packs_1_T_68_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_src1_valid = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_src1_valid : _io_o_issue_packs_1_T_68_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_phy_rs1 = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_68_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_arch_rs1 = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_68_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_src2_valid = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_src2_valid : _io_o_issue_packs_1_T_68_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_phy_rs2 = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_68_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_arch_rs2 = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_68_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_rob_idx = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_rob_idx : _io_o_issue_packs_1_T_68_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_imm = _issued_age_pack_issued_ages_1_T_58 ? reservation_station_58_io_o_uop_imm
     : _io_o_issue_packs_1_T_68_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_src1_value = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_src1_value : _io_o_issue_packs_1_T_68_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_src2_value = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_src2_value : _io_o_issue_packs_1_T_68_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_69_op1_sel = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_op1_sel : _io_o_issue_packs_1_T_68_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_69_op2_sel = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_op2_sel : _io_o_issue_packs_1_T_68_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_alu_sel = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_alu_sel : _io_o_issue_packs_1_T_68_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_69_branch_type = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_branch_type : _io_o_issue_packs_1_T_68_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_69_mem_type = _issued_age_pack_issued_ages_1_T_58 ?
    reservation_station_58_io_o_uop_mem_type : _io_o_issue_packs_1_T_68_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_70_pc = _issued_age_pack_issued_ages_1_T_57 ? reservation_station_57_io_o_uop_pc :
    _io_o_issue_packs_1_T_69_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_70_inst = _issued_age_pack_issued_ages_1_T_57 ? reservation_station_57_io_o_uop_inst
     : _io_o_issue_packs_1_T_69_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_func_code = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_func_code : _io_o_issue_packs_1_T_69_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_69_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_69_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_70_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_69_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_69_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_69_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_phy_dst = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_phy_dst : _io_o_issue_packs_1_T_69_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_stale_dst = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_stale_dst : _io_o_issue_packs_1_T_69_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_arch_dst = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_arch_dst : _io_o_issue_packs_1_T_69_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_70_inst_type = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_inst_type : _io_o_issue_packs_1_T_69_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_regWen = _issued_age_pack_issued_ages_1_T_57 ? reservation_station_57_io_o_uop_regWen
     : _io_o_issue_packs_1_T_69_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_src1_valid = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_src1_valid : _io_o_issue_packs_1_T_69_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_phy_rs1 = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_69_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_arch_rs1 = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_69_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_src2_valid = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_src2_valid : _io_o_issue_packs_1_T_69_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_phy_rs2 = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_69_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_arch_rs2 = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_69_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_rob_idx = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_rob_idx : _io_o_issue_packs_1_T_69_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_imm = _issued_age_pack_issued_ages_1_T_57 ? reservation_station_57_io_o_uop_imm
     : _io_o_issue_packs_1_T_69_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_src1_value = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_src1_value : _io_o_issue_packs_1_T_69_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_src2_value = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_src2_value : _io_o_issue_packs_1_T_69_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_70_op1_sel = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_op1_sel : _io_o_issue_packs_1_T_69_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_70_op2_sel = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_op2_sel : _io_o_issue_packs_1_T_69_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_alu_sel = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_alu_sel : _io_o_issue_packs_1_T_69_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_70_branch_type = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_branch_type : _io_o_issue_packs_1_T_69_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_70_mem_type = _issued_age_pack_issued_ages_1_T_57 ?
    reservation_station_57_io_o_uop_mem_type : _io_o_issue_packs_1_T_69_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_71_pc = _issued_age_pack_issued_ages_1_T_56 ? reservation_station_56_io_o_uop_pc :
    _io_o_issue_packs_1_T_70_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_71_inst = _issued_age_pack_issued_ages_1_T_56 ? reservation_station_56_io_o_uop_inst
     : _io_o_issue_packs_1_T_70_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_func_code = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_func_code : _io_o_issue_packs_1_T_70_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_70_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_70_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_71_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_70_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_70_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_70_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_phy_dst = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_phy_dst : _io_o_issue_packs_1_T_70_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_stale_dst = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_stale_dst : _io_o_issue_packs_1_T_70_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_arch_dst = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_arch_dst : _io_o_issue_packs_1_T_70_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_71_inst_type = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_inst_type : _io_o_issue_packs_1_T_70_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_regWen = _issued_age_pack_issued_ages_1_T_56 ? reservation_station_56_io_o_uop_regWen
     : _io_o_issue_packs_1_T_70_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_src1_valid = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_src1_valid : _io_o_issue_packs_1_T_70_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_phy_rs1 = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_70_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_arch_rs1 = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_70_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_src2_valid = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_src2_valid : _io_o_issue_packs_1_T_70_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_phy_rs2 = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_70_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_arch_rs2 = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_70_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_rob_idx = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_rob_idx : _io_o_issue_packs_1_T_70_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_imm = _issued_age_pack_issued_ages_1_T_56 ? reservation_station_56_io_o_uop_imm
     : _io_o_issue_packs_1_T_70_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_src1_value = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_src1_value : _io_o_issue_packs_1_T_70_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_src2_value = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_src2_value : _io_o_issue_packs_1_T_70_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_71_op1_sel = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_op1_sel : _io_o_issue_packs_1_T_70_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_71_op2_sel = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_op2_sel : _io_o_issue_packs_1_T_70_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_alu_sel = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_alu_sel : _io_o_issue_packs_1_T_70_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_71_branch_type = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_branch_type : _io_o_issue_packs_1_T_70_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_71_mem_type = _issued_age_pack_issued_ages_1_T_56 ?
    reservation_station_56_io_o_uop_mem_type : _io_o_issue_packs_1_T_70_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_72_pc = _issued_age_pack_issued_ages_1_T_55 ? reservation_station_55_io_o_uop_pc :
    _io_o_issue_packs_1_T_71_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_72_inst = _issued_age_pack_issued_ages_1_T_55 ? reservation_station_55_io_o_uop_inst
     : _io_o_issue_packs_1_T_71_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_func_code = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_func_code : _io_o_issue_packs_1_T_71_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_71_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_71_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_72_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_71_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_71_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_71_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_phy_dst = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_phy_dst : _io_o_issue_packs_1_T_71_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_stale_dst = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_stale_dst : _io_o_issue_packs_1_T_71_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_arch_dst = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_arch_dst : _io_o_issue_packs_1_T_71_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_72_inst_type = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_inst_type : _io_o_issue_packs_1_T_71_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_regWen = _issued_age_pack_issued_ages_1_T_55 ? reservation_station_55_io_o_uop_regWen
     : _io_o_issue_packs_1_T_71_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_src1_valid = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_src1_valid : _io_o_issue_packs_1_T_71_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_phy_rs1 = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_71_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_arch_rs1 = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_71_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_src2_valid = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_src2_valid : _io_o_issue_packs_1_T_71_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_phy_rs2 = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_71_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_arch_rs2 = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_71_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_rob_idx = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_rob_idx : _io_o_issue_packs_1_T_71_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_imm = _issued_age_pack_issued_ages_1_T_55 ? reservation_station_55_io_o_uop_imm
     : _io_o_issue_packs_1_T_71_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_src1_value = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_src1_value : _io_o_issue_packs_1_T_71_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_src2_value = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_src2_value : _io_o_issue_packs_1_T_71_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_72_op1_sel = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_op1_sel : _io_o_issue_packs_1_T_71_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_72_op2_sel = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_op2_sel : _io_o_issue_packs_1_T_71_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_alu_sel = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_alu_sel : _io_o_issue_packs_1_T_71_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_72_branch_type = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_branch_type : _io_o_issue_packs_1_T_71_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_72_mem_type = _issued_age_pack_issued_ages_1_T_55 ?
    reservation_station_55_io_o_uop_mem_type : _io_o_issue_packs_1_T_71_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_73_pc = _issued_age_pack_issued_ages_1_T_54 ? reservation_station_54_io_o_uop_pc :
    _io_o_issue_packs_1_T_72_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_73_inst = _issued_age_pack_issued_ages_1_T_54 ? reservation_station_54_io_o_uop_inst
     : _io_o_issue_packs_1_T_72_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_func_code = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_func_code : _io_o_issue_packs_1_T_72_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_72_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_72_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_73_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_72_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_72_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_72_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_phy_dst = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_phy_dst : _io_o_issue_packs_1_T_72_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_stale_dst = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_stale_dst : _io_o_issue_packs_1_T_72_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_arch_dst = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_arch_dst : _io_o_issue_packs_1_T_72_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_73_inst_type = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_inst_type : _io_o_issue_packs_1_T_72_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_regWen = _issued_age_pack_issued_ages_1_T_54 ? reservation_station_54_io_o_uop_regWen
     : _io_o_issue_packs_1_T_72_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_src1_valid = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_src1_valid : _io_o_issue_packs_1_T_72_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_phy_rs1 = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_72_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_arch_rs1 = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_72_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_src2_valid = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_src2_valid : _io_o_issue_packs_1_T_72_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_phy_rs2 = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_72_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_arch_rs2 = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_72_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_rob_idx = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_rob_idx : _io_o_issue_packs_1_T_72_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_imm = _issued_age_pack_issued_ages_1_T_54 ? reservation_station_54_io_o_uop_imm
     : _io_o_issue_packs_1_T_72_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_src1_value = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_src1_value : _io_o_issue_packs_1_T_72_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_src2_value = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_src2_value : _io_o_issue_packs_1_T_72_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_73_op1_sel = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_op1_sel : _io_o_issue_packs_1_T_72_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_73_op2_sel = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_op2_sel : _io_o_issue_packs_1_T_72_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_alu_sel = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_alu_sel : _io_o_issue_packs_1_T_72_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_73_branch_type = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_branch_type : _io_o_issue_packs_1_T_72_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_73_mem_type = _issued_age_pack_issued_ages_1_T_54 ?
    reservation_station_54_io_o_uop_mem_type : _io_o_issue_packs_1_T_72_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_74_pc = _issued_age_pack_issued_ages_1_T_53 ? reservation_station_53_io_o_uop_pc :
    _io_o_issue_packs_1_T_73_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_74_inst = _issued_age_pack_issued_ages_1_T_53 ? reservation_station_53_io_o_uop_inst
     : _io_o_issue_packs_1_T_73_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_func_code = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_func_code : _io_o_issue_packs_1_T_73_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_73_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_73_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_74_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_73_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_73_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_73_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_phy_dst = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_phy_dst : _io_o_issue_packs_1_T_73_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_stale_dst = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_stale_dst : _io_o_issue_packs_1_T_73_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_arch_dst = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_arch_dst : _io_o_issue_packs_1_T_73_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_74_inst_type = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_inst_type : _io_o_issue_packs_1_T_73_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_regWen = _issued_age_pack_issued_ages_1_T_53 ? reservation_station_53_io_o_uop_regWen
     : _io_o_issue_packs_1_T_73_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_src1_valid = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_src1_valid : _io_o_issue_packs_1_T_73_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_phy_rs1 = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_73_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_arch_rs1 = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_73_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_src2_valid = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_src2_valid : _io_o_issue_packs_1_T_73_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_phy_rs2 = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_73_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_arch_rs2 = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_73_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_rob_idx = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_rob_idx : _io_o_issue_packs_1_T_73_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_imm = _issued_age_pack_issued_ages_1_T_53 ? reservation_station_53_io_o_uop_imm
     : _io_o_issue_packs_1_T_73_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_src1_value = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_src1_value : _io_o_issue_packs_1_T_73_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_src2_value = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_src2_value : _io_o_issue_packs_1_T_73_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_74_op1_sel = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_op1_sel : _io_o_issue_packs_1_T_73_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_74_op2_sel = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_op2_sel : _io_o_issue_packs_1_T_73_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_alu_sel = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_alu_sel : _io_o_issue_packs_1_T_73_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_74_branch_type = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_branch_type : _io_o_issue_packs_1_T_73_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_74_mem_type = _issued_age_pack_issued_ages_1_T_53 ?
    reservation_station_53_io_o_uop_mem_type : _io_o_issue_packs_1_T_73_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_75_pc = _issued_age_pack_issued_ages_1_T_52 ? reservation_station_52_io_o_uop_pc :
    _io_o_issue_packs_1_T_74_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_75_inst = _issued_age_pack_issued_ages_1_T_52 ? reservation_station_52_io_o_uop_inst
     : _io_o_issue_packs_1_T_74_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_func_code = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_func_code : _io_o_issue_packs_1_T_74_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_74_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_74_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_75_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_74_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_74_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_74_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_phy_dst = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_phy_dst : _io_o_issue_packs_1_T_74_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_stale_dst = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_stale_dst : _io_o_issue_packs_1_T_74_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_arch_dst = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_arch_dst : _io_o_issue_packs_1_T_74_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_75_inst_type = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_inst_type : _io_o_issue_packs_1_T_74_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_regWen = _issued_age_pack_issued_ages_1_T_52 ? reservation_station_52_io_o_uop_regWen
     : _io_o_issue_packs_1_T_74_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_src1_valid = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_src1_valid : _io_o_issue_packs_1_T_74_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_phy_rs1 = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_74_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_arch_rs1 = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_74_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_src2_valid = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_src2_valid : _io_o_issue_packs_1_T_74_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_phy_rs2 = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_74_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_arch_rs2 = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_74_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_rob_idx = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_rob_idx : _io_o_issue_packs_1_T_74_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_imm = _issued_age_pack_issued_ages_1_T_52 ? reservation_station_52_io_o_uop_imm
     : _io_o_issue_packs_1_T_74_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_src1_value = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_src1_value : _io_o_issue_packs_1_T_74_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_src2_value = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_src2_value : _io_o_issue_packs_1_T_74_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_75_op1_sel = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_op1_sel : _io_o_issue_packs_1_T_74_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_75_op2_sel = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_op2_sel : _io_o_issue_packs_1_T_74_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_alu_sel = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_alu_sel : _io_o_issue_packs_1_T_74_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_75_branch_type = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_branch_type : _io_o_issue_packs_1_T_74_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_75_mem_type = _issued_age_pack_issued_ages_1_T_52 ?
    reservation_station_52_io_o_uop_mem_type : _io_o_issue_packs_1_T_74_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_76_pc = _issued_age_pack_issued_ages_1_T_51 ? reservation_station_51_io_o_uop_pc :
    _io_o_issue_packs_1_T_75_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_76_inst = _issued_age_pack_issued_ages_1_T_51 ? reservation_station_51_io_o_uop_inst
     : _io_o_issue_packs_1_T_75_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_func_code = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_func_code : _io_o_issue_packs_1_T_75_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_75_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_75_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_76_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_75_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_75_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_75_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_phy_dst = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_phy_dst : _io_o_issue_packs_1_T_75_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_stale_dst = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_stale_dst : _io_o_issue_packs_1_T_75_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_arch_dst = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_arch_dst : _io_o_issue_packs_1_T_75_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_76_inst_type = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_inst_type : _io_o_issue_packs_1_T_75_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_regWen = _issued_age_pack_issued_ages_1_T_51 ? reservation_station_51_io_o_uop_regWen
     : _io_o_issue_packs_1_T_75_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_src1_valid = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_src1_valid : _io_o_issue_packs_1_T_75_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_phy_rs1 = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_75_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_arch_rs1 = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_75_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_src2_valid = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_src2_valid : _io_o_issue_packs_1_T_75_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_phy_rs2 = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_75_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_arch_rs2 = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_75_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_rob_idx = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_rob_idx : _io_o_issue_packs_1_T_75_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_imm = _issued_age_pack_issued_ages_1_T_51 ? reservation_station_51_io_o_uop_imm
     : _io_o_issue_packs_1_T_75_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_src1_value = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_src1_value : _io_o_issue_packs_1_T_75_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_src2_value = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_src2_value : _io_o_issue_packs_1_T_75_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_76_op1_sel = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_op1_sel : _io_o_issue_packs_1_T_75_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_76_op2_sel = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_op2_sel : _io_o_issue_packs_1_T_75_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_alu_sel = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_alu_sel : _io_o_issue_packs_1_T_75_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_76_branch_type = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_branch_type : _io_o_issue_packs_1_T_75_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_76_mem_type = _issued_age_pack_issued_ages_1_T_51 ?
    reservation_station_51_io_o_uop_mem_type : _io_o_issue_packs_1_T_75_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_77_pc = _issued_age_pack_issued_ages_1_T_50 ? reservation_station_50_io_o_uop_pc :
    _io_o_issue_packs_1_T_76_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_77_inst = _issued_age_pack_issued_ages_1_T_50 ? reservation_station_50_io_o_uop_inst
     : _io_o_issue_packs_1_T_76_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_func_code = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_func_code : _io_o_issue_packs_1_T_76_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_76_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_76_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_77_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_76_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_76_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_76_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_phy_dst = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_phy_dst : _io_o_issue_packs_1_T_76_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_stale_dst = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_stale_dst : _io_o_issue_packs_1_T_76_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_arch_dst = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_arch_dst : _io_o_issue_packs_1_T_76_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_77_inst_type = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_inst_type : _io_o_issue_packs_1_T_76_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_regWen = _issued_age_pack_issued_ages_1_T_50 ? reservation_station_50_io_o_uop_regWen
     : _io_o_issue_packs_1_T_76_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_src1_valid = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_src1_valid : _io_o_issue_packs_1_T_76_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_phy_rs1 = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_76_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_arch_rs1 = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_76_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_src2_valid = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_src2_valid : _io_o_issue_packs_1_T_76_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_phy_rs2 = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_76_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_arch_rs2 = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_76_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_rob_idx = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_rob_idx : _io_o_issue_packs_1_T_76_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_imm = _issued_age_pack_issued_ages_1_T_50 ? reservation_station_50_io_o_uop_imm
     : _io_o_issue_packs_1_T_76_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_src1_value = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_src1_value : _io_o_issue_packs_1_T_76_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_src2_value = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_src2_value : _io_o_issue_packs_1_T_76_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_77_op1_sel = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_op1_sel : _io_o_issue_packs_1_T_76_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_77_op2_sel = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_op2_sel : _io_o_issue_packs_1_T_76_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_alu_sel = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_alu_sel : _io_o_issue_packs_1_T_76_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_77_branch_type = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_branch_type : _io_o_issue_packs_1_T_76_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_77_mem_type = _issued_age_pack_issued_ages_1_T_50 ?
    reservation_station_50_io_o_uop_mem_type : _io_o_issue_packs_1_T_76_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_78_pc = _issued_age_pack_issued_ages_1_T_49 ? reservation_station_49_io_o_uop_pc :
    _io_o_issue_packs_1_T_77_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_78_inst = _issued_age_pack_issued_ages_1_T_49 ? reservation_station_49_io_o_uop_inst
     : _io_o_issue_packs_1_T_77_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_func_code = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_func_code : _io_o_issue_packs_1_T_77_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_77_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_77_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_78_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_77_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_77_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_77_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_phy_dst = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_phy_dst : _io_o_issue_packs_1_T_77_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_stale_dst = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_stale_dst : _io_o_issue_packs_1_T_77_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_arch_dst = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_arch_dst : _io_o_issue_packs_1_T_77_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_78_inst_type = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_inst_type : _io_o_issue_packs_1_T_77_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_regWen = _issued_age_pack_issued_ages_1_T_49 ? reservation_station_49_io_o_uop_regWen
     : _io_o_issue_packs_1_T_77_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_src1_valid = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_src1_valid : _io_o_issue_packs_1_T_77_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_phy_rs1 = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_77_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_arch_rs1 = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_77_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_src2_valid = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_src2_valid : _io_o_issue_packs_1_T_77_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_phy_rs2 = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_77_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_arch_rs2 = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_77_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_rob_idx = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_rob_idx : _io_o_issue_packs_1_T_77_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_imm = _issued_age_pack_issued_ages_1_T_49 ? reservation_station_49_io_o_uop_imm
     : _io_o_issue_packs_1_T_77_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_src1_value = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_src1_value : _io_o_issue_packs_1_T_77_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_src2_value = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_src2_value : _io_o_issue_packs_1_T_77_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_78_op1_sel = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_op1_sel : _io_o_issue_packs_1_T_77_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_78_op2_sel = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_op2_sel : _io_o_issue_packs_1_T_77_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_alu_sel = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_alu_sel : _io_o_issue_packs_1_T_77_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_78_branch_type = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_branch_type : _io_o_issue_packs_1_T_77_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_78_mem_type = _issued_age_pack_issued_ages_1_T_49 ?
    reservation_station_49_io_o_uop_mem_type : _io_o_issue_packs_1_T_77_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_79_pc = _issued_age_pack_issued_ages_1_T_48 ? reservation_station_48_io_o_uop_pc :
    _io_o_issue_packs_1_T_78_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_79_inst = _issued_age_pack_issued_ages_1_T_48 ? reservation_station_48_io_o_uop_inst
     : _io_o_issue_packs_1_T_78_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_func_code = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_func_code : _io_o_issue_packs_1_T_78_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_78_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_78_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_79_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_78_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_78_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_78_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_phy_dst = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_phy_dst : _io_o_issue_packs_1_T_78_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_stale_dst = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_stale_dst : _io_o_issue_packs_1_T_78_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_arch_dst = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_arch_dst : _io_o_issue_packs_1_T_78_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_79_inst_type = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_inst_type : _io_o_issue_packs_1_T_78_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_regWen = _issued_age_pack_issued_ages_1_T_48 ? reservation_station_48_io_o_uop_regWen
     : _io_o_issue_packs_1_T_78_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_src1_valid = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_src1_valid : _io_o_issue_packs_1_T_78_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_phy_rs1 = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_78_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_arch_rs1 = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_78_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_src2_valid = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_src2_valid : _io_o_issue_packs_1_T_78_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_phy_rs2 = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_78_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_arch_rs2 = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_78_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_rob_idx = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_rob_idx : _io_o_issue_packs_1_T_78_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_imm = _issued_age_pack_issued_ages_1_T_48 ? reservation_station_48_io_o_uop_imm
     : _io_o_issue_packs_1_T_78_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_src1_value = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_src1_value : _io_o_issue_packs_1_T_78_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_src2_value = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_src2_value : _io_o_issue_packs_1_T_78_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_79_op1_sel = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_op1_sel : _io_o_issue_packs_1_T_78_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_79_op2_sel = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_op2_sel : _io_o_issue_packs_1_T_78_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_alu_sel = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_alu_sel : _io_o_issue_packs_1_T_78_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_79_branch_type = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_branch_type : _io_o_issue_packs_1_T_78_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_79_mem_type = _issued_age_pack_issued_ages_1_T_48 ?
    reservation_station_48_io_o_uop_mem_type : _io_o_issue_packs_1_T_78_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_80_pc = _issued_age_pack_issued_ages_1_T_47 ? reservation_station_47_io_o_uop_pc :
    _io_o_issue_packs_1_T_79_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_80_inst = _issued_age_pack_issued_ages_1_T_47 ? reservation_station_47_io_o_uop_inst
     : _io_o_issue_packs_1_T_79_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_func_code = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_func_code : _io_o_issue_packs_1_T_79_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_79_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_79_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_80_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_79_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_79_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_79_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_phy_dst = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_phy_dst : _io_o_issue_packs_1_T_79_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_stale_dst = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_stale_dst : _io_o_issue_packs_1_T_79_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_arch_dst = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_arch_dst : _io_o_issue_packs_1_T_79_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_80_inst_type = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_inst_type : _io_o_issue_packs_1_T_79_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_regWen = _issued_age_pack_issued_ages_1_T_47 ? reservation_station_47_io_o_uop_regWen
     : _io_o_issue_packs_1_T_79_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_src1_valid = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_src1_valid : _io_o_issue_packs_1_T_79_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_phy_rs1 = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_79_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_arch_rs1 = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_79_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_src2_valid = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_src2_valid : _io_o_issue_packs_1_T_79_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_phy_rs2 = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_79_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_arch_rs2 = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_79_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_rob_idx = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_rob_idx : _io_o_issue_packs_1_T_79_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_imm = _issued_age_pack_issued_ages_1_T_47 ? reservation_station_47_io_o_uop_imm
     : _io_o_issue_packs_1_T_79_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_src1_value = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_src1_value : _io_o_issue_packs_1_T_79_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_src2_value = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_src2_value : _io_o_issue_packs_1_T_79_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_80_op1_sel = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_op1_sel : _io_o_issue_packs_1_T_79_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_80_op2_sel = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_op2_sel : _io_o_issue_packs_1_T_79_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_alu_sel = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_alu_sel : _io_o_issue_packs_1_T_79_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_80_branch_type = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_branch_type : _io_o_issue_packs_1_T_79_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_80_mem_type = _issued_age_pack_issued_ages_1_T_47 ?
    reservation_station_47_io_o_uop_mem_type : _io_o_issue_packs_1_T_79_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_81_pc = _issued_age_pack_issued_ages_1_T_46 ? reservation_station_46_io_o_uop_pc :
    _io_o_issue_packs_1_T_80_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_81_inst = _issued_age_pack_issued_ages_1_T_46 ? reservation_station_46_io_o_uop_inst
     : _io_o_issue_packs_1_T_80_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_func_code = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_func_code : _io_o_issue_packs_1_T_80_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_80_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_80_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_81_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_80_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_80_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_80_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_phy_dst = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_phy_dst : _io_o_issue_packs_1_T_80_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_stale_dst = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_stale_dst : _io_o_issue_packs_1_T_80_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_arch_dst = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_arch_dst : _io_o_issue_packs_1_T_80_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_81_inst_type = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_inst_type : _io_o_issue_packs_1_T_80_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_regWen = _issued_age_pack_issued_ages_1_T_46 ? reservation_station_46_io_o_uop_regWen
     : _io_o_issue_packs_1_T_80_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_src1_valid = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_src1_valid : _io_o_issue_packs_1_T_80_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_phy_rs1 = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_80_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_arch_rs1 = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_80_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_src2_valid = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_src2_valid : _io_o_issue_packs_1_T_80_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_phy_rs2 = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_80_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_arch_rs2 = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_80_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_rob_idx = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_rob_idx : _io_o_issue_packs_1_T_80_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_imm = _issued_age_pack_issued_ages_1_T_46 ? reservation_station_46_io_o_uop_imm
     : _io_o_issue_packs_1_T_80_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_src1_value = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_src1_value : _io_o_issue_packs_1_T_80_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_src2_value = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_src2_value : _io_o_issue_packs_1_T_80_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_81_op1_sel = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_op1_sel : _io_o_issue_packs_1_T_80_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_81_op2_sel = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_op2_sel : _io_o_issue_packs_1_T_80_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_alu_sel = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_alu_sel : _io_o_issue_packs_1_T_80_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_81_branch_type = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_branch_type : _io_o_issue_packs_1_T_80_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_81_mem_type = _issued_age_pack_issued_ages_1_T_46 ?
    reservation_station_46_io_o_uop_mem_type : _io_o_issue_packs_1_T_80_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_82_pc = _issued_age_pack_issued_ages_1_T_45 ? reservation_station_45_io_o_uop_pc :
    _io_o_issue_packs_1_T_81_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_82_inst = _issued_age_pack_issued_ages_1_T_45 ? reservation_station_45_io_o_uop_inst
     : _io_o_issue_packs_1_T_81_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_func_code = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_func_code : _io_o_issue_packs_1_T_81_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_81_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_81_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_82_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_81_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_81_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_81_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_phy_dst = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_phy_dst : _io_o_issue_packs_1_T_81_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_stale_dst = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_stale_dst : _io_o_issue_packs_1_T_81_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_arch_dst = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_arch_dst : _io_o_issue_packs_1_T_81_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_82_inst_type = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_inst_type : _io_o_issue_packs_1_T_81_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_regWen = _issued_age_pack_issued_ages_1_T_45 ? reservation_station_45_io_o_uop_regWen
     : _io_o_issue_packs_1_T_81_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_src1_valid = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_src1_valid : _io_o_issue_packs_1_T_81_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_phy_rs1 = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_81_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_arch_rs1 = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_81_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_src2_valid = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_src2_valid : _io_o_issue_packs_1_T_81_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_phy_rs2 = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_81_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_arch_rs2 = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_81_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_rob_idx = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_rob_idx : _io_o_issue_packs_1_T_81_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_imm = _issued_age_pack_issued_ages_1_T_45 ? reservation_station_45_io_o_uop_imm
     : _io_o_issue_packs_1_T_81_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_src1_value = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_src1_value : _io_o_issue_packs_1_T_81_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_src2_value = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_src2_value : _io_o_issue_packs_1_T_81_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_82_op1_sel = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_op1_sel : _io_o_issue_packs_1_T_81_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_82_op2_sel = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_op2_sel : _io_o_issue_packs_1_T_81_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_alu_sel = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_alu_sel : _io_o_issue_packs_1_T_81_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_82_branch_type = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_branch_type : _io_o_issue_packs_1_T_81_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_82_mem_type = _issued_age_pack_issued_ages_1_T_45 ?
    reservation_station_45_io_o_uop_mem_type : _io_o_issue_packs_1_T_81_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_83_pc = _issued_age_pack_issued_ages_1_T_44 ? reservation_station_44_io_o_uop_pc :
    _io_o_issue_packs_1_T_82_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_83_inst = _issued_age_pack_issued_ages_1_T_44 ? reservation_station_44_io_o_uop_inst
     : _io_o_issue_packs_1_T_82_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_func_code = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_func_code : _io_o_issue_packs_1_T_82_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_82_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_82_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_83_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_82_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_82_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_82_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_phy_dst = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_phy_dst : _io_o_issue_packs_1_T_82_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_stale_dst = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_stale_dst : _io_o_issue_packs_1_T_82_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_arch_dst = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_arch_dst : _io_o_issue_packs_1_T_82_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_83_inst_type = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_inst_type : _io_o_issue_packs_1_T_82_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_regWen = _issued_age_pack_issued_ages_1_T_44 ? reservation_station_44_io_o_uop_regWen
     : _io_o_issue_packs_1_T_82_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_src1_valid = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_src1_valid : _io_o_issue_packs_1_T_82_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_phy_rs1 = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_82_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_arch_rs1 = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_82_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_src2_valid = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_src2_valid : _io_o_issue_packs_1_T_82_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_phy_rs2 = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_82_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_arch_rs2 = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_82_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_rob_idx = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_rob_idx : _io_o_issue_packs_1_T_82_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_imm = _issued_age_pack_issued_ages_1_T_44 ? reservation_station_44_io_o_uop_imm
     : _io_o_issue_packs_1_T_82_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_src1_value = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_src1_value : _io_o_issue_packs_1_T_82_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_src2_value = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_src2_value : _io_o_issue_packs_1_T_82_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_83_op1_sel = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_op1_sel : _io_o_issue_packs_1_T_82_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_83_op2_sel = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_op2_sel : _io_o_issue_packs_1_T_82_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_alu_sel = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_alu_sel : _io_o_issue_packs_1_T_82_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_83_branch_type = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_branch_type : _io_o_issue_packs_1_T_82_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_83_mem_type = _issued_age_pack_issued_ages_1_T_44 ?
    reservation_station_44_io_o_uop_mem_type : _io_o_issue_packs_1_T_82_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_84_pc = _issued_age_pack_issued_ages_1_T_43 ? reservation_station_43_io_o_uop_pc :
    _io_o_issue_packs_1_T_83_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_84_inst = _issued_age_pack_issued_ages_1_T_43 ? reservation_station_43_io_o_uop_inst
     : _io_o_issue_packs_1_T_83_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_func_code = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_func_code : _io_o_issue_packs_1_T_83_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_83_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_83_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_84_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_83_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_83_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_83_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_phy_dst = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_phy_dst : _io_o_issue_packs_1_T_83_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_stale_dst = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_stale_dst : _io_o_issue_packs_1_T_83_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_arch_dst = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_arch_dst : _io_o_issue_packs_1_T_83_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_84_inst_type = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_inst_type : _io_o_issue_packs_1_T_83_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_regWen = _issued_age_pack_issued_ages_1_T_43 ? reservation_station_43_io_o_uop_regWen
     : _io_o_issue_packs_1_T_83_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_src1_valid = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_src1_valid : _io_o_issue_packs_1_T_83_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_phy_rs1 = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_83_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_arch_rs1 = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_83_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_src2_valid = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_src2_valid : _io_o_issue_packs_1_T_83_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_phy_rs2 = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_83_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_arch_rs2 = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_83_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_rob_idx = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_rob_idx : _io_o_issue_packs_1_T_83_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_imm = _issued_age_pack_issued_ages_1_T_43 ? reservation_station_43_io_o_uop_imm
     : _io_o_issue_packs_1_T_83_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_src1_value = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_src1_value : _io_o_issue_packs_1_T_83_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_src2_value = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_src2_value : _io_o_issue_packs_1_T_83_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_84_op1_sel = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_op1_sel : _io_o_issue_packs_1_T_83_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_84_op2_sel = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_op2_sel : _io_o_issue_packs_1_T_83_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_alu_sel = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_alu_sel : _io_o_issue_packs_1_T_83_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_84_branch_type = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_branch_type : _io_o_issue_packs_1_T_83_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_84_mem_type = _issued_age_pack_issued_ages_1_T_43 ?
    reservation_station_43_io_o_uop_mem_type : _io_o_issue_packs_1_T_83_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_85_pc = _issued_age_pack_issued_ages_1_T_42 ? reservation_station_42_io_o_uop_pc :
    _io_o_issue_packs_1_T_84_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_85_inst = _issued_age_pack_issued_ages_1_T_42 ? reservation_station_42_io_o_uop_inst
     : _io_o_issue_packs_1_T_84_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_func_code = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_func_code : _io_o_issue_packs_1_T_84_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_84_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_84_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_85_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_84_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_84_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_84_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_phy_dst = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_phy_dst : _io_o_issue_packs_1_T_84_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_stale_dst = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_stale_dst : _io_o_issue_packs_1_T_84_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_arch_dst = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_arch_dst : _io_o_issue_packs_1_T_84_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_85_inst_type = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_inst_type : _io_o_issue_packs_1_T_84_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_regWen = _issued_age_pack_issued_ages_1_T_42 ? reservation_station_42_io_o_uop_regWen
     : _io_o_issue_packs_1_T_84_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_src1_valid = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_src1_valid : _io_o_issue_packs_1_T_84_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_phy_rs1 = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_84_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_arch_rs1 = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_84_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_src2_valid = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_src2_valid : _io_o_issue_packs_1_T_84_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_phy_rs2 = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_84_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_arch_rs2 = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_84_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_rob_idx = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_rob_idx : _io_o_issue_packs_1_T_84_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_imm = _issued_age_pack_issued_ages_1_T_42 ? reservation_station_42_io_o_uop_imm
     : _io_o_issue_packs_1_T_84_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_src1_value = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_src1_value : _io_o_issue_packs_1_T_84_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_src2_value = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_src2_value : _io_o_issue_packs_1_T_84_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_85_op1_sel = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_op1_sel : _io_o_issue_packs_1_T_84_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_85_op2_sel = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_op2_sel : _io_o_issue_packs_1_T_84_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_alu_sel = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_alu_sel : _io_o_issue_packs_1_T_84_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_85_branch_type = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_branch_type : _io_o_issue_packs_1_T_84_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_85_mem_type = _issued_age_pack_issued_ages_1_T_42 ?
    reservation_station_42_io_o_uop_mem_type : _io_o_issue_packs_1_T_84_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_86_pc = _issued_age_pack_issued_ages_1_T_41 ? reservation_station_41_io_o_uop_pc :
    _io_o_issue_packs_1_T_85_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_86_inst = _issued_age_pack_issued_ages_1_T_41 ? reservation_station_41_io_o_uop_inst
     : _io_o_issue_packs_1_T_85_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_func_code = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_func_code : _io_o_issue_packs_1_T_85_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_85_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_85_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_86_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_85_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_85_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_85_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_phy_dst = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_phy_dst : _io_o_issue_packs_1_T_85_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_stale_dst = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_stale_dst : _io_o_issue_packs_1_T_85_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_arch_dst = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_arch_dst : _io_o_issue_packs_1_T_85_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_86_inst_type = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_inst_type : _io_o_issue_packs_1_T_85_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_regWen = _issued_age_pack_issued_ages_1_T_41 ? reservation_station_41_io_o_uop_regWen
     : _io_o_issue_packs_1_T_85_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_src1_valid = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_src1_valid : _io_o_issue_packs_1_T_85_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_phy_rs1 = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_85_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_arch_rs1 = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_85_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_src2_valid = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_src2_valid : _io_o_issue_packs_1_T_85_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_phy_rs2 = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_85_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_arch_rs2 = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_85_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_rob_idx = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_rob_idx : _io_o_issue_packs_1_T_85_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_imm = _issued_age_pack_issued_ages_1_T_41 ? reservation_station_41_io_o_uop_imm
     : _io_o_issue_packs_1_T_85_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_src1_value = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_src1_value : _io_o_issue_packs_1_T_85_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_src2_value = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_src2_value : _io_o_issue_packs_1_T_85_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_86_op1_sel = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_op1_sel : _io_o_issue_packs_1_T_85_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_86_op2_sel = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_op2_sel : _io_o_issue_packs_1_T_85_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_alu_sel = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_alu_sel : _io_o_issue_packs_1_T_85_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_86_branch_type = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_branch_type : _io_o_issue_packs_1_T_85_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_86_mem_type = _issued_age_pack_issued_ages_1_T_41 ?
    reservation_station_41_io_o_uop_mem_type : _io_o_issue_packs_1_T_85_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_87_pc = _issued_age_pack_issued_ages_1_T_40 ? reservation_station_40_io_o_uop_pc :
    _io_o_issue_packs_1_T_86_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_87_inst = _issued_age_pack_issued_ages_1_T_40 ? reservation_station_40_io_o_uop_inst
     : _io_o_issue_packs_1_T_86_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_func_code = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_func_code : _io_o_issue_packs_1_T_86_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_86_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_86_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_87_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_86_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_86_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_86_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_phy_dst = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_phy_dst : _io_o_issue_packs_1_T_86_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_stale_dst = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_stale_dst : _io_o_issue_packs_1_T_86_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_arch_dst = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_arch_dst : _io_o_issue_packs_1_T_86_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_87_inst_type = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_inst_type : _io_o_issue_packs_1_T_86_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_regWen = _issued_age_pack_issued_ages_1_T_40 ? reservation_station_40_io_o_uop_regWen
     : _io_o_issue_packs_1_T_86_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_src1_valid = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_src1_valid : _io_o_issue_packs_1_T_86_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_phy_rs1 = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_86_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_arch_rs1 = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_86_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_src2_valid = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_src2_valid : _io_o_issue_packs_1_T_86_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_phy_rs2 = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_86_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_arch_rs2 = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_86_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_rob_idx = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_rob_idx : _io_o_issue_packs_1_T_86_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_imm = _issued_age_pack_issued_ages_1_T_40 ? reservation_station_40_io_o_uop_imm
     : _io_o_issue_packs_1_T_86_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_src1_value = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_src1_value : _io_o_issue_packs_1_T_86_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_src2_value = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_src2_value : _io_o_issue_packs_1_T_86_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_87_op1_sel = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_op1_sel : _io_o_issue_packs_1_T_86_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_87_op2_sel = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_op2_sel : _io_o_issue_packs_1_T_86_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_alu_sel = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_alu_sel : _io_o_issue_packs_1_T_86_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_87_branch_type = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_branch_type : _io_o_issue_packs_1_T_86_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_87_mem_type = _issued_age_pack_issued_ages_1_T_40 ?
    reservation_station_40_io_o_uop_mem_type : _io_o_issue_packs_1_T_86_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_88_pc = _issued_age_pack_issued_ages_1_T_39 ? reservation_station_39_io_o_uop_pc :
    _io_o_issue_packs_1_T_87_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_88_inst = _issued_age_pack_issued_ages_1_T_39 ? reservation_station_39_io_o_uop_inst
     : _io_o_issue_packs_1_T_87_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_func_code = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_func_code : _io_o_issue_packs_1_T_87_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_87_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_87_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_88_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_87_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_87_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_87_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_phy_dst = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_phy_dst : _io_o_issue_packs_1_T_87_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_stale_dst = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_stale_dst : _io_o_issue_packs_1_T_87_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_arch_dst = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_arch_dst : _io_o_issue_packs_1_T_87_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_88_inst_type = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_inst_type : _io_o_issue_packs_1_T_87_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_regWen = _issued_age_pack_issued_ages_1_T_39 ? reservation_station_39_io_o_uop_regWen
     : _io_o_issue_packs_1_T_87_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_src1_valid = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_src1_valid : _io_o_issue_packs_1_T_87_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_phy_rs1 = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_87_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_arch_rs1 = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_87_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_src2_valid = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_src2_valid : _io_o_issue_packs_1_T_87_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_phy_rs2 = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_87_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_arch_rs2 = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_87_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_rob_idx = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_rob_idx : _io_o_issue_packs_1_T_87_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_imm = _issued_age_pack_issued_ages_1_T_39 ? reservation_station_39_io_o_uop_imm
     : _io_o_issue_packs_1_T_87_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_src1_value = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_src1_value : _io_o_issue_packs_1_T_87_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_src2_value = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_src2_value : _io_o_issue_packs_1_T_87_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_88_op1_sel = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_op1_sel : _io_o_issue_packs_1_T_87_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_88_op2_sel = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_op2_sel : _io_o_issue_packs_1_T_87_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_alu_sel = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_alu_sel : _io_o_issue_packs_1_T_87_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_88_branch_type = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_branch_type : _io_o_issue_packs_1_T_87_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_88_mem_type = _issued_age_pack_issued_ages_1_T_39 ?
    reservation_station_39_io_o_uop_mem_type : _io_o_issue_packs_1_T_87_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_89_pc = _issued_age_pack_issued_ages_1_T_38 ? reservation_station_38_io_o_uop_pc :
    _io_o_issue_packs_1_T_88_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_89_inst = _issued_age_pack_issued_ages_1_T_38 ? reservation_station_38_io_o_uop_inst
     : _io_o_issue_packs_1_T_88_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_func_code = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_func_code : _io_o_issue_packs_1_T_88_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_88_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_88_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_89_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_88_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_88_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_88_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_phy_dst = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_phy_dst : _io_o_issue_packs_1_T_88_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_stale_dst = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_stale_dst : _io_o_issue_packs_1_T_88_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_arch_dst = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_arch_dst : _io_o_issue_packs_1_T_88_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_89_inst_type = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_inst_type : _io_o_issue_packs_1_T_88_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_regWen = _issued_age_pack_issued_ages_1_T_38 ? reservation_station_38_io_o_uop_regWen
     : _io_o_issue_packs_1_T_88_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_src1_valid = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_src1_valid : _io_o_issue_packs_1_T_88_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_phy_rs1 = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_88_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_arch_rs1 = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_88_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_src2_valid = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_src2_valid : _io_o_issue_packs_1_T_88_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_phy_rs2 = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_88_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_arch_rs2 = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_88_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_rob_idx = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_rob_idx : _io_o_issue_packs_1_T_88_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_imm = _issued_age_pack_issued_ages_1_T_38 ? reservation_station_38_io_o_uop_imm
     : _io_o_issue_packs_1_T_88_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_src1_value = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_src1_value : _io_o_issue_packs_1_T_88_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_src2_value = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_src2_value : _io_o_issue_packs_1_T_88_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_89_op1_sel = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_op1_sel : _io_o_issue_packs_1_T_88_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_89_op2_sel = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_op2_sel : _io_o_issue_packs_1_T_88_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_alu_sel = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_alu_sel : _io_o_issue_packs_1_T_88_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_89_branch_type = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_branch_type : _io_o_issue_packs_1_T_88_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_89_mem_type = _issued_age_pack_issued_ages_1_T_38 ?
    reservation_station_38_io_o_uop_mem_type : _io_o_issue_packs_1_T_88_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_90_pc = _issued_age_pack_issued_ages_1_T_37 ? reservation_station_37_io_o_uop_pc :
    _io_o_issue_packs_1_T_89_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_90_inst = _issued_age_pack_issued_ages_1_T_37 ? reservation_station_37_io_o_uop_inst
     : _io_o_issue_packs_1_T_89_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_func_code = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_func_code : _io_o_issue_packs_1_T_89_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_89_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_89_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_90_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_89_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_89_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_89_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_phy_dst = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_phy_dst : _io_o_issue_packs_1_T_89_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_stale_dst = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_stale_dst : _io_o_issue_packs_1_T_89_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_arch_dst = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_arch_dst : _io_o_issue_packs_1_T_89_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_90_inst_type = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_inst_type : _io_o_issue_packs_1_T_89_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_regWen = _issued_age_pack_issued_ages_1_T_37 ? reservation_station_37_io_o_uop_regWen
     : _io_o_issue_packs_1_T_89_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_src1_valid = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_src1_valid : _io_o_issue_packs_1_T_89_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_phy_rs1 = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_89_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_arch_rs1 = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_89_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_src2_valid = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_src2_valid : _io_o_issue_packs_1_T_89_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_phy_rs2 = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_89_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_arch_rs2 = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_89_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_rob_idx = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_rob_idx : _io_o_issue_packs_1_T_89_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_imm = _issued_age_pack_issued_ages_1_T_37 ? reservation_station_37_io_o_uop_imm
     : _io_o_issue_packs_1_T_89_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_src1_value = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_src1_value : _io_o_issue_packs_1_T_89_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_src2_value = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_src2_value : _io_o_issue_packs_1_T_89_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_90_op1_sel = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_op1_sel : _io_o_issue_packs_1_T_89_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_90_op2_sel = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_op2_sel : _io_o_issue_packs_1_T_89_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_alu_sel = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_alu_sel : _io_o_issue_packs_1_T_89_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_90_branch_type = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_branch_type : _io_o_issue_packs_1_T_89_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_90_mem_type = _issued_age_pack_issued_ages_1_T_37 ?
    reservation_station_37_io_o_uop_mem_type : _io_o_issue_packs_1_T_89_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_91_pc = _issued_age_pack_issued_ages_1_T_36 ? reservation_station_36_io_o_uop_pc :
    _io_o_issue_packs_1_T_90_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_91_inst = _issued_age_pack_issued_ages_1_T_36 ? reservation_station_36_io_o_uop_inst
     : _io_o_issue_packs_1_T_90_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_func_code = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_func_code : _io_o_issue_packs_1_T_90_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_90_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_90_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_91_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_90_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_90_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_90_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_phy_dst = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_phy_dst : _io_o_issue_packs_1_T_90_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_stale_dst = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_stale_dst : _io_o_issue_packs_1_T_90_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_arch_dst = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_arch_dst : _io_o_issue_packs_1_T_90_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_91_inst_type = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_inst_type : _io_o_issue_packs_1_T_90_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_regWen = _issued_age_pack_issued_ages_1_T_36 ? reservation_station_36_io_o_uop_regWen
     : _io_o_issue_packs_1_T_90_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_src1_valid = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_src1_valid : _io_o_issue_packs_1_T_90_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_phy_rs1 = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_90_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_arch_rs1 = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_90_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_src2_valid = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_src2_valid : _io_o_issue_packs_1_T_90_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_phy_rs2 = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_90_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_arch_rs2 = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_90_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_rob_idx = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_rob_idx : _io_o_issue_packs_1_T_90_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_imm = _issued_age_pack_issued_ages_1_T_36 ? reservation_station_36_io_o_uop_imm
     : _io_o_issue_packs_1_T_90_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_src1_value = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_src1_value : _io_o_issue_packs_1_T_90_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_src2_value = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_src2_value : _io_o_issue_packs_1_T_90_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_91_op1_sel = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_op1_sel : _io_o_issue_packs_1_T_90_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_91_op2_sel = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_op2_sel : _io_o_issue_packs_1_T_90_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_alu_sel = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_alu_sel : _io_o_issue_packs_1_T_90_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_91_branch_type = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_branch_type : _io_o_issue_packs_1_T_90_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_91_mem_type = _issued_age_pack_issued_ages_1_T_36 ?
    reservation_station_36_io_o_uop_mem_type : _io_o_issue_packs_1_T_90_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_92_pc = _issued_age_pack_issued_ages_1_T_35 ? reservation_station_35_io_o_uop_pc :
    _io_o_issue_packs_1_T_91_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_92_inst = _issued_age_pack_issued_ages_1_T_35 ? reservation_station_35_io_o_uop_inst
     : _io_o_issue_packs_1_T_91_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_func_code = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_func_code : _io_o_issue_packs_1_T_91_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_91_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_91_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_92_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_91_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_91_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_91_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_phy_dst = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_phy_dst : _io_o_issue_packs_1_T_91_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_stale_dst = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_stale_dst : _io_o_issue_packs_1_T_91_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_arch_dst = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_arch_dst : _io_o_issue_packs_1_T_91_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_92_inst_type = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_inst_type : _io_o_issue_packs_1_T_91_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_regWen = _issued_age_pack_issued_ages_1_T_35 ? reservation_station_35_io_o_uop_regWen
     : _io_o_issue_packs_1_T_91_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_src1_valid = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_src1_valid : _io_o_issue_packs_1_T_91_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_phy_rs1 = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_91_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_arch_rs1 = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_91_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_src2_valid = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_src2_valid : _io_o_issue_packs_1_T_91_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_phy_rs2 = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_91_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_arch_rs2 = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_91_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_rob_idx = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_rob_idx : _io_o_issue_packs_1_T_91_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_imm = _issued_age_pack_issued_ages_1_T_35 ? reservation_station_35_io_o_uop_imm
     : _io_o_issue_packs_1_T_91_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_src1_value = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_src1_value : _io_o_issue_packs_1_T_91_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_src2_value = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_src2_value : _io_o_issue_packs_1_T_91_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_92_op1_sel = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_op1_sel : _io_o_issue_packs_1_T_91_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_92_op2_sel = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_op2_sel : _io_o_issue_packs_1_T_91_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_alu_sel = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_alu_sel : _io_o_issue_packs_1_T_91_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_92_branch_type = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_branch_type : _io_o_issue_packs_1_T_91_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_92_mem_type = _issued_age_pack_issued_ages_1_T_35 ?
    reservation_station_35_io_o_uop_mem_type : _io_o_issue_packs_1_T_91_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_93_pc = _issued_age_pack_issued_ages_1_T_34 ? reservation_station_34_io_o_uop_pc :
    _io_o_issue_packs_1_T_92_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_93_inst = _issued_age_pack_issued_ages_1_T_34 ? reservation_station_34_io_o_uop_inst
     : _io_o_issue_packs_1_T_92_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_func_code = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_func_code : _io_o_issue_packs_1_T_92_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_92_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_92_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_93_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_92_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_92_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_92_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_phy_dst = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_phy_dst : _io_o_issue_packs_1_T_92_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_stale_dst = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_stale_dst : _io_o_issue_packs_1_T_92_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_arch_dst = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_arch_dst : _io_o_issue_packs_1_T_92_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_93_inst_type = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_inst_type : _io_o_issue_packs_1_T_92_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_regWen = _issued_age_pack_issued_ages_1_T_34 ? reservation_station_34_io_o_uop_regWen
     : _io_o_issue_packs_1_T_92_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_src1_valid = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_src1_valid : _io_o_issue_packs_1_T_92_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_phy_rs1 = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_92_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_arch_rs1 = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_92_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_src2_valid = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_src2_valid : _io_o_issue_packs_1_T_92_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_phy_rs2 = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_92_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_arch_rs2 = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_92_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_rob_idx = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_rob_idx : _io_o_issue_packs_1_T_92_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_imm = _issued_age_pack_issued_ages_1_T_34 ? reservation_station_34_io_o_uop_imm
     : _io_o_issue_packs_1_T_92_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_src1_value = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_src1_value : _io_o_issue_packs_1_T_92_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_src2_value = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_src2_value : _io_o_issue_packs_1_T_92_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_93_op1_sel = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_op1_sel : _io_o_issue_packs_1_T_92_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_93_op2_sel = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_op2_sel : _io_o_issue_packs_1_T_92_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_alu_sel = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_alu_sel : _io_o_issue_packs_1_T_92_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_93_branch_type = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_branch_type : _io_o_issue_packs_1_T_92_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_93_mem_type = _issued_age_pack_issued_ages_1_T_34 ?
    reservation_station_34_io_o_uop_mem_type : _io_o_issue_packs_1_T_92_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_94_pc = _issued_age_pack_issued_ages_1_T_33 ? reservation_station_33_io_o_uop_pc :
    _io_o_issue_packs_1_T_93_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_94_inst = _issued_age_pack_issued_ages_1_T_33 ? reservation_station_33_io_o_uop_inst
     : _io_o_issue_packs_1_T_93_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_func_code = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_func_code : _io_o_issue_packs_1_T_93_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_93_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_93_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_94_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_93_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_93_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_93_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_phy_dst = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_phy_dst : _io_o_issue_packs_1_T_93_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_stale_dst = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_stale_dst : _io_o_issue_packs_1_T_93_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_arch_dst = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_arch_dst : _io_o_issue_packs_1_T_93_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_94_inst_type = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_inst_type : _io_o_issue_packs_1_T_93_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_regWen = _issued_age_pack_issued_ages_1_T_33 ? reservation_station_33_io_o_uop_regWen
     : _io_o_issue_packs_1_T_93_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_src1_valid = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_src1_valid : _io_o_issue_packs_1_T_93_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_phy_rs1 = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_93_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_arch_rs1 = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_93_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_src2_valid = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_src2_valid : _io_o_issue_packs_1_T_93_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_phy_rs2 = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_93_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_arch_rs2 = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_93_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_rob_idx = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_rob_idx : _io_o_issue_packs_1_T_93_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_imm = _issued_age_pack_issued_ages_1_T_33 ? reservation_station_33_io_o_uop_imm
     : _io_o_issue_packs_1_T_93_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_src1_value = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_src1_value : _io_o_issue_packs_1_T_93_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_src2_value = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_src2_value : _io_o_issue_packs_1_T_93_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_94_op1_sel = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_op1_sel : _io_o_issue_packs_1_T_93_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_94_op2_sel = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_op2_sel : _io_o_issue_packs_1_T_93_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_alu_sel = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_alu_sel : _io_o_issue_packs_1_T_93_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_94_branch_type = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_branch_type : _io_o_issue_packs_1_T_93_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_94_mem_type = _issued_age_pack_issued_ages_1_T_33 ?
    reservation_station_33_io_o_uop_mem_type : _io_o_issue_packs_1_T_93_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_95_pc = _issued_age_pack_issued_ages_1_T_32 ? reservation_station_32_io_o_uop_pc :
    _io_o_issue_packs_1_T_94_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_95_inst = _issued_age_pack_issued_ages_1_T_32 ? reservation_station_32_io_o_uop_inst
     : _io_o_issue_packs_1_T_94_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_func_code = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_func_code : _io_o_issue_packs_1_T_94_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_94_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_94_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_95_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_94_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_94_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_94_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_phy_dst = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_phy_dst : _io_o_issue_packs_1_T_94_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_stale_dst = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_stale_dst : _io_o_issue_packs_1_T_94_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_arch_dst = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_arch_dst : _io_o_issue_packs_1_T_94_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_95_inst_type = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_inst_type : _io_o_issue_packs_1_T_94_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_regWen = _issued_age_pack_issued_ages_1_T_32 ? reservation_station_32_io_o_uop_regWen
     : _io_o_issue_packs_1_T_94_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_src1_valid = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_src1_valid : _io_o_issue_packs_1_T_94_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_phy_rs1 = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_94_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_arch_rs1 = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_94_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_src2_valid = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_src2_valid : _io_o_issue_packs_1_T_94_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_phy_rs2 = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_94_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_arch_rs2 = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_94_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_rob_idx = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_rob_idx : _io_o_issue_packs_1_T_94_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_imm = _issued_age_pack_issued_ages_1_T_32 ? reservation_station_32_io_o_uop_imm
     : _io_o_issue_packs_1_T_94_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_src1_value = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_src1_value : _io_o_issue_packs_1_T_94_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_src2_value = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_src2_value : _io_o_issue_packs_1_T_94_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_95_op1_sel = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_op1_sel : _io_o_issue_packs_1_T_94_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_95_op2_sel = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_op2_sel : _io_o_issue_packs_1_T_94_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_alu_sel = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_alu_sel : _io_o_issue_packs_1_T_94_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_95_branch_type = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_branch_type : _io_o_issue_packs_1_T_94_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_95_mem_type = _issued_age_pack_issued_ages_1_T_32 ?
    reservation_station_32_io_o_uop_mem_type : _io_o_issue_packs_1_T_94_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_96_pc = _issued_age_pack_issued_ages_1_T_31 ? reservation_station_31_io_o_uop_pc :
    _io_o_issue_packs_1_T_95_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_96_inst = _issued_age_pack_issued_ages_1_T_31 ? reservation_station_31_io_o_uop_inst
     : _io_o_issue_packs_1_T_95_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_func_code = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_func_code : _io_o_issue_packs_1_T_95_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_95_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_95_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_96_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_95_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_95_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_95_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_phy_dst = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_phy_dst : _io_o_issue_packs_1_T_95_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_stale_dst = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_stale_dst : _io_o_issue_packs_1_T_95_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_arch_dst = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_arch_dst : _io_o_issue_packs_1_T_95_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_96_inst_type = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_inst_type : _io_o_issue_packs_1_T_95_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_regWen = _issued_age_pack_issued_ages_1_T_31 ? reservation_station_31_io_o_uop_regWen
     : _io_o_issue_packs_1_T_95_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_src1_valid = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_src1_valid : _io_o_issue_packs_1_T_95_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_phy_rs1 = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_95_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_arch_rs1 = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_95_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_src2_valid = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_src2_valid : _io_o_issue_packs_1_T_95_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_phy_rs2 = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_95_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_arch_rs2 = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_95_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_rob_idx = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_rob_idx : _io_o_issue_packs_1_T_95_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_imm = _issued_age_pack_issued_ages_1_T_31 ? reservation_station_31_io_o_uop_imm
     : _io_o_issue_packs_1_T_95_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_src1_value = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_src1_value : _io_o_issue_packs_1_T_95_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_src2_value = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_src2_value : _io_o_issue_packs_1_T_95_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_96_op1_sel = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_op1_sel : _io_o_issue_packs_1_T_95_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_96_op2_sel = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_op2_sel : _io_o_issue_packs_1_T_95_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_alu_sel = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_alu_sel : _io_o_issue_packs_1_T_95_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_96_branch_type = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_branch_type : _io_o_issue_packs_1_T_95_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_96_mem_type = _issued_age_pack_issued_ages_1_T_31 ?
    reservation_station_31_io_o_uop_mem_type : _io_o_issue_packs_1_T_95_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_97_pc = _issued_age_pack_issued_ages_1_T_30 ? reservation_station_30_io_o_uop_pc :
    _io_o_issue_packs_1_T_96_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_97_inst = _issued_age_pack_issued_ages_1_T_30 ? reservation_station_30_io_o_uop_inst
     : _io_o_issue_packs_1_T_96_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_func_code = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_func_code : _io_o_issue_packs_1_T_96_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_96_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_96_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_97_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_96_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_96_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_96_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_phy_dst = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_phy_dst : _io_o_issue_packs_1_T_96_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_stale_dst = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_stale_dst : _io_o_issue_packs_1_T_96_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_arch_dst = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_arch_dst : _io_o_issue_packs_1_T_96_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_97_inst_type = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_inst_type : _io_o_issue_packs_1_T_96_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_regWen = _issued_age_pack_issued_ages_1_T_30 ? reservation_station_30_io_o_uop_regWen
     : _io_o_issue_packs_1_T_96_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_src1_valid = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_src1_valid : _io_o_issue_packs_1_T_96_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_phy_rs1 = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_96_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_arch_rs1 = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_96_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_src2_valid = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_src2_valid : _io_o_issue_packs_1_T_96_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_phy_rs2 = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_96_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_arch_rs2 = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_96_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_rob_idx = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_rob_idx : _io_o_issue_packs_1_T_96_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_imm = _issued_age_pack_issued_ages_1_T_30 ? reservation_station_30_io_o_uop_imm
     : _io_o_issue_packs_1_T_96_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_src1_value = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_src1_value : _io_o_issue_packs_1_T_96_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_src2_value = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_src2_value : _io_o_issue_packs_1_T_96_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_97_op1_sel = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_op1_sel : _io_o_issue_packs_1_T_96_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_97_op2_sel = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_op2_sel : _io_o_issue_packs_1_T_96_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_alu_sel = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_alu_sel : _io_o_issue_packs_1_T_96_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_97_branch_type = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_branch_type : _io_o_issue_packs_1_T_96_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_97_mem_type = _issued_age_pack_issued_ages_1_T_30 ?
    reservation_station_30_io_o_uop_mem_type : _io_o_issue_packs_1_T_96_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_98_pc = _issued_age_pack_issued_ages_1_T_29 ? reservation_station_29_io_o_uop_pc :
    _io_o_issue_packs_1_T_97_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_98_inst = _issued_age_pack_issued_ages_1_T_29 ? reservation_station_29_io_o_uop_inst
     : _io_o_issue_packs_1_T_97_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_func_code = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_func_code : _io_o_issue_packs_1_T_97_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_97_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_97_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_98_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_97_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_97_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_97_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_phy_dst = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_phy_dst : _io_o_issue_packs_1_T_97_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_stale_dst = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_stale_dst : _io_o_issue_packs_1_T_97_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_arch_dst = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_arch_dst : _io_o_issue_packs_1_T_97_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_98_inst_type = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_inst_type : _io_o_issue_packs_1_T_97_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_regWen = _issued_age_pack_issued_ages_1_T_29 ? reservation_station_29_io_o_uop_regWen
     : _io_o_issue_packs_1_T_97_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_src1_valid = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_src1_valid : _io_o_issue_packs_1_T_97_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_phy_rs1 = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_97_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_arch_rs1 = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_97_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_src2_valid = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_src2_valid : _io_o_issue_packs_1_T_97_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_phy_rs2 = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_97_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_arch_rs2 = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_97_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_rob_idx = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_rob_idx : _io_o_issue_packs_1_T_97_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_imm = _issued_age_pack_issued_ages_1_T_29 ? reservation_station_29_io_o_uop_imm
     : _io_o_issue_packs_1_T_97_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_src1_value = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_src1_value : _io_o_issue_packs_1_T_97_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_src2_value = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_src2_value : _io_o_issue_packs_1_T_97_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_98_op1_sel = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_op1_sel : _io_o_issue_packs_1_T_97_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_98_op2_sel = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_op2_sel : _io_o_issue_packs_1_T_97_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_alu_sel = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_alu_sel : _io_o_issue_packs_1_T_97_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_98_branch_type = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_branch_type : _io_o_issue_packs_1_T_97_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_98_mem_type = _issued_age_pack_issued_ages_1_T_29 ?
    reservation_station_29_io_o_uop_mem_type : _io_o_issue_packs_1_T_97_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_99_pc = _issued_age_pack_issued_ages_1_T_28 ? reservation_station_28_io_o_uop_pc :
    _io_o_issue_packs_1_T_98_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_99_inst = _issued_age_pack_issued_ages_1_T_28 ? reservation_station_28_io_o_uop_inst
     : _io_o_issue_packs_1_T_98_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_func_code = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_func_code : _io_o_issue_packs_1_T_98_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_98_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_98_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_99_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_98_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_98_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_98_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_phy_dst = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_phy_dst : _io_o_issue_packs_1_T_98_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_stale_dst = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_stale_dst : _io_o_issue_packs_1_T_98_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_arch_dst = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_arch_dst : _io_o_issue_packs_1_T_98_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_99_inst_type = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_inst_type : _io_o_issue_packs_1_T_98_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_regWen = _issued_age_pack_issued_ages_1_T_28 ? reservation_station_28_io_o_uop_regWen
     : _io_o_issue_packs_1_T_98_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_src1_valid = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_src1_valid : _io_o_issue_packs_1_T_98_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_phy_rs1 = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_98_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_arch_rs1 = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_98_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_src2_valid = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_src2_valid : _io_o_issue_packs_1_T_98_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_phy_rs2 = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_98_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_arch_rs2 = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_98_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_rob_idx = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_rob_idx : _io_o_issue_packs_1_T_98_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_imm = _issued_age_pack_issued_ages_1_T_28 ? reservation_station_28_io_o_uop_imm
     : _io_o_issue_packs_1_T_98_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_src1_value = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_src1_value : _io_o_issue_packs_1_T_98_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_src2_value = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_src2_value : _io_o_issue_packs_1_T_98_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_99_op1_sel = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_op1_sel : _io_o_issue_packs_1_T_98_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_99_op2_sel = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_op2_sel : _io_o_issue_packs_1_T_98_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_alu_sel = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_alu_sel : _io_o_issue_packs_1_T_98_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_99_branch_type = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_branch_type : _io_o_issue_packs_1_T_98_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_99_mem_type = _issued_age_pack_issued_ages_1_T_28 ?
    reservation_station_28_io_o_uop_mem_type : _io_o_issue_packs_1_T_98_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_100_pc = _issued_age_pack_issued_ages_1_T_27 ? reservation_station_27_io_o_uop_pc :
    _io_o_issue_packs_1_T_99_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_100_inst = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_inst : _io_o_issue_packs_1_T_99_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_func_code = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_func_code : _io_o_issue_packs_1_T_99_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_99_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_99_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_100_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_99_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_99_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_99_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_phy_dst = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_phy_dst : _io_o_issue_packs_1_T_99_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_stale_dst = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_stale_dst : _io_o_issue_packs_1_T_99_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_arch_dst = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_arch_dst : _io_o_issue_packs_1_T_99_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_100_inst_type = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_inst_type : _io_o_issue_packs_1_T_99_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_regWen = _issued_age_pack_issued_ages_1_T_27 ? reservation_station_27_io_o_uop_regWen
     : _io_o_issue_packs_1_T_99_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_src1_valid = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_src1_valid : _io_o_issue_packs_1_T_99_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_phy_rs1 = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_99_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_arch_rs1 = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_99_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_src2_valid = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_src2_valid : _io_o_issue_packs_1_T_99_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_phy_rs2 = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_99_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_arch_rs2 = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_99_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_rob_idx = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_rob_idx : _io_o_issue_packs_1_T_99_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_imm = _issued_age_pack_issued_ages_1_T_27 ? reservation_station_27_io_o_uop_imm
     : _io_o_issue_packs_1_T_99_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_src1_value = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_src1_value : _io_o_issue_packs_1_T_99_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_src2_value = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_src2_value : _io_o_issue_packs_1_T_99_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_100_op1_sel = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_op1_sel : _io_o_issue_packs_1_T_99_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_100_op2_sel = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_op2_sel : _io_o_issue_packs_1_T_99_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_alu_sel = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_alu_sel : _io_o_issue_packs_1_T_99_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_100_branch_type = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_branch_type : _io_o_issue_packs_1_T_99_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_100_mem_type = _issued_age_pack_issued_ages_1_T_27 ?
    reservation_station_27_io_o_uop_mem_type : _io_o_issue_packs_1_T_99_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_101_pc = _issued_age_pack_issued_ages_1_T_26 ? reservation_station_26_io_o_uop_pc :
    _io_o_issue_packs_1_T_100_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_101_inst = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_inst : _io_o_issue_packs_1_T_100_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_func_code = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_func_code : _io_o_issue_packs_1_T_100_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_100_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_100_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_101_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_100_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_100_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_100_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_phy_dst = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_phy_dst : _io_o_issue_packs_1_T_100_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_stale_dst = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_stale_dst : _io_o_issue_packs_1_T_100_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_arch_dst = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_arch_dst : _io_o_issue_packs_1_T_100_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_101_inst_type = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_inst_type : _io_o_issue_packs_1_T_100_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_regWen = _issued_age_pack_issued_ages_1_T_26 ? reservation_station_26_io_o_uop_regWen
     : _io_o_issue_packs_1_T_100_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_src1_valid = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_src1_valid : _io_o_issue_packs_1_T_100_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_phy_rs1 = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_100_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_arch_rs1 = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_100_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_src2_valid = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_src2_valid : _io_o_issue_packs_1_T_100_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_phy_rs2 = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_100_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_arch_rs2 = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_100_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_rob_idx = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_rob_idx : _io_o_issue_packs_1_T_100_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_imm = _issued_age_pack_issued_ages_1_T_26 ? reservation_station_26_io_o_uop_imm
     : _io_o_issue_packs_1_T_100_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_src1_value = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_src1_value : _io_o_issue_packs_1_T_100_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_src2_value = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_src2_value : _io_o_issue_packs_1_T_100_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_101_op1_sel = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_op1_sel : _io_o_issue_packs_1_T_100_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_101_op2_sel = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_op2_sel : _io_o_issue_packs_1_T_100_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_alu_sel = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_alu_sel : _io_o_issue_packs_1_T_100_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_101_branch_type = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_branch_type : _io_o_issue_packs_1_T_100_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_101_mem_type = _issued_age_pack_issued_ages_1_T_26 ?
    reservation_station_26_io_o_uop_mem_type : _io_o_issue_packs_1_T_100_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_102_pc = _issued_age_pack_issued_ages_1_T_25 ? reservation_station_25_io_o_uop_pc :
    _io_o_issue_packs_1_T_101_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_102_inst = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_inst : _io_o_issue_packs_1_T_101_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_func_code = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_func_code : _io_o_issue_packs_1_T_101_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_101_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_101_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_102_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_101_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_101_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_101_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_phy_dst = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_phy_dst : _io_o_issue_packs_1_T_101_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_stale_dst = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_stale_dst : _io_o_issue_packs_1_T_101_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_arch_dst = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_arch_dst : _io_o_issue_packs_1_T_101_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_102_inst_type = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_inst_type : _io_o_issue_packs_1_T_101_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_regWen = _issued_age_pack_issued_ages_1_T_25 ? reservation_station_25_io_o_uop_regWen
     : _io_o_issue_packs_1_T_101_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_src1_valid = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_src1_valid : _io_o_issue_packs_1_T_101_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_phy_rs1 = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_101_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_arch_rs1 = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_101_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_src2_valid = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_src2_valid : _io_o_issue_packs_1_T_101_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_phy_rs2 = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_101_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_arch_rs2 = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_101_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_rob_idx = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_rob_idx : _io_o_issue_packs_1_T_101_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_imm = _issued_age_pack_issued_ages_1_T_25 ? reservation_station_25_io_o_uop_imm
     : _io_o_issue_packs_1_T_101_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_src1_value = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_src1_value : _io_o_issue_packs_1_T_101_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_src2_value = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_src2_value : _io_o_issue_packs_1_T_101_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_102_op1_sel = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_op1_sel : _io_o_issue_packs_1_T_101_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_102_op2_sel = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_op2_sel : _io_o_issue_packs_1_T_101_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_alu_sel = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_alu_sel : _io_o_issue_packs_1_T_101_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_102_branch_type = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_branch_type : _io_o_issue_packs_1_T_101_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_102_mem_type = _issued_age_pack_issued_ages_1_T_25 ?
    reservation_station_25_io_o_uop_mem_type : _io_o_issue_packs_1_T_101_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_103_pc = _issued_age_pack_issued_ages_1_T_24 ? reservation_station_24_io_o_uop_pc :
    _io_o_issue_packs_1_T_102_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_103_inst = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_inst : _io_o_issue_packs_1_T_102_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_func_code = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_func_code : _io_o_issue_packs_1_T_102_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_102_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_102_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_103_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_102_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_102_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_102_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_phy_dst = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_phy_dst : _io_o_issue_packs_1_T_102_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_stale_dst = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_stale_dst : _io_o_issue_packs_1_T_102_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_arch_dst = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_arch_dst : _io_o_issue_packs_1_T_102_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_103_inst_type = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_inst_type : _io_o_issue_packs_1_T_102_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_regWen = _issued_age_pack_issued_ages_1_T_24 ? reservation_station_24_io_o_uop_regWen
     : _io_o_issue_packs_1_T_102_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_src1_valid = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_src1_valid : _io_o_issue_packs_1_T_102_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_phy_rs1 = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_102_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_arch_rs1 = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_102_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_src2_valid = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_src2_valid : _io_o_issue_packs_1_T_102_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_phy_rs2 = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_102_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_arch_rs2 = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_102_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_rob_idx = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_rob_idx : _io_o_issue_packs_1_T_102_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_imm = _issued_age_pack_issued_ages_1_T_24 ? reservation_station_24_io_o_uop_imm
     : _io_o_issue_packs_1_T_102_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_src1_value = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_src1_value : _io_o_issue_packs_1_T_102_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_src2_value = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_src2_value : _io_o_issue_packs_1_T_102_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_103_op1_sel = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_op1_sel : _io_o_issue_packs_1_T_102_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_103_op2_sel = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_op2_sel : _io_o_issue_packs_1_T_102_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_alu_sel = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_alu_sel : _io_o_issue_packs_1_T_102_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_103_branch_type = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_branch_type : _io_o_issue_packs_1_T_102_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_103_mem_type = _issued_age_pack_issued_ages_1_T_24 ?
    reservation_station_24_io_o_uop_mem_type : _io_o_issue_packs_1_T_102_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_104_pc = _issued_age_pack_issued_ages_1_T_23 ? reservation_station_23_io_o_uop_pc :
    _io_o_issue_packs_1_T_103_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_104_inst = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_inst : _io_o_issue_packs_1_T_103_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_func_code = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_func_code : _io_o_issue_packs_1_T_103_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_103_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_103_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_104_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_103_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_103_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_103_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_phy_dst = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_phy_dst : _io_o_issue_packs_1_T_103_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_stale_dst = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_stale_dst : _io_o_issue_packs_1_T_103_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_arch_dst = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_arch_dst : _io_o_issue_packs_1_T_103_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_104_inst_type = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_inst_type : _io_o_issue_packs_1_T_103_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_regWen = _issued_age_pack_issued_ages_1_T_23 ? reservation_station_23_io_o_uop_regWen
     : _io_o_issue_packs_1_T_103_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_src1_valid = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_src1_valid : _io_o_issue_packs_1_T_103_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_phy_rs1 = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_103_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_arch_rs1 = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_103_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_src2_valid = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_src2_valid : _io_o_issue_packs_1_T_103_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_phy_rs2 = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_103_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_arch_rs2 = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_103_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_rob_idx = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_rob_idx : _io_o_issue_packs_1_T_103_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_imm = _issued_age_pack_issued_ages_1_T_23 ? reservation_station_23_io_o_uop_imm
     : _io_o_issue_packs_1_T_103_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_src1_value = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_src1_value : _io_o_issue_packs_1_T_103_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_src2_value = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_src2_value : _io_o_issue_packs_1_T_103_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_104_op1_sel = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_op1_sel : _io_o_issue_packs_1_T_103_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_104_op2_sel = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_op2_sel : _io_o_issue_packs_1_T_103_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_alu_sel = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_alu_sel : _io_o_issue_packs_1_T_103_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_104_branch_type = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_branch_type : _io_o_issue_packs_1_T_103_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_104_mem_type = _issued_age_pack_issued_ages_1_T_23 ?
    reservation_station_23_io_o_uop_mem_type : _io_o_issue_packs_1_T_103_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_105_pc = _issued_age_pack_issued_ages_1_T_22 ? reservation_station_22_io_o_uop_pc :
    _io_o_issue_packs_1_T_104_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_105_inst = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_inst : _io_o_issue_packs_1_T_104_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_func_code = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_func_code : _io_o_issue_packs_1_T_104_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_104_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_104_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_105_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_104_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_104_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_104_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_phy_dst = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_phy_dst : _io_o_issue_packs_1_T_104_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_stale_dst = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_stale_dst : _io_o_issue_packs_1_T_104_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_arch_dst = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_arch_dst : _io_o_issue_packs_1_T_104_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_105_inst_type = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_inst_type : _io_o_issue_packs_1_T_104_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_regWen = _issued_age_pack_issued_ages_1_T_22 ? reservation_station_22_io_o_uop_regWen
     : _io_o_issue_packs_1_T_104_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_src1_valid = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_src1_valid : _io_o_issue_packs_1_T_104_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_phy_rs1 = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_104_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_arch_rs1 = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_104_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_src2_valid = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_src2_valid : _io_o_issue_packs_1_T_104_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_phy_rs2 = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_104_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_arch_rs2 = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_104_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_rob_idx = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_rob_idx : _io_o_issue_packs_1_T_104_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_imm = _issued_age_pack_issued_ages_1_T_22 ? reservation_station_22_io_o_uop_imm
     : _io_o_issue_packs_1_T_104_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_src1_value = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_src1_value : _io_o_issue_packs_1_T_104_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_src2_value = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_src2_value : _io_o_issue_packs_1_T_104_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_105_op1_sel = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_op1_sel : _io_o_issue_packs_1_T_104_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_105_op2_sel = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_op2_sel : _io_o_issue_packs_1_T_104_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_alu_sel = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_alu_sel : _io_o_issue_packs_1_T_104_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_105_branch_type = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_branch_type : _io_o_issue_packs_1_T_104_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_105_mem_type = _issued_age_pack_issued_ages_1_T_22 ?
    reservation_station_22_io_o_uop_mem_type : _io_o_issue_packs_1_T_104_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_106_pc = _issued_age_pack_issued_ages_1_T_21 ? reservation_station_21_io_o_uop_pc :
    _io_o_issue_packs_1_T_105_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_106_inst = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_inst : _io_o_issue_packs_1_T_105_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_func_code = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_func_code : _io_o_issue_packs_1_T_105_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_105_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_105_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_106_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_105_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_105_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_105_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_phy_dst = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_phy_dst : _io_o_issue_packs_1_T_105_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_stale_dst = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_stale_dst : _io_o_issue_packs_1_T_105_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_arch_dst = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_arch_dst : _io_o_issue_packs_1_T_105_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_106_inst_type = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_inst_type : _io_o_issue_packs_1_T_105_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_regWen = _issued_age_pack_issued_ages_1_T_21 ? reservation_station_21_io_o_uop_regWen
     : _io_o_issue_packs_1_T_105_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_src1_valid = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_src1_valid : _io_o_issue_packs_1_T_105_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_phy_rs1 = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_105_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_arch_rs1 = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_105_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_src2_valid = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_src2_valid : _io_o_issue_packs_1_T_105_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_phy_rs2 = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_105_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_arch_rs2 = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_105_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_rob_idx = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_rob_idx : _io_o_issue_packs_1_T_105_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_imm = _issued_age_pack_issued_ages_1_T_21 ? reservation_station_21_io_o_uop_imm
     : _io_o_issue_packs_1_T_105_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_src1_value = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_src1_value : _io_o_issue_packs_1_T_105_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_src2_value = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_src2_value : _io_o_issue_packs_1_T_105_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_106_op1_sel = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_op1_sel : _io_o_issue_packs_1_T_105_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_106_op2_sel = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_op2_sel : _io_o_issue_packs_1_T_105_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_alu_sel = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_alu_sel : _io_o_issue_packs_1_T_105_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_106_branch_type = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_branch_type : _io_o_issue_packs_1_T_105_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_106_mem_type = _issued_age_pack_issued_ages_1_T_21 ?
    reservation_station_21_io_o_uop_mem_type : _io_o_issue_packs_1_T_105_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_107_pc = _issued_age_pack_issued_ages_1_T_20 ? reservation_station_20_io_o_uop_pc :
    _io_o_issue_packs_1_T_106_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_107_inst = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_inst : _io_o_issue_packs_1_T_106_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_func_code = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_func_code : _io_o_issue_packs_1_T_106_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_106_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_106_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_107_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_106_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_106_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_106_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_phy_dst = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_phy_dst : _io_o_issue_packs_1_T_106_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_stale_dst = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_stale_dst : _io_o_issue_packs_1_T_106_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_arch_dst = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_arch_dst : _io_o_issue_packs_1_T_106_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_107_inst_type = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_inst_type : _io_o_issue_packs_1_T_106_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_regWen = _issued_age_pack_issued_ages_1_T_20 ? reservation_station_20_io_o_uop_regWen
     : _io_o_issue_packs_1_T_106_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_src1_valid = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_src1_valid : _io_o_issue_packs_1_T_106_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_phy_rs1 = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_106_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_arch_rs1 = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_106_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_src2_valid = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_src2_valid : _io_o_issue_packs_1_T_106_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_phy_rs2 = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_106_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_arch_rs2 = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_106_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_rob_idx = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_rob_idx : _io_o_issue_packs_1_T_106_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_imm = _issued_age_pack_issued_ages_1_T_20 ? reservation_station_20_io_o_uop_imm
     : _io_o_issue_packs_1_T_106_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_src1_value = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_src1_value : _io_o_issue_packs_1_T_106_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_src2_value = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_src2_value : _io_o_issue_packs_1_T_106_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_107_op1_sel = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_op1_sel : _io_o_issue_packs_1_T_106_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_107_op2_sel = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_op2_sel : _io_o_issue_packs_1_T_106_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_alu_sel = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_alu_sel : _io_o_issue_packs_1_T_106_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_107_branch_type = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_branch_type : _io_o_issue_packs_1_T_106_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_107_mem_type = _issued_age_pack_issued_ages_1_T_20 ?
    reservation_station_20_io_o_uop_mem_type : _io_o_issue_packs_1_T_106_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_108_pc = _issued_age_pack_issued_ages_1_T_19 ? reservation_station_19_io_o_uop_pc :
    _io_o_issue_packs_1_T_107_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_108_inst = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_inst : _io_o_issue_packs_1_T_107_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_func_code = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_func_code : _io_o_issue_packs_1_T_107_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_107_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_107_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_108_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_107_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_107_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_107_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_phy_dst = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_phy_dst : _io_o_issue_packs_1_T_107_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_stale_dst = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_stale_dst : _io_o_issue_packs_1_T_107_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_arch_dst = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_arch_dst : _io_o_issue_packs_1_T_107_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_108_inst_type = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_inst_type : _io_o_issue_packs_1_T_107_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_regWen = _issued_age_pack_issued_ages_1_T_19 ? reservation_station_19_io_o_uop_regWen
     : _io_o_issue_packs_1_T_107_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_src1_valid = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_src1_valid : _io_o_issue_packs_1_T_107_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_phy_rs1 = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_107_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_arch_rs1 = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_107_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_src2_valid = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_src2_valid : _io_o_issue_packs_1_T_107_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_phy_rs2 = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_107_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_arch_rs2 = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_107_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_rob_idx = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_rob_idx : _io_o_issue_packs_1_T_107_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_imm = _issued_age_pack_issued_ages_1_T_19 ? reservation_station_19_io_o_uop_imm
     : _io_o_issue_packs_1_T_107_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_src1_value = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_src1_value : _io_o_issue_packs_1_T_107_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_src2_value = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_src2_value : _io_o_issue_packs_1_T_107_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_108_op1_sel = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_op1_sel : _io_o_issue_packs_1_T_107_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_108_op2_sel = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_op2_sel : _io_o_issue_packs_1_T_107_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_alu_sel = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_alu_sel : _io_o_issue_packs_1_T_107_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_108_branch_type = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_branch_type : _io_o_issue_packs_1_T_107_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_108_mem_type = _issued_age_pack_issued_ages_1_T_19 ?
    reservation_station_19_io_o_uop_mem_type : _io_o_issue_packs_1_T_107_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_109_pc = _issued_age_pack_issued_ages_1_T_18 ? reservation_station_18_io_o_uop_pc :
    _io_o_issue_packs_1_T_108_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_109_inst = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_inst : _io_o_issue_packs_1_T_108_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_func_code = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_func_code : _io_o_issue_packs_1_T_108_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_108_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_108_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_109_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_108_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_108_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_108_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_phy_dst = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_phy_dst : _io_o_issue_packs_1_T_108_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_stale_dst = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_stale_dst : _io_o_issue_packs_1_T_108_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_arch_dst = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_arch_dst : _io_o_issue_packs_1_T_108_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_109_inst_type = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_inst_type : _io_o_issue_packs_1_T_108_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_regWen = _issued_age_pack_issued_ages_1_T_18 ? reservation_station_18_io_o_uop_regWen
     : _io_o_issue_packs_1_T_108_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_src1_valid = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_src1_valid : _io_o_issue_packs_1_T_108_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_phy_rs1 = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_108_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_arch_rs1 = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_108_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_src2_valid = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_src2_valid : _io_o_issue_packs_1_T_108_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_phy_rs2 = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_108_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_arch_rs2 = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_108_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_rob_idx = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_rob_idx : _io_o_issue_packs_1_T_108_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_imm = _issued_age_pack_issued_ages_1_T_18 ? reservation_station_18_io_o_uop_imm
     : _io_o_issue_packs_1_T_108_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_src1_value = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_src1_value : _io_o_issue_packs_1_T_108_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_src2_value = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_src2_value : _io_o_issue_packs_1_T_108_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_109_op1_sel = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_op1_sel : _io_o_issue_packs_1_T_108_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_109_op2_sel = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_op2_sel : _io_o_issue_packs_1_T_108_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_alu_sel = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_alu_sel : _io_o_issue_packs_1_T_108_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_109_branch_type = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_branch_type : _io_o_issue_packs_1_T_108_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_109_mem_type = _issued_age_pack_issued_ages_1_T_18 ?
    reservation_station_18_io_o_uop_mem_type : _io_o_issue_packs_1_T_108_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_110_pc = _issued_age_pack_issued_ages_1_T_17 ? reservation_station_17_io_o_uop_pc :
    _io_o_issue_packs_1_T_109_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_110_inst = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_inst : _io_o_issue_packs_1_T_109_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_func_code = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_func_code : _io_o_issue_packs_1_T_109_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_109_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_109_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_110_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_109_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_109_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_109_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_phy_dst = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_phy_dst : _io_o_issue_packs_1_T_109_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_stale_dst = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_stale_dst : _io_o_issue_packs_1_T_109_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_arch_dst = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_arch_dst : _io_o_issue_packs_1_T_109_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_110_inst_type = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_inst_type : _io_o_issue_packs_1_T_109_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_regWen = _issued_age_pack_issued_ages_1_T_17 ? reservation_station_17_io_o_uop_regWen
     : _io_o_issue_packs_1_T_109_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_src1_valid = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_src1_valid : _io_o_issue_packs_1_T_109_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_phy_rs1 = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_109_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_arch_rs1 = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_109_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_src2_valid = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_src2_valid : _io_o_issue_packs_1_T_109_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_phy_rs2 = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_109_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_arch_rs2 = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_109_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_rob_idx = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_rob_idx : _io_o_issue_packs_1_T_109_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_imm = _issued_age_pack_issued_ages_1_T_17 ? reservation_station_17_io_o_uop_imm
     : _io_o_issue_packs_1_T_109_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_src1_value = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_src1_value : _io_o_issue_packs_1_T_109_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_src2_value = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_src2_value : _io_o_issue_packs_1_T_109_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_110_op1_sel = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_op1_sel : _io_o_issue_packs_1_T_109_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_110_op2_sel = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_op2_sel : _io_o_issue_packs_1_T_109_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_alu_sel = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_alu_sel : _io_o_issue_packs_1_T_109_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_110_branch_type = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_branch_type : _io_o_issue_packs_1_T_109_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_110_mem_type = _issued_age_pack_issued_ages_1_T_17 ?
    reservation_station_17_io_o_uop_mem_type : _io_o_issue_packs_1_T_109_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_111_pc = _issued_age_pack_issued_ages_1_T_16 ? reservation_station_16_io_o_uop_pc :
    _io_o_issue_packs_1_T_110_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_111_inst = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_inst : _io_o_issue_packs_1_T_110_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_func_code = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_func_code : _io_o_issue_packs_1_T_110_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_110_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_110_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_111_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_110_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_110_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_110_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_phy_dst = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_phy_dst : _io_o_issue_packs_1_T_110_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_stale_dst = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_stale_dst : _io_o_issue_packs_1_T_110_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_arch_dst = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_arch_dst : _io_o_issue_packs_1_T_110_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_111_inst_type = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_inst_type : _io_o_issue_packs_1_T_110_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_regWen = _issued_age_pack_issued_ages_1_T_16 ? reservation_station_16_io_o_uop_regWen
     : _io_o_issue_packs_1_T_110_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_src1_valid = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_src1_valid : _io_o_issue_packs_1_T_110_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_phy_rs1 = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_110_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_arch_rs1 = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_110_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_src2_valid = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_src2_valid : _io_o_issue_packs_1_T_110_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_phy_rs2 = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_110_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_arch_rs2 = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_110_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_rob_idx = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_rob_idx : _io_o_issue_packs_1_T_110_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_imm = _issued_age_pack_issued_ages_1_T_16 ? reservation_station_16_io_o_uop_imm
     : _io_o_issue_packs_1_T_110_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_src1_value = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_src1_value : _io_o_issue_packs_1_T_110_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_src2_value = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_src2_value : _io_o_issue_packs_1_T_110_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_111_op1_sel = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_op1_sel : _io_o_issue_packs_1_T_110_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_111_op2_sel = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_op2_sel : _io_o_issue_packs_1_T_110_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_alu_sel = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_alu_sel : _io_o_issue_packs_1_T_110_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_111_branch_type = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_branch_type : _io_o_issue_packs_1_T_110_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_111_mem_type = _issued_age_pack_issued_ages_1_T_16 ?
    reservation_station_16_io_o_uop_mem_type : _io_o_issue_packs_1_T_110_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_112_pc = _issued_age_pack_issued_ages_1_T_15 ? reservation_station_15_io_o_uop_pc :
    _io_o_issue_packs_1_T_111_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_112_inst = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_inst : _io_o_issue_packs_1_T_111_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_func_code = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_func_code : _io_o_issue_packs_1_T_111_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_111_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_111_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_112_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_111_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_111_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_111_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_phy_dst = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_phy_dst : _io_o_issue_packs_1_T_111_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_stale_dst = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_stale_dst : _io_o_issue_packs_1_T_111_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_arch_dst = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_arch_dst : _io_o_issue_packs_1_T_111_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_112_inst_type = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_inst_type : _io_o_issue_packs_1_T_111_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_regWen = _issued_age_pack_issued_ages_1_T_15 ? reservation_station_15_io_o_uop_regWen
     : _io_o_issue_packs_1_T_111_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_src1_valid = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_src1_valid : _io_o_issue_packs_1_T_111_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_phy_rs1 = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_111_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_arch_rs1 = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_111_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_src2_valid = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_src2_valid : _io_o_issue_packs_1_T_111_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_phy_rs2 = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_111_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_arch_rs2 = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_111_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_rob_idx = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_rob_idx : _io_o_issue_packs_1_T_111_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_imm = _issued_age_pack_issued_ages_1_T_15 ? reservation_station_15_io_o_uop_imm
     : _io_o_issue_packs_1_T_111_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_src1_value = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_src1_value : _io_o_issue_packs_1_T_111_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_src2_value = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_src2_value : _io_o_issue_packs_1_T_111_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_112_op1_sel = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_op1_sel : _io_o_issue_packs_1_T_111_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_112_op2_sel = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_op2_sel : _io_o_issue_packs_1_T_111_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_alu_sel = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_alu_sel : _io_o_issue_packs_1_T_111_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_112_branch_type = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_branch_type : _io_o_issue_packs_1_T_111_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_112_mem_type = _issued_age_pack_issued_ages_1_T_15 ?
    reservation_station_15_io_o_uop_mem_type : _io_o_issue_packs_1_T_111_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_113_pc = _issued_age_pack_issued_ages_1_T_14 ? reservation_station_14_io_o_uop_pc :
    _io_o_issue_packs_1_T_112_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_113_inst = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_inst : _io_o_issue_packs_1_T_112_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_func_code = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_func_code : _io_o_issue_packs_1_T_112_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_112_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_112_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_113_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_112_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_112_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_112_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_phy_dst = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_phy_dst : _io_o_issue_packs_1_T_112_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_stale_dst = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_stale_dst : _io_o_issue_packs_1_T_112_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_arch_dst = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_arch_dst : _io_o_issue_packs_1_T_112_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_113_inst_type = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_inst_type : _io_o_issue_packs_1_T_112_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_regWen = _issued_age_pack_issued_ages_1_T_14 ? reservation_station_14_io_o_uop_regWen
     : _io_o_issue_packs_1_T_112_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_src1_valid = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_src1_valid : _io_o_issue_packs_1_T_112_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_phy_rs1 = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_112_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_arch_rs1 = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_112_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_src2_valid = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_src2_valid : _io_o_issue_packs_1_T_112_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_phy_rs2 = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_112_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_arch_rs2 = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_112_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_rob_idx = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_rob_idx : _io_o_issue_packs_1_T_112_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_imm = _issued_age_pack_issued_ages_1_T_14 ? reservation_station_14_io_o_uop_imm
     : _io_o_issue_packs_1_T_112_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_src1_value = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_src1_value : _io_o_issue_packs_1_T_112_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_src2_value = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_src2_value : _io_o_issue_packs_1_T_112_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_113_op1_sel = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_op1_sel : _io_o_issue_packs_1_T_112_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_113_op2_sel = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_op2_sel : _io_o_issue_packs_1_T_112_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_alu_sel = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_alu_sel : _io_o_issue_packs_1_T_112_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_113_branch_type = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_branch_type : _io_o_issue_packs_1_T_112_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_113_mem_type = _issued_age_pack_issued_ages_1_T_14 ?
    reservation_station_14_io_o_uop_mem_type : _io_o_issue_packs_1_T_112_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_114_pc = _issued_age_pack_issued_ages_1_T_13 ? reservation_station_13_io_o_uop_pc :
    _io_o_issue_packs_1_T_113_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_114_inst = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_inst : _io_o_issue_packs_1_T_113_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_func_code = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_func_code : _io_o_issue_packs_1_T_113_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_113_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_113_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_114_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_113_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_113_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_113_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_phy_dst = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_phy_dst : _io_o_issue_packs_1_T_113_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_stale_dst = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_stale_dst : _io_o_issue_packs_1_T_113_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_arch_dst = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_arch_dst : _io_o_issue_packs_1_T_113_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_114_inst_type = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_inst_type : _io_o_issue_packs_1_T_113_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_regWen = _issued_age_pack_issued_ages_1_T_13 ? reservation_station_13_io_o_uop_regWen
     : _io_o_issue_packs_1_T_113_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_src1_valid = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_src1_valid : _io_o_issue_packs_1_T_113_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_phy_rs1 = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_113_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_arch_rs1 = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_113_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_src2_valid = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_src2_valid : _io_o_issue_packs_1_T_113_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_phy_rs2 = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_113_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_arch_rs2 = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_113_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_rob_idx = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_rob_idx : _io_o_issue_packs_1_T_113_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_imm = _issued_age_pack_issued_ages_1_T_13 ? reservation_station_13_io_o_uop_imm
     : _io_o_issue_packs_1_T_113_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_src1_value = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_src1_value : _io_o_issue_packs_1_T_113_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_src2_value = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_src2_value : _io_o_issue_packs_1_T_113_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_114_op1_sel = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_op1_sel : _io_o_issue_packs_1_T_113_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_114_op2_sel = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_op2_sel : _io_o_issue_packs_1_T_113_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_alu_sel = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_alu_sel : _io_o_issue_packs_1_T_113_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_114_branch_type = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_branch_type : _io_o_issue_packs_1_T_113_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_114_mem_type = _issued_age_pack_issued_ages_1_T_13 ?
    reservation_station_13_io_o_uop_mem_type : _io_o_issue_packs_1_T_113_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_115_pc = _issued_age_pack_issued_ages_1_T_12 ? reservation_station_12_io_o_uop_pc :
    _io_o_issue_packs_1_T_114_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_115_inst = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_inst : _io_o_issue_packs_1_T_114_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_func_code = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_func_code : _io_o_issue_packs_1_T_114_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_114_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_114_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_115_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_114_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_114_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_114_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_phy_dst = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_phy_dst : _io_o_issue_packs_1_T_114_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_stale_dst = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_stale_dst : _io_o_issue_packs_1_T_114_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_arch_dst = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_arch_dst : _io_o_issue_packs_1_T_114_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_115_inst_type = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_inst_type : _io_o_issue_packs_1_T_114_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_regWen = _issued_age_pack_issued_ages_1_T_12 ? reservation_station_12_io_o_uop_regWen
     : _io_o_issue_packs_1_T_114_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_src1_valid = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_src1_valid : _io_o_issue_packs_1_T_114_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_phy_rs1 = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_114_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_arch_rs1 = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_114_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_src2_valid = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_src2_valid : _io_o_issue_packs_1_T_114_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_phy_rs2 = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_114_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_arch_rs2 = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_114_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_rob_idx = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_rob_idx : _io_o_issue_packs_1_T_114_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_imm = _issued_age_pack_issued_ages_1_T_12 ? reservation_station_12_io_o_uop_imm
     : _io_o_issue_packs_1_T_114_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_src1_value = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_src1_value : _io_o_issue_packs_1_T_114_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_src2_value = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_src2_value : _io_o_issue_packs_1_T_114_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_115_op1_sel = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_op1_sel : _io_o_issue_packs_1_T_114_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_115_op2_sel = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_op2_sel : _io_o_issue_packs_1_T_114_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_alu_sel = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_alu_sel : _io_o_issue_packs_1_T_114_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_115_branch_type = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_branch_type : _io_o_issue_packs_1_T_114_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_115_mem_type = _issued_age_pack_issued_ages_1_T_12 ?
    reservation_station_12_io_o_uop_mem_type : _io_o_issue_packs_1_T_114_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_116_pc = _issued_age_pack_issued_ages_1_T_11 ? reservation_station_11_io_o_uop_pc :
    _io_o_issue_packs_1_T_115_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_116_inst = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_inst : _io_o_issue_packs_1_T_115_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_func_code = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_func_code : _io_o_issue_packs_1_T_115_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_115_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_115_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_116_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_115_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_115_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_115_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_phy_dst = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_phy_dst : _io_o_issue_packs_1_T_115_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_stale_dst = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_stale_dst : _io_o_issue_packs_1_T_115_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_arch_dst = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_arch_dst : _io_o_issue_packs_1_T_115_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_116_inst_type = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_inst_type : _io_o_issue_packs_1_T_115_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_regWen = _issued_age_pack_issued_ages_1_T_11 ? reservation_station_11_io_o_uop_regWen
     : _io_o_issue_packs_1_T_115_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_src1_valid = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_src1_valid : _io_o_issue_packs_1_T_115_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_phy_rs1 = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_115_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_arch_rs1 = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_115_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_src2_valid = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_src2_valid : _io_o_issue_packs_1_T_115_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_phy_rs2 = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_115_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_arch_rs2 = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_115_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_rob_idx = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_rob_idx : _io_o_issue_packs_1_T_115_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_imm = _issued_age_pack_issued_ages_1_T_11 ? reservation_station_11_io_o_uop_imm
     : _io_o_issue_packs_1_T_115_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_src1_value = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_src1_value : _io_o_issue_packs_1_T_115_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_src2_value = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_src2_value : _io_o_issue_packs_1_T_115_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_116_op1_sel = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_op1_sel : _io_o_issue_packs_1_T_115_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_116_op2_sel = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_op2_sel : _io_o_issue_packs_1_T_115_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_alu_sel = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_alu_sel : _io_o_issue_packs_1_T_115_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_116_branch_type = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_branch_type : _io_o_issue_packs_1_T_115_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_116_mem_type = _issued_age_pack_issued_ages_1_T_11 ?
    reservation_station_11_io_o_uop_mem_type : _io_o_issue_packs_1_T_115_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_117_pc = _issued_age_pack_issued_ages_1_T_10 ? reservation_station_10_io_o_uop_pc :
    _io_o_issue_packs_1_T_116_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_117_inst = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_inst : _io_o_issue_packs_1_T_116_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_func_code = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_func_code : _io_o_issue_packs_1_T_116_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_116_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_116_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_117_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_116_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_116_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_116_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_phy_dst = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_phy_dst : _io_o_issue_packs_1_T_116_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_stale_dst = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_stale_dst : _io_o_issue_packs_1_T_116_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_arch_dst = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_arch_dst : _io_o_issue_packs_1_T_116_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_117_inst_type = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_inst_type : _io_o_issue_packs_1_T_116_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_regWen = _issued_age_pack_issued_ages_1_T_10 ? reservation_station_10_io_o_uop_regWen
     : _io_o_issue_packs_1_T_116_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_src1_valid = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_src1_valid : _io_o_issue_packs_1_T_116_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_phy_rs1 = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_116_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_arch_rs1 = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_116_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_src2_valid = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_src2_valid : _io_o_issue_packs_1_T_116_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_phy_rs2 = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_116_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_arch_rs2 = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_116_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_rob_idx = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_rob_idx : _io_o_issue_packs_1_T_116_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_imm = _issued_age_pack_issued_ages_1_T_10 ? reservation_station_10_io_o_uop_imm
     : _io_o_issue_packs_1_T_116_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_src1_value = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_src1_value : _io_o_issue_packs_1_T_116_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_src2_value = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_src2_value : _io_o_issue_packs_1_T_116_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_117_op1_sel = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_op1_sel : _io_o_issue_packs_1_T_116_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_117_op2_sel = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_op2_sel : _io_o_issue_packs_1_T_116_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_alu_sel = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_alu_sel : _io_o_issue_packs_1_T_116_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_117_branch_type = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_branch_type : _io_o_issue_packs_1_T_116_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_117_mem_type = _issued_age_pack_issued_ages_1_T_10 ?
    reservation_station_10_io_o_uop_mem_type : _io_o_issue_packs_1_T_116_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_118_pc = _issued_age_pack_issued_ages_1_T_9 ? reservation_station_9_io_o_uop_pc :
    _io_o_issue_packs_1_T_117_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_118_inst = _issued_age_pack_issued_ages_1_T_9 ? reservation_station_9_io_o_uop_inst
     : _io_o_issue_packs_1_T_117_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_func_code = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_func_code : _io_o_issue_packs_1_T_117_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_117_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_117_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_118_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_117_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_117_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_117_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_phy_dst = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_phy_dst : _io_o_issue_packs_1_T_117_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_stale_dst = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_stale_dst : _io_o_issue_packs_1_T_117_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_arch_dst = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_arch_dst : _io_o_issue_packs_1_T_117_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_118_inst_type = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_inst_type : _io_o_issue_packs_1_T_117_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_regWen = _issued_age_pack_issued_ages_1_T_9 ? reservation_station_9_io_o_uop_regWen :
    _io_o_issue_packs_1_T_117_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_src1_valid = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_src1_valid : _io_o_issue_packs_1_T_117_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_phy_rs1 = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_117_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_arch_rs1 = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_117_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_src2_valid = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_src2_valid : _io_o_issue_packs_1_T_117_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_phy_rs2 = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_117_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_arch_rs2 = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_117_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_rob_idx = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_rob_idx : _io_o_issue_packs_1_T_117_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_imm = _issued_age_pack_issued_ages_1_T_9 ? reservation_station_9_io_o_uop_imm :
    _io_o_issue_packs_1_T_117_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_src1_value = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_src1_value : _io_o_issue_packs_1_T_117_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_src2_value = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_src2_value : _io_o_issue_packs_1_T_117_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_118_op1_sel = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_op1_sel : _io_o_issue_packs_1_T_117_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_118_op2_sel = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_op2_sel : _io_o_issue_packs_1_T_117_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_alu_sel = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_alu_sel : _io_o_issue_packs_1_T_117_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_118_branch_type = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_branch_type : _io_o_issue_packs_1_T_117_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_118_mem_type = _issued_age_pack_issued_ages_1_T_9 ?
    reservation_station_9_io_o_uop_mem_type : _io_o_issue_packs_1_T_117_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_119_pc = _issued_age_pack_issued_ages_1_T_8 ? reservation_station_8_io_o_uop_pc :
    _io_o_issue_packs_1_T_118_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_119_inst = _issued_age_pack_issued_ages_1_T_8 ? reservation_station_8_io_o_uop_inst
     : _io_o_issue_packs_1_T_118_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_func_code = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_func_code : _io_o_issue_packs_1_T_118_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_118_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_118_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_119_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_118_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_118_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_118_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_phy_dst = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_phy_dst : _io_o_issue_packs_1_T_118_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_stale_dst = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_stale_dst : _io_o_issue_packs_1_T_118_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_arch_dst = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_arch_dst : _io_o_issue_packs_1_T_118_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_119_inst_type = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_inst_type : _io_o_issue_packs_1_T_118_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_regWen = _issued_age_pack_issued_ages_1_T_8 ? reservation_station_8_io_o_uop_regWen :
    _io_o_issue_packs_1_T_118_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_src1_valid = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_src1_valid : _io_o_issue_packs_1_T_118_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_phy_rs1 = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_118_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_arch_rs1 = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_118_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_src2_valid = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_src2_valid : _io_o_issue_packs_1_T_118_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_phy_rs2 = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_118_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_arch_rs2 = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_118_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_rob_idx = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_rob_idx : _io_o_issue_packs_1_T_118_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_imm = _issued_age_pack_issued_ages_1_T_8 ? reservation_station_8_io_o_uop_imm :
    _io_o_issue_packs_1_T_118_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_src1_value = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_src1_value : _io_o_issue_packs_1_T_118_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_src2_value = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_src2_value : _io_o_issue_packs_1_T_118_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_119_op1_sel = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_op1_sel : _io_o_issue_packs_1_T_118_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_119_op2_sel = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_op2_sel : _io_o_issue_packs_1_T_118_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_alu_sel = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_alu_sel : _io_o_issue_packs_1_T_118_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_119_branch_type = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_branch_type : _io_o_issue_packs_1_T_118_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_119_mem_type = _issued_age_pack_issued_ages_1_T_8 ?
    reservation_station_8_io_o_uop_mem_type : _io_o_issue_packs_1_T_118_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_120_pc = _issued_age_pack_issued_ages_1_T_7 ? reservation_station_7_io_o_uop_pc :
    _io_o_issue_packs_1_T_119_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_120_inst = _issued_age_pack_issued_ages_1_T_7 ? reservation_station_7_io_o_uop_inst
     : _io_o_issue_packs_1_T_119_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_func_code = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_func_code : _io_o_issue_packs_1_T_119_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_119_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_119_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_120_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_119_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_119_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_119_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_phy_dst = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_phy_dst : _io_o_issue_packs_1_T_119_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_stale_dst = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_stale_dst : _io_o_issue_packs_1_T_119_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_arch_dst = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_arch_dst : _io_o_issue_packs_1_T_119_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_120_inst_type = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_inst_type : _io_o_issue_packs_1_T_119_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_regWen = _issued_age_pack_issued_ages_1_T_7 ? reservation_station_7_io_o_uop_regWen :
    _io_o_issue_packs_1_T_119_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_src1_valid = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_src1_valid : _io_o_issue_packs_1_T_119_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_phy_rs1 = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_119_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_arch_rs1 = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_119_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_src2_valid = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_src2_valid : _io_o_issue_packs_1_T_119_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_phy_rs2 = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_119_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_arch_rs2 = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_119_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_rob_idx = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_rob_idx : _io_o_issue_packs_1_T_119_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_imm = _issued_age_pack_issued_ages_1_T_7 ? reservation_station_7_io_o_uop_imm :
    _io_o_issue_packs_1_T_119_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_src1_value = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_src1_value : _io_o_issue_packs_1_T_119_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_src2_value = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_src2_value : _io_o_issue_packs_1_T_119_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_120_op1_sel = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_op1_sel : _io_o_issue_packs_1_T_119_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_120_op2_sel = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_op2_sel : _io_o_issue_packs_1_T_119_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_alu_sel = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_alu_sel : _io_o_issue_packs_1_T_119_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_120_branch_type = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_branch_type : _io_o_issue_packs_1_T_119_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_120_mem_type = _issued_age_pack_issued_ages_1_T_7 ?
    reservation_station_7_io_o_uop_mem_type : _io_o_issue_packs_1_T_119_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_121_pc = _issued_age_pack_issued_ages_1_T_6 ? reservation_station_6_io_o_uop_pc :
    _io_o_issue_packs_1_T_120_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_121_inst = _issued_age_pack_issued_ages_1_T_6 ? reservation_station_6_io_o_uop_inst
     : _io_o_issue_packs_1_T_120_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_func_code = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_func_code : _io_o_issue_packs_1_T_120_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_120_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_120_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_121_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_120_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_120_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_120_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_phy_dst = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_phy_dst : _io_o_issue_packs_1_T_120_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_stale_dst = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_stale_dst : _io_o_issue_packs_1_T_120_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_arch_dst = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_arch_dst : _io_o_issue_packs_1_T_120_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_121_inst_type = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_inst_type : _io_o_issue_packs_1_T_120_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_regWen = _issued_age_pack_issued_ages_1_T_6 ? reservation_station_6_io_o_uop_regWen :
    _io_o_issue_packs_1_T_120_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_src1_valid = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_src1_valid : _io_o_issue_packs_1_T_120_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_phy_rs1 = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_120_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_arch_rs1 = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_120_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_src2_valid = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_src2_valid : _io_o_issue_packs_1_T_120_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_phy_rs2 = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_120_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_arch_rs2 = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_120_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_rob_idx = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_rob_idx : _io_o_issue_packs_1_T_120_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_imm = _issued_age_pack_issued_ages_1_T_6 ? reservation_station_6_io_o_uop_imm :
    _io_o_issue_packs_1_T_120_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_src1_value = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_src1_value : _io_o_issue_packs_1_T_120_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_src2_value = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_src2_value : _io_o_issue_packs_1_T_120_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_121_op1_sel = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_op1_sel : _io_o_issue_packs_1_T_120_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_121_op2_sel = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_op2_sel : _io_o_issue_packs_1_T_120_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_alu_sel = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_alu_sel : _io_o_issue_packs_1_T_120_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_121_branch_type = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_branch_type : _io_o_issue_packs_1_T_120_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_121_mem_type = _issued_age_pack_issued_ages_1_T_6 ?
    reservation_station_6_io_o_uop_mem_type : _io_o_issue_packs_1_T_120_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_122_pc = _issued_age_pack_issued_ages_1_T_5 ? reservation_station_5_io_o_uop_pc :
    _io_o_issue_packs_1_T_121_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_122_inst = _issued_age_pack_issued_ages_1_T_5 ? reservation_station_5_io_o_uop_inst
     : _io_o_issue_packs_1_T_121_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_func_code = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_func_code : _io_o_issue_packs_1_T_121_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_121_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_121_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_122_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_121_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_121_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_121_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_phy_dst = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_phy_dst : _io_o_issue_packs_1_T_121_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_stale_dst = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_stale_dst : _io_o_issue_packs_1_T_121_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_arch_dst = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_arch_dst : _io_o_issue_packs_1_T_121_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_122_inst_type = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_inst_type : _io_o_issue_packs_1_T_121_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_regWen = _issued_age_pack_issued_ages_1_T_5 ? reservation_station_5_io_o_uop_regWen :
    _io_o_issue_packs_1_T_121_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_src1_valid = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_src1_valid : _io_o_issue_packs_1_T_121_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_phy_rs1 = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_121_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_arch_rs1 = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_121_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_src2_valid = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_src2_valid : _io_o_issue_packs_1_T_121_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_phy_rs2 = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_121_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_arch_rs2 = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_121_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_rob_idx = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_rob_idx : _io_o_issue_packs_1_T_121_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_imm = _issued_age_pack_issued_ages_1_T_5 ? reservation_station_5_io_o_uop_imm :
    _io_o_issue_packs_1_T_121_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_src1_value = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_src1_value : _io_o_issue_packs_1_T_121_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_src2_value = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_src2_value : _io_o_issue_packs_1_T_121_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_122_op1_sel = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_op1_sel : _io_o_issue_packs_1_T_121_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_122_op2_sel = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_op2_sel : _io_o_issue_packs_1_T_121_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_alu_sel = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_alu_sel : _io_o_issue_packs_1_T_121_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_122_branch_type = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_branch_type : _io_o_issue_packs_1_T_121_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_122_mem_type = _issued_age_pack_issued_ages_1_T_5 ?
    reservation_station_5_io_o_uop_mem_type : _io_o_issue_packs_1_T_121_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_123_pc = _issued_age_pack_issued_ages_1_T_4 ? reservation_station_4_io_o_uop_pc :
    _io_o_issue_packs_1_T_122_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_123_inst = _issued_age_pack_issued_ages_1_T_4 ? reservation_station_4_io_o_uop_inst
     : _io_o_issue_packs_1_T_122_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_func_code = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_func_code : _io_o_issue_packs_1_T_122_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_122_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_122_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_123_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_122_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_122_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_122_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_phy_dst = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_phy_dst : _io_o_issue_packs_1_T_122_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_stale_dst = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_stale_dst : _io_o_issue_packs_1_T_122_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_arch_dst = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_arch_dst : _io_o_issue_packs_1_T_122_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_123_inst_type = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_inst_type : _io_o_issue_packs_1_T_122_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_regWen = _issued_age_pack_issued_ages_1_T_4 ? reservation_station_4_io_o_uop_regWen :
    _io_o_issue_packs_1_T_122_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_src1_valid = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_src1_valid : _io_o_issue_packs_1_T_122_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_phy_rs1 = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_122_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_arch_rs1 = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_122_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_src2_valid = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_src2_valid : _io_o_issue_packs_1_T_122_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_phy_rs2 = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_122_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_arch_rs2 = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_122_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_rob_idx = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_rob_idx : _io_o_issue_packs_1_T_122_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_imm = _issued_age_pack_issued_ages_1_T_4 ? reservation_station_4_io_o_uop_imm :
    _io_o_issue_packs_1_T_122_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_src1_value = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_src1_value : _io_o_issue_packs_1_T_122_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_src2_value = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_src2_value : _io_o_issue_packs_1_T_122_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_123_op1_sel = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_op1_sel : _io_o_issue_packs_1_T_122_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_123_op2_sel = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_op2_sel : _io_o_issue_packs_1_T_122_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_alu_sel = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_alu_sel : _io_o_issue_packs_1_T_122_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_123_branch_type = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_branch_type : _io_o_issue_packs_1_T_122_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_123_mem_type = _issued_age_pack_issued_ages_1_T_4 ?
    reservation_station_4_io_o_uop_mem_type : _io_o_issue_packs_1_T_122_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_124_pc = _issued_age_pack_issued_ages_1_T_3 ? reservation_station_3_io_o_uop_pc :
    _io_o_issue_packs_1_T_123_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_124_inst = _issued_age_pack_issued_ages_1_T_3 ? reservation_station_3_io_o_uop_inst
     : _io_o_issue_packs_1_T_123_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_func_code = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_func_code : _io_o_issue_packs_1_T_123_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_123_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_123_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_124_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_123_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_123_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_123_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_phy_dst = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_phy_dst : _io_o_issue_packs_1_T_123_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_stale_dst = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_stale_dst : _io_o_issue_packs_1_T_123_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_arch_dst = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_arch_dst : _io_o_issue_packs_1_T_123_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_124_inst_type = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_inst_type : _io_o_issue_packs_1_T_123_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_regWen = _issued_age_pack_issued_ages_1_T_3 ? reservation_station_3_io_o_uop_regWen :
    _io_o_issue_packs_1_T_123_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_src1_valid = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_src1_valid : _io_o_issue_packs_1_T_123_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_phy_rs1 = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_123_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_arch_rs1 = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_123_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_src2_valid = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_src2_valid : _io_o_issue_packs_1_T_123_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_phy_rs2 = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_123_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_arch_rs2 = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_123_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_rob_idx = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_rob_idx : _io_o_issue_packs_1_T_123_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_imm = _issued_age_pack_issued_ages_1_T_3 ? reservation_station_3_io_o_uop_imm :
    _io_o_issue_packs_1_T_123_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_src1_value = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_src1_value : _io_o_issue_packs_1_T_123_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_src2_value = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_src2_value : _io_o_issue_packs_1_T_123_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_124_op1_sel = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_op1_sel : _io_o_issue_packs_1_T_123_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_124_op2_sel = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_op2_sel : _io_o_issue_packs_1_T_123_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_alu_sel = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_alu_sel : _io_o_issue_packs_1_T_123_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_124_branch_type = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_branch_type : _io_o_issue_packs_1_T_123_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_124_mem_type = _issued_age_pack_issued_ages_1_T_3 ?
    reservation_station_3_io_o_uop_mem_type : _io_o_issue_packs_1_T_123_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_125_pc = _issued_age_pack_issued_ages_1_T_2 ? reservation_station_2_io_o_uop_pc :
    _io_o_issue_packs_1_T_124_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_125_inst = _issued_age_pack_issued_ages_1_T_2 ? reservation_station_2_io_o_uop_inst
     : _io_o_issue_packs_1_T_124_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_func_code = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_func_code : _io_o_issue_packs_1_T_124_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_124_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_124_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_125_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_124_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_124_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_124_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_phy_dst = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_phy_dst : _io_o_issue_packs_1_T_124_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_stale_dst = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_stale_dst : _io_o_issue_packs_1_T_124_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_arch_dst = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_arch_dst : _io_o_issue_packs_1_T_124_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_125_inst_type = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_inst_type : _io_o_issue_packs_1_T_124_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_regWen = _issued_age_pack_issued_ages_1_T_2 ? reservation_station_2_io_o_uop_regWen :
    _io_o_issue_packs_1_T_124_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_src1_valid = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_src1_valid : _io_o_issue_packs_1_T_124_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_phy_rs1 = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_124_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_arch_rs1 = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_124_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_src2_valid = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_src2_valid : _io_o_issue_packs_1_T_124_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_phy_rs2 = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_124_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_arch_rs2 = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_124_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_rob_idx = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_rob_idx : _io_o_issue_packs_1_T_124_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_imm = _issued_age_pack_issued_ages_1_T_2 ? reservation_station_2_io_o_uop_imm :
    _io_o_issue_packs_1_T_124_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_src1_value = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_src1_value : _io_o_issue_packs_1_T_124_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_src2_value = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_src2_value : _io_o_issue_packs_1_T_124_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_125_op1_sel = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_op1_sel : _io_o_issue_packs_1_T_124_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_125_op2_sel = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_op2_sel : _io_o_issue_packs_1_T_124_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_alu_sel = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_alu_sel : _io_o_issue_packs_1_T_124_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_125_branch_type = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_branch_type : _io_o_issue_packs_1_T_124_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_125_mem_type = _issued_age_pack_issued_ages_1_T_2 ?
    reservation_station_2_io_o_uop_mem_type : _io_o_issue_packs_1_T_124_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_126_pc = _issued_age_pack_issued_ages_1_T_1 ? reservation_station_1_io_o_uop_pc :
    _io_o_issue_packs_1_T_125_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_126_inst = _issued_age_pack_issued_ages_1_T_1 ? reservation_station_1_io_o_uop_inst
     : _io_o_issue_packs_1_T_125_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_func_code = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_func_code : _io_o_issue_packs_1_T_125_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_125_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_125_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_126_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_125_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_125_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_125_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_phy_dst = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_phy_dst : _io_o_issue_packs_1_T_125_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_stale_dst = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_stale_dst : _io_o_issue_packs_1_T_125_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_arch_dst = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_arch_dst : _io_o_issue_packs_1_T_125_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_126_inst_type = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_inst_type : _io_o_issue_packs_1_T_125_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_regWen = _issued_age_pack_issued_ages_1_T_1 ? reservation_station_1_io_o_uop_regWen :
    _io_o_issue_packs_1_T_125_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_src1_valid = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_src1_valid : _io_o_issue_packs_1_T_125_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_phy_rs1 = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_phy_rs1 : _io_o_issue_packs_1_T_125_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_arch_rs1 = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_arch_rs1 : _io_o_issue_packs_1_T_125_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_src2_valid = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_src2_valid : _io_o_issue_packs_1_T_125_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_phy_rs2 = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_phy_rs2 : _io_o_issue_packs_1_T_125_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_arch_rs2 = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_arch_rs2 : _io_o_issue_packs_1_T_125_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_rob_idx = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_rob_idx : _io_o_issue_packs_1_T_125_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_imm = _issued_age_pack_issued_ages_1_T_1 ? reservation_station_1_io_o_uop_imm :
    _io_o_issue_packs_1_T_125_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_src1_value = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_src1_value : _io_o_issue_packs_1_T_125_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_src2_value = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_src2_value : _io_o_issue_packs_1_T_125_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_126_op1_sel = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_op1_sel : _io_o_issue_packs_1_T_125_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_126_op2_sel = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_op2_sel : _io_o_issue_packs_1_T_125_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_alu_sel = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_alu_sel : _io_o_issue_packs_1_T_125_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_126_branch_type = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_branch_type : _io_o_issue_packs_1_T_125_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_126_mem_type = _issued_age_pack_issued_ages_1_T_1 ?
    reservation_station_1_io_o_uop_mem_type : _io_o_issue_packs_1_T_125_mem_type; // @[Mux.scala 101:16]
  wire  _reservation_station_0_io_i_write_slot_T = 6'h0 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_0_io_i_write_slot_T_1 = 6'h0 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_1_io_i_write_slot_T = 6'h1 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_1_io_i_write_slot_T_1 = 6'h1 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_2_io_i_write_slot_T = 6'h2 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_2_io_i_write_slot_T_1 = 6'h2 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_3_io_i_write_slot_T = 6'h3 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_3_io_i_write_slot_T_1 = 6'h3 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_4_io_i_write_slot_T = 6'h4 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_4_io_i_write_slot_T_1 = 6'h4 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_5_io_i_write_slot_T = 6'h5 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_5_io_i_write_slot_T_1 = 6'h5 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_6_io_i_write_slot_T = 6'h6 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_6_io_i_write_slot_T_1 = 6'h6 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_7_io_i_write_slot_T = 6'h7 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_7_io_i_write_slot_T_1 = 6'h7 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_8_io_i_write_slot_T = 6'h8 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_8_io_i_write_slot_T_1 = 6'h8 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_9_io_i_write_slot_T = 6'h9 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_9_io_i_write_slot_T_1 = 6'h9 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_10_io_i_write_slot_T = 6'ha == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_10_io_i_write_slot_T_1 = 6'ha == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_11_io_i_write_slot_T = 6'hb == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_11_io_i_write_slot_T_1 = 6'hb == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_12_io_i_write_slot_T = 6'hc == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_12_io_i_write_slot_T_1 = 6'hc == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_13_io_i_write_slot_T = 6'hd == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_13_io_i_write_slot_T_1 = 6'hd == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_14_io_i_write_slot_T = 6'he == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_14_io_i_write_slot_T_1 = 6'he == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_15_io_i_write_slot_T = 6'hf == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_15_io_i_write_slot_T_1 = 6'hf == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_16_io_i_write_slot_T = 6'h10 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_16_io_i_write_slot_T_1 = 6'h10 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_17_io_i_write_slot_T = 6'h11 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_17_io_i_write_slot_T_1 = 6'h11 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_18_io_i_write_slot_T = 6'h12 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_18_io_i_write_slot_T_1 = 6'h12 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_19_io_i_write_slot_T = 6'h13 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_19_io_i_write_slot_T_1 = 6'h13 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_20_io_i_write_slot_T = 6'h14 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_20_io_i_write_slot_T_1 = 6'h14 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_21_io_i_write_slot_T = 6'h15 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_21_io_i_write_slot_T_1 = 6'h15 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_22_io_i_write_slot_T = 6'h16 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_22_io_i_write_slot_T_1 = 6'h16 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_23_io_i_write_slot_T = 6'h17 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_23_io_i_write_slot_T_1 = 6'h17 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_24_io_i_write_slot_T = 6'h18 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_24_io_i_write_slot_T_1 = 6'h18 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_25_io_i_write_slot_T = 6'h19 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_25_io_i_write_slot_T_1 = 6'h19 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_26_io_i_write_slot_T = 6'h1a == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_26_io_i_write_slot_T_1 = 6'h1a == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_27_io_i_write_slot_T = 6'h1b == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_27_io_i_write_slot_T_1 = 6'h1b == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_28_io_i_write_slot_T = 6'h1c == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_28_io_i_write_slot_T_1 = 6'h1c == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_29_io_i_write_slot_T = 6'h1d == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_29_io_i_write_slot_T_1 = 6'h1d == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_30_io_i_write_slot_T = 6'h1e == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_30_io_i_write_slot_T_1 = 6'h1e == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_31_io_i_write_slot_T = 6'h1f == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_31_io_i_write_slot_T_1 = 6'h1f == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_32_io_i_write_slot_T = 6'h20 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_32_io_i_write_slot_T_1 = 6'h20 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_33_io_i_write_slot_T = 6'h21 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_33_io_i_write_slot_T_1 = 6'h21 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_34_io_i_write_slot_T = 6'h22 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_34_io_i_write_slot_T_1 = 6'h22 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_35_io_i_write_slot_T = 6'h23 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_35_io_i_write_slot_T_1 = 6'h23 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_36_io_i_write_slot_T = 6'h24 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_36_io_i_write_slot_T_1 = 6'h24 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_37_io_i_write_slot_T = 6'h25 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_37_io_i_write_slot_T_1 = 6'h25 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_38_io_i_write_slot_T = 6'h26 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_38_io_i_write_slot_T_1 = 6'h26 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_39_io_i_write_slot_T = 6'h27 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_39_io_i_write_slot_T_1 = 6'h27 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_40_io_i_write_slot_T = 6'h28 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_40_io_i_write_slot_T_1 = 6'h28 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_41_io_i_write_slot_T = 6'h29 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_41_io_i_write_slot_T_1 = 6'h29 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_42_io_i_write_slot_T = 6'h2a == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_42_io_i_write_slot_T_1 = 6'h2a == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_43_io_i_write_slot_T = 6'h2b == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_43_io_i_write_slot_T_1 = 6'h2b == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_44_io_i_write_slot_T = 6'h2c == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_44_io_i_write_slot_T_1 = 6'h2c == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_45_io_i_write_slot_T = 6'h2d == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_45_io_i_write_slot_T_1 = 6'h2d == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_46_io_i_write_slot_T = 6'h2e == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_46_io_i_write_slot_T_1 = 6'h2e == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_47_io_i_write_slot_T = 6'h2f == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_47_io_i_write_slot_T_1 = 6'h2f == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_48_io_i_write_slot_T = 6'h30 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_48_io_i_write_slot_T_1 = 6'h30 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_49_io_i_write_slot_T = 6'h31 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_49_io_i_write_slot_T_1 = 6'h31 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_50_io_i_write_slot_T = 6'h32 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_50_io_i_write_slot_T_1 = 6'h32 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_51_io_i_write_slot_T = 6'h33 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_51_io_i_write_slot_T_1 = 6'h33 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_52_io_i_write_slot_T = 6'h34 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_52_io_i_write_slot_T_1 = 6'h34 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_53_io_i_write_slot_T = 6'h35 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_53_io_i_write_slot_T_1 = 6'h35 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_54_io_i_write_slot_T = 6'h36 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_54_io_i_write_slot_T_1 = 6'h36 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_55_io_i_write_slot_T = 6'h37 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_55_io_i_write_slot_T_1 = 6'h37 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_56_io_i_write_slot_T = 6'h38 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_56_io_i_write_slot_T_1 = 6'h38 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_57_io_i_write_slot_T = 6'h39 == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_57_io_i_write_slot_T_1 = 6'h39 == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_58_io_i_write_slot_T = 6'h3a == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_58_io_i_write_slot_T_1 = 6'h3a == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_59_io_i_write_slot_T = 6'h3b == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_59_io_i_write_slot_T_1 = 6'h3b == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_60_io_i_write_slot_T = 6'h3c == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_60_io_i_write_slot_T_1 = 6'h3c == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_61_io_i_write_slot_T = 6'h3d == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_61_io_i_write_slot_T_1 = 6'h3d == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_62_io_i_write_slot_T = 6'h3e == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_62_io_i_write_slot_T_1 = 6'h3e == write_idx2; // @[reservation_station.scala 249:13]
  wire  _reservation_station_63_io_i_write_slot_T = 6'h3f == write_idx1; // @[reservation_station.scala 248:13]
  wire  _reservation_station_63_io_i_write_slot_T_1 = 6'h3f == write_idx2; // @[reservation_station.scala 249:13]
  Reservation_Station_Slot reservation_station_0 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_0_clock),
    .reset(reservation_station_0_reset),
    .io_o_valid(reservation_station_0_io_o_valid),
    .io_o_ready_to_issue(reservation_station_0_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_0_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_0_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_0_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_0_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_0_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_0_io_i_exception),
    .io_i_write_slot(reservation_station_0_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_0_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_0_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_0_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_0_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_0_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_0_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_0_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_0_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_0_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_0_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_0_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_0_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_0_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_0_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_0_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_0_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_0_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_0_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_0_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_0_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_0_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_0_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_0_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_0_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_0_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_0_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_0_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_0_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_0_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_0_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_0_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_0_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_0_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_0_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_0_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_0_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_0_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_0_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_0_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_0_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_0_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_0_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_0_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_0_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_0_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_0_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_0_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_0_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_0_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_0_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_0_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_0_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_0_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_0_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_0_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_0_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_0_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_0_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_0_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_0_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_0_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_0_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_0_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_0_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_0_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_0_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_0_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_0_io_o_age),
    .io_i_ROB_first_entry(reservation_station_0_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_1 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_1_clock),
    .reset(reservation_station_1_reset),
    .io_o_valid(reservation_station_1_io_o_valid),
    .io_o_ready_to_issue(reservation_station_1_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_1_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_1_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_1_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_1_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_1_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_1_io_i_exception),
    .io_i_write_slot(reservation_station_1_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_1_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_1_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_1_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_1_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_1_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_1_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_1_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_1_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_1_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_1_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_1_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_1_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_1_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_1_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_1_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_1_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_1_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_1_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_1_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_1_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_1_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_1_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_1_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_1_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_1_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_1_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_1_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_1_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_1_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_1_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_1_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_1_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_1_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_1_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_1_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_1_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_1_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_1_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_1_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_1_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_1_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_1_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_1_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_1_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_1_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_1_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_1_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_1_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_1_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_1_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_1_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_1_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_1_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_1_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_1_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_1_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_1_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_1_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_1_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_1_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_1_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_1_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_1_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_1_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_1_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_1_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_1_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_1_io_o_age),
    .io_i_ROB_first_entry(reservation_station_1_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_2 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_2_clock),
    .reset(reservation_station_2_reset),
    .io_o_valid(reservation_station_2_io_o_valid),
    .io_o_ready_to_issue(reservation_station_2_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_2_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_2_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_2_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_2_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_2_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_2_io_i_exception),
    .io_i_write_slot(reservation_station_2_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_2_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_2_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_2_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_2_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_2_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_2_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_2_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_2_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_2_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_2_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_2_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_2_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_2_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_2_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_2_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_2_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_2_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_2_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_2_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_2_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_2_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_2_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_2_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_2_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_2_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_2_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_2_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_2_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_2_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_2_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_2_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_2_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_2_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_2_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_2_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_2_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_2_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_2_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_2_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_2_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_2_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_2_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_2_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_2_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_2_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_2_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_2_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_2_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_2_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_2_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_2_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_2_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_2_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_2_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_2_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_2_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_2_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_2_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_2_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_2_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_2_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_2_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_2_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_2_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_2_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_2_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_2_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_2_io_o_age),
    .io_i_ROB_first_entry(reservation_station_2_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_3 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_3_clock),
    .reset(reservation_station_3_reset),
    .io_o_valid(reservation_station_3_io_o_valid),
    .io_o_ready_to_issue(reservation_station_3_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_3_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_3_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_3_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_3_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_3_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_3_io_i_exception),
    .io_i_write_slot(reservation_station_3_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_3_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_3_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_3_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_3_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_3_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_3_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_3_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_3_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_3_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_3_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_3_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_3_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_3_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_3_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_3_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_3_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_3_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_3_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_3_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_3_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_3_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_3_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_3_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_3_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_3_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_3_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_3_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_3_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_3_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_3_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_3_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_3_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_3_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_3_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_3_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_3_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_3_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_3_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_3_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_3_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_3_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_3_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_3_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_3_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_3_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_3_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_3_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_3_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_3_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_3_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_3_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_3_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_3_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_3_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_3_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_3_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_3_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_3_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_3_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_3_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_3_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_3_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_3_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_3_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_3_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_3_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_3_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_3_io_o_age),
    .io_i_ROB_first_entry(reservation_station_3_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_4 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_4_clock),
    .reset(reservation_station_4_reset),
    .io_o_valid(reservation_station_4_io_o_valid),
    .io_o_ready_to_issue(reservation_station_4_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_4_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_4_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_4_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_4_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_4_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_4_io_i_exception),
    .io_i_write_slot(reservation_station_4_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_4_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_4_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_4_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_4_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_4_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_4_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_4_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_4_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_4_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_4_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_4_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_4_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_4_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_4_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_4_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_4_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_4_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_4_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_4_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_4_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_4_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_4_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_4_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_4_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_4_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_4_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_4_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_4_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_4_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_4_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_4_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_4_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_4_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_4_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_4_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_4_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_4_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_4_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_4_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_4_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_4_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_4_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_4_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_4_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_4_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_4_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_4_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_4_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_4_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_4_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_4_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_4_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_4_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_4_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_4_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_4_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_4_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_4_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_4_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_4_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_4_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_4_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_4_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_4_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_4_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_4_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_4_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_4_io_o_age),
    .io_i_ROB_first_entry(reservation_station_4_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_5 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_5_clock),
    .reset(reservation_station_5_reset),
    .io_o_valid(reservation_station_5_io_o_valid),
    .io_o_ready_to_issue(reservation_station_5_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_5_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_5_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_5_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_5_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_5_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_5_io_i_exception),
    .io_i_write_slot(reservation_station_5_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_5_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_5_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_5_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_5_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_5_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_5_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_5_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_5_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_5_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_5_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_5_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_5_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_5_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_5_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_5_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_5_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_5_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_5_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_5_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_5_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_5_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_5_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_5_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_5_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_5_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_5_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_5_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_5_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_5_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_5_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_5_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_5_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_5_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_5_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_5_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_5_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_5_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_5_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_5_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_5_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_5_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_5_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_5_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_5_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_5_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_5_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_5_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_5_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_5_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_5_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_5_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_5_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_5_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_5_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_5_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_5_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_5_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_5_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_5_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_5_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_5_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_5_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_5_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_5_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_5_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_5_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_5_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_5_io_o_age),
    .io_i_ROB_first_entry(reservation_station_5_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_6 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_6_clock),
    .reset(reservation_station_6_reset),
    .io_o_valid(reservation_station_6_io_o_valid),
    .io_o_ready_to_issue(reservation_station_6_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_6_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_6_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_6_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_6_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_6_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_6_io_i_exception),
    .io_i_write_slot(reservation_station_6_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_6_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_6_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_6_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_6_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_6_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_6_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_6_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_6_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_6_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_6_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_6_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_6_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_6_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_6_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_6_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_6_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_6_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_6_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_6_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_6_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_6_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_6_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_6_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_6_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_6_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_6_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_6_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_6_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_6_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_6_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_6_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_6_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_6_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_6_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_6_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_6_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_6_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_6_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_6_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_6_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_6_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_6_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_6_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_6_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_6_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_6_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_6_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_6_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_6_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_6_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_6_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_6_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_6_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_6_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_6_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_6_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_6_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_6_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_6_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_6_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_6_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_6_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_6_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_6_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_6_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_6_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_6_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_6_io_o_age),
    .io_i_ROB_first_entry(reservation_station_6_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_7 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_7_clock),
    .reset(reservation_station_7_reset),
    .io_o_valid(reservation_station_7_io_o_valid),
    .io_o_ready_to_issue(reservation_station_7_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_7_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_7_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_7_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_7_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_7_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_7_io_i_exception),
    .io_i_write_slot(reservation_station_7_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_7_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_7_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_7_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_7_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_7_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_7_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_7_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_7_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_7_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_7_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_7_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_7_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_7_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_7_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_7_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_7_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_7_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_7_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_7_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_7_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_7_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_7_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_7_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_7_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_7_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_7_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_7_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_7_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_7_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_7_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_7_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_7_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_7_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_7_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_7_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_7_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_7_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_7_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_7_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_7_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_7_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_7_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_7_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_7_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_7_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_7_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_7_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_7_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_7_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_7_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_7_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_7_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_7_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_7_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_7_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_7_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_7_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_7_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_7_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_7_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_7_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_7_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_7_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_7_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_7_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_7_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_7_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_7_io_o_age),
    .io_i_ROB_first_entry(reservation_station_7_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_8 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_8_clock),
    .reset(reservation_station_8_reset),
    .io_o_valid(reservation_station_8_io_o_valid),
    .io_o_ready_to_issue(reservation_station_8_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_8_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_8_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_8_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_8_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_8_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_8_io_i_exception),
    .io_i_write_slot(reservation_station_8_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_8_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_8_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_8_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_8_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_8_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_8_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_8_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_8_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_8_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_8_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_8_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_8_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_8_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_8_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_8_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_8_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_8_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_8_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_8_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_8_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_8_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_8_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_8_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_8_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_8_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_8_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_8_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_8_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_8_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_8_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_8_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_8_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_8_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_8_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_8_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_8_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_8_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_8_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_8_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_8_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_8_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_8_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_8_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_8_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_8_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_8_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_8_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_8_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_8_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_8_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_8_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_8_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_8_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_8_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_8_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_8_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_8_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_8_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_8_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_8_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_8_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_8_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_8_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_8_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_8_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_8_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_8_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_8_io_o_age),
    .io_i_ROB_first_entry(reservation_station_8_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_9 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_9_clock),
    .reset(reservation_station_9_reset),
    .io_o_valid(reservation_station_9_io_o_valid),
    .io_o_ready_to_issue(reservation_station_9_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_9_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_9_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_9_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_9_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_9_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_9_io_i_exception),
    .io_i_write_slot(reservation_station_9_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_9_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_9_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_9_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_9_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_9_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_9_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_9_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_9_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_9_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_9_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_9_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_9_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_9_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_9_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_9_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_9_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_9_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_9_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_9_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_9_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_9_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_9_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_9_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_9_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_9_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_9_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_9_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_9_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_9_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_9_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_9_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_9_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_9_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_9_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_9_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_9_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_9_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_9_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_9_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_9_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_9_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_9_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_9_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_9_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_9_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_9_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_9_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_9_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_9_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_9_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_9_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_9_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_9_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_9_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_9_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_9_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_9_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_9_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_9_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_9_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_9_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_9_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_9_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_9_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_9_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_9_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_9_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_9_io_o_age),
    .io_i_ROB_first_entry(reservation_station_9_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_10 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_10_clock),
    .reset(reservation_station_10_reset),
    .io_o_valid(reservation_station_10_io_o_valid),
    .io_o_ready_to_issue(reservation_station_10_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_10_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_10_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_10_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_10_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_10_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_10_io_i_exception),
    .io_i_write_slot(reservation_station_10_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_10_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_10_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_10_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_10_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_10_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_10_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_10_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_10_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_10_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_10_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_10_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_10_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_10_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_10_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_10_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_10_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_10_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_10_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_10_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_10_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_10_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_10_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_10_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_10_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_10_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_10_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_10_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_10_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_10_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_10_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_10_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_10_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_10_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_10_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_10_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_10_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_10_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_10_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_10_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_10_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_10_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_10_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_10_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_10_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_10_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_10_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_10_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_10_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_10_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_10_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_10_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_10_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_10_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_10_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_10_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_10_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_10_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_10_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_10_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_10_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_10_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_10_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_10_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_10_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_10_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_10_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_10_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_10_io_o_age),
    .io_i_ROB_first_entry(reservation_station_10_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_11 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_11_clock),
    .reset(reservation_station_11_reset),
    .io_o_valid(reservation_station_11_io_o_valid),
    .io_o_ready_to_issue(reservation_station_11_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_11_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_11_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_11_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_11_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_11_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_11_io_i_exception),
    .io_i_write_slot(reservation_station_11_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_11_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_11_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_11_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_11_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_11_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_11_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_11_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_11_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_11_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_11_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_11_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_11_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_11_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_11_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_11_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_11_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_11_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_11_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_11_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_11_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_11_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_11_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_11_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_11_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_11_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_11_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_11_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_11_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_11_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_11_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_11_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_11_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_11_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_11_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_11_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_11_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_11_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_11_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_11_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_11_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_11_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_11_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_11_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_11_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_11_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_11_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_11_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_11_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_11_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_11_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_11_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_11_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_11_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_11_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_11_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_11_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_11_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_11_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_11_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_11_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_11_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_11_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_11_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_11_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_11_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_11_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_11_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_11_io_o_age),
    .io_i_ROB_first_entry(reservation_station_11_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_12 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_12_clock),
    .reset(reservation_station_12_reset),
    .io_o_valid(reservation_station_12_io_o_valid),
    .io_o_ready_to_issue(reservation_station_12_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_12_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_12_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_12_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_12_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_12_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_12_io_i_exception),
    .io_i_write_slot(reservation_station_12_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_12_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_12_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_12_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_12_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_12_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_12_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_12_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_12_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_12_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_12_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_12_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_12_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_12_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_12_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_12_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_12_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_12_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_12_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_12_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_12_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_12_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_12_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_12_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_12_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_12_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_12_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_12_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_12_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_12_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_12_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_12_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_12_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_12_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_12_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_12_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_12_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_12_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_12_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_12_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_12_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_12_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_12_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_12_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_12_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_12_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_12_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_12_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_12_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_12_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_12_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_12_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_12_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_12_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_12_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_12_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_12_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_12_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_12_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_12_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_12_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_12_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_12_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_12_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_12_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_12_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_12_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_12_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_12_io_o_age),
    .io_i_ROB_first_entry(reservation_station_12_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_13 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_13_clock),
    .reset(reservation_station_13_reset),
    .io_o_valid(reservation_station_13_io_o_valid),
    .io_o_ready_to_issue(reservation_station_13_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_13_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_13_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_13_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_13_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_13_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_13_io_i_exception),
    .io_i_write_slot(reservation_station_13_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_13_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_13_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_13_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_13_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_13_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_13_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_13_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_13_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_13_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_13_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_13_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_13_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_13_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_13_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_13_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_13_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_13_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_13_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_13_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_13_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_13_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_13_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_13_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_13_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_13_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_13_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_13_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_13_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_13_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_13_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_13_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_13_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_13_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_13_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_13_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_13_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_13_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_13_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_13_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_13_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_13_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_13_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_13_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_13_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_13_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_13_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_13_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_13_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_13_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_13_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_13_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_13_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_13_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_13_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_13_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_13_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_13_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_13_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_13_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_13_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_13_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_13_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_13_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_13_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_13_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_13_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_13_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_13_io_o_age),
    .io_i_ROB_first_entry(reservation_station_13_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_14 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_14_clock),
    .reset(reservation_station_14_reset),
    .io_o_valid(reservation_station_14_io_o_valid),
    .io_o_ready_to_issue(reservation_station_14_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_14_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_14_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_14_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_14_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_14_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_14_io_i_exception),
    .io_i_write_slot(reservation_station_14_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_14_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_14_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_14_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_14_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_14_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_14_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_14_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_14_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_14_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_14_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_14_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_14_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_14_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_14_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_14_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_14_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_14_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_14_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_14_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_14_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_14_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_14_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_14_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_14_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_14_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_14_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_14_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_14_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_14_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_14_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_14_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_14_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_14_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_14_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_14_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_14_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_14_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_14_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_14_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_14_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_14_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_14_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_14_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_14_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_14_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_14_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_14_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_14_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_14_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_14_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_14_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_14_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_14_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_14_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_14_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_14_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_14_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_14_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_14_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_14_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_14_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_14_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_14_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_14_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_14_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_14_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_14_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_14_io_o_age),
    .io_i_ROB_first_entry(reservation_station_14_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_15 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_15_clock),
    .reset(reservation_station_15_reset),
    .io_o_valid(reservation_station_15_io_o_valid),
    .io_o_ready_to_issue(reservation_station_15_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_15_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_15_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_15_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_15_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_15_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_15_io_i_exception),
    .io_i_write_slot(reservation_station_15_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_15_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_15_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_15_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_15_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_15_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_15_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_15_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_15_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_15_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_15_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_15_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_15_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_15_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_15_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_15_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_15_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_15_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_15_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_15_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_15_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_15_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_15_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_15_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_15_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_15_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_15_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_15_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_15_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_15_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_15_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_15_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_15_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_15_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_15_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_15_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_15_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_15_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_15_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_15_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_15_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_15_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_15_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_15_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_15_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_15_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_15_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_15_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_15_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_15_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_15_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_15_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_15_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_15_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_15_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_15_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_15_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_15_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_15_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_15_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_15_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_15_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_15_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_15_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_15_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_15_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_15_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_15_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_15_io_o_age),
    .io_i_ROB_first_entry(reservation_station_15_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_16 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_16_clock),
    .reset(reservation_station_16_reset),
    .io_o_valid(reservation_station_16_io_o_valid),
    .io_o_ready_to_issue(reservation_station_16_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_16_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_16_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_16_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_16_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_16_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_16_io_i_exception),
    .io_i_write_slot(reservation_station_16_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_16_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_16_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_16_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_16_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_16_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_16_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_16_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_16_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_16_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_16_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_16_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_16_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_16_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_16_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_16_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_16_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_16_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_16_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_16_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_16_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_16_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_16_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_16_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_16_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_16_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_16_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_16_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_16_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_16_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_16_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_16_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_16_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_16_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_16_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_16_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_16_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_16_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_16_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_16_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_16_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_16_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_16_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_16_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_16_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_16_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_16_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_16_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_16_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_16_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_16_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_16_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_16_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_16_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_16_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_16_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_16_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_16_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_16_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_16_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_16_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_16_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_16_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_16_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_16_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_16_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_16_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_16_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_16_io_o_age),
    .io_i_ROB_first_entry(reservation_station_16_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_17 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_17_clock),
    .reset(reservation_station_17_reset),
    .io_o_valid(reservation_station_17_io_o_valid),
    .io_o_ready_to_issue(reservation_station_17_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_17_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_17_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_17_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_17_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_17_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_17_io_i_exception),
    .io_i_write_slot(reservation_station_17_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_17_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_17_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_17_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_17_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_17_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_17_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_17_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_17_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_17_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_17_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_17_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_17_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_17_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_17_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_17_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_17_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_17_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_17_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_17_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_17_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_17_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_17_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_17_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_17_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_17_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_17_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_17_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_17_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_17_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_17_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_17_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_17_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_17_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_17_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_17_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_17_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_17_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_17_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_17_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_17_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_17_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_17_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_17_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_17_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_17_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_17_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_17_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_17_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_17_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_17_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_17_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_17_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_17_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_17_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_17_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_17_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_17_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_17_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_17_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_17_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_17_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_17_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_17_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_17_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_17_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_17_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_17_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_17_io_o_age),
    .io_i_ROB_first_entry(reservation_station_17_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_18 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_18_clock),
    .reset(reservation_station_18_reset),
    .io_o_valid(reservation_station_18_io_o_valid),
    .io_o_ready_to_issue(reservation_station_18_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_18_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_18_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_18_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_18_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_18_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_18_io_i_exception),
    .io_i_write_slot(reservation_station_18_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_18_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_18_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_18_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_18_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_18_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_18_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_18_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_18_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_18_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_18_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_18_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_18_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_18_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_18_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_18_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_18_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_18_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_18_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_18_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_18_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_18_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_18_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_18_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_18_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_18_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_18_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_18_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_18_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_18_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_18_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_18_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_18_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_18_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_18_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_18_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_18_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_18_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_18_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_18_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_18_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_18_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_18_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_18_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_18_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_18_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_18_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_18_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_18_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_18_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_18_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_18_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_18_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_18_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_18_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_18_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_18_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_18_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_18_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_18_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_18_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_18_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_18_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_18_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_18_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_18_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_18_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_18_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_18_io_o_age),
    .io_i_ROB_first_entry(reservation_station_18_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_19 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_19_clock),
    .reset(reservation_station_19_reset),
    .io_o_valid(reservation_station_19_io_o_valid),
    .io_o_ready_to_issue(reservation_station_19_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_19_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_19_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_19_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_19_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_19_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_19_io_i_exception),
    .io_i_write_slot(reservation_station_19_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_19_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_19_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_19_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_19_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_19_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_19_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_19_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_19_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_19_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_19_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_19_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_19_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_19_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_19_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_19_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_19_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_19_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_19_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_19_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_19_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_19_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_19_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_19_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_19_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_19_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_19_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_19_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_19_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_19_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_19_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_19_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_19_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_19_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_19_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_19_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_19_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_19_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_19_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_19_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_19_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_19_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_19_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_19_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_19_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_19_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_19_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_19_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_19_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_19_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_19_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_19_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_19_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_19_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_19_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_19_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_19_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_19_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_19_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_19_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_19_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_19_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_19_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_19_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_19_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_19_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_19_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_19_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_19_io_o_age),
    .io_i_ROB_first_entry(reservation_station_19_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_20 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_20_clock),
    .reset(reservation_station_20_reset),
    .io_o_valid(reservation_station_20_io_o_valid),
    .io_o_ready_to_issue(reservation_station_20_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_20_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_20_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_20_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_20_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_20_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_20_io_i_exception),
    .io_i_write_slot(reservation_station_20_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_20_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_20_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_20_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_20_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_20_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_20_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_20_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_20_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_20_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_20_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_20_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_20_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_20_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_20_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_20_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_20_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_20_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_20_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_20_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_20_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_20_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_20_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_20_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_20_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_20_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_20_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_20_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_20_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_20_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_20_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_20_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_20_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_20_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_20_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_20_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_20_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_20_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_20_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_20_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_20_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_20_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_20_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_20_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_20_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_20_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_20_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_20_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_20_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_20_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_20_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_20_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_20_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_20_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_20_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_20_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_20_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_20_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_20_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_20_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_20_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_20_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_20_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_20_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_20_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_20_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_20_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_20_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_20_io_o_age),
    .io_i_ROB_first_entry(reservation_station_20_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_21 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_21_clock),
    .reset(reservation_station_21_reset),
    .io_o_valid(reservation_station_21_io_o_valid),
    .io_o_ready_to_issue(reservation_station_21_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_21_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_21_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_21_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_21_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_21_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_21_io_i_exception),
    .io_i_write_slot(reservation_station_21_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_21_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_21_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_21_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_21_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_21_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_21_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_21_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_21_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_21_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_21_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_21_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_21_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_21_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_21_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_21_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_21_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_21_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_21_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_21_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_21_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_21_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_21_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_21_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_21_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_21_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_21_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_21_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_21_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_21_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_21_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_21_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_21_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_21_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_21_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_21_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_21_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_21_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_21_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_21_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_21_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_21_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_21_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_21_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_21_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_21_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_21_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_21_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_21_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_21_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_21_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_21_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_21_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_21_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_21_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_21_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_21_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_21_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_21_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_21_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_21_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_21_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_21_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_21_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_21_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_21_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_21_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_21_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_21_io_o_age),
    .io_i_ROB_first_entry(reservation_station_21_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_22 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_22_clock),
    .reset(reservation_station_22_reset),
    .io_o_valid(reservation_station_22_io_o_valid),
    .io_o_ready_to_issue(reservation_station_22_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_22_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_22_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_22_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_22_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_22_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_22_io_i_exception),
    .io_i_write_slot(reservation_station_22_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_22_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_22_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_22_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_22_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_22_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_22_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_22_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_22_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_22_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_22_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_22_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_22_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_22_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_22_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_22_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_22_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_22_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_22_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_22_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_22_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_22_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_22_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_22_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_22_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_22_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_22_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_22_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_22_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_22_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_22_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_22_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_22_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_22_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_22_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_22_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_22_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_22_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_22_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_22_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_22_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_22_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_22_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_22_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_22_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_22_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_22_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_22_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_22_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_22_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_22_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_22_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_22_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_22_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_22_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_22_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_22_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_22_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_22_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_22_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_22_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_22_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_22_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_22_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_22_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_22_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_22_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_22_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_22_io_o_age),
    .io_i_ROB_first_entry(reservation_station_22_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_23 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_23_clock),
    .reset(reservation_station_23_reset),
    .io_o_valid(reservation_station_23_io_o_valid),
    .io_o_ready_to_issue(reservation_station_23_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_23_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_23_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_23_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_23_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_23_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_23_io_i_exception),
    .io_i_write_slot(reservation_station_23_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_23_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_23_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_23_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_23_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_23_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_23_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_23_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_23_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_23_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_23_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_23_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_23_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_23_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_23_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_23_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_23_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_23_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_23_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_23_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_23_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_23_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_23_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_23_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_23_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_23_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_23_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_23_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_23_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_23_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_23_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_23_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_23_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_23_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_23_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_23_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_23_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_23_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_23_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_23_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_23_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_23_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_23_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_23_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_23_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_23_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_23_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_23_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_23_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_23_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_23_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_23_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_23_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_23_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_23_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_23_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_23_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_23_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_23_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_23_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_23_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_23_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_23_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_23_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_23_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_23_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_23_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_23_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_23_io_o_age),
    .io_i_ROB_first_entry(reservation_station_23_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_24 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_24_clock),
    .reset(reservation_station_24_reset),
    .io_o_valid(reservation_station_24_io_o_valid),
    .io_o_ready_to_issue(reservation_station_24_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_24_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_24_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_24_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_24_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_24_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_24_io_i_exception),
    .io_i_write_slot(reservation_station_24_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_24_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_24_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_24_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_24_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_24_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_24_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_24_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_24_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_24_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_24_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_24_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_24_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_24_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_24_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_24_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_24_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_24_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_24_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_24_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_24_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_24_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_24_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_24_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_24_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_24_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_24_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_24_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_24_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_24_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_24_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_24_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_24_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_24_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_24_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_24_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_24_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_24_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_24_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_24_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_24_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_24_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_24_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_24_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_24_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_24_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_24_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_24_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_24_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_24_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_24_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_24_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_24_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_24_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_24_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_24_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_24_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_24_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_24_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_24_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_24_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_24_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_24_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_24_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_24_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_24_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_24_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_24_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_24_io_o_age),
    .io_i_ROB_first_entry(reservation_station_24_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_25 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_25_clock),
    .reset(reservation_station_25_reset),
    .io_o_valid(reservation_station_25_io_o_valid),
    .io_o_ready_to_issue(reservation_station_25_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_25_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_25_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_25_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_25_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_25_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_25_io_i_exception),
    .io_i_write_slot(reservation_station_25_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_25_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_25_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_25_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_25_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_25_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_25_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_25_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_25_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_25_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_25_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_25_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_25_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_25_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_25_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_25_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_25_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_25_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_25_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_25_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_25_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_25_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_25_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_25_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_25_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_25_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_25_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_25_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_25_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_25_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_25_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_25_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_25_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_25_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_25_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_25_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_25_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_25_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_25_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_25_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_25_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_25_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_25_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_25_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_25_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_25_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_25_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_25_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_25_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_25_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_25_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_25_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_25_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_25_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_25_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_25_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_25_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_25_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_25_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_25_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_25_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_25_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_25_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_25_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_25_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_25_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_25_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_25_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_25_io_o_age),
    .io_i_ROB_first_entry(reservation_station_25_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_26 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_26_clock),
    .reset(reservation_station_26_reset),
    .io_o_valid(reservation_station_26_io_o_valid),
    .io_o_ready_to_issue(reservation_station_26_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_26_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_26_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_26_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_26_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_26_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_26_io_i_exception),
    .io_i_write_slot(reservation_station_26_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_26_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_26_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_26_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_26_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_26_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_26_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_26_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_26_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_26_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_26_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_26_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_26_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_26_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_26_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_26_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_26_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_26_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_26_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_26_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_26_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_26_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_26_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_26_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_26_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_26_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_26_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_26_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_26_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_26_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_26_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_26_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_26_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_26_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_26_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_26_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_26_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_26_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_26_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_26_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_26_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_26_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_26_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_26_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_26_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_26_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_26_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_26_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_26_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_26_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_26_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_26_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_26_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_26_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_26_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_26_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_26_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_26_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_26_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_26_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_26_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_26_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_26_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_26_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_26_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_26_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_26_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_26_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_26_io_o_age),
    .io_i_ROB_first_entry(reservation_station_26_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_27 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_27_clock),
    .reset(reservation_station_27_reset),
    .io_o_valid(reservation_station_27_io_o_valid),
    .io_o_ready_to_issue(reservation_station_27_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_27_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_27_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_27_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_27_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_27_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_27_io_i_exception),
    .io_i_write_slot(reservation_station_27_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_27_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_27_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_27_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_27_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_27_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_27_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_27_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_27_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_27_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_27_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_27_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_27_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_27_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_27_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_27_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_27_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_27_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_27_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_27_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_27_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_27_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_27_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_27_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_27_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_27_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_27_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_27_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_27_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_27_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_27_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_27_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_27_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_27_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_27_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_27_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_27_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_27_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_27_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_27_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_27_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_27_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_27_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_27_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_27_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_27_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_27_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_27_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_27_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_27_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_27_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_27_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_27_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_27_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_27_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_27_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_27_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_27_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_27_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_27_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_27_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_27_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_27_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_27_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_27_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_27_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_27_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_27_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_27_io_o_age),
    .io_i_ROB_first_entry(reservation_station_27_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_28 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_28_clock),
    .reset(reservation_station_28_reset),
    .io_o_valid(reservation_station_28_io_o_valid),
    .io_o_ready_to_issue(reservation_station_28_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_28_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_28_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_28_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_28_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_28_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_28_io_i_exception),
    .io_i_write_slot(reservation_station_28_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_28_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_28_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_28_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_28_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_28_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_28_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_28_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_28_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_28_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_28_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_28_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_28_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_28_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_28_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_28_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_28_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_28_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_28_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_28_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_28_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_28_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_28_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_28_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_28_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_28_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_28_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_28_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_28_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_28_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_28_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_28_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_28_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_28_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_28_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_28_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_28_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_28_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_28_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_28_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_28_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_28_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_28_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_28_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_28_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_28_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_28_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_28_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_28_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_28_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_28_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_28_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_28_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_28_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_28_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_28_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_28_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_28_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_28_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_28_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_28_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_28_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_28_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_28_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_28_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_28_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_28_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_28_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_28_io_o_age),
    .io_i_ROB_first_entry(reservation_station_28_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_29 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_29_clock),
    .reset(reservation_station_29_reset),
    .io_o_valid(reservation_station_29_io_o_valid),
    .io_o_ready_to_issue(reservation_station_29_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_29_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_29_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_29_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_29_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_29_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_29_io_i_exception),
    .io_i_write_slot(reservation_station_29_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_29_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_29_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_29_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_29_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_29_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_29_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_29_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_29_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_29_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_29_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_29_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_29_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_29_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_29_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_29_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_29_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_29_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_29_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_29_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_29_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_29_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_29_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_29_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_29_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_29_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_29_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_29_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_29_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_29_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_29_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_29_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_29_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_29_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_29_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_29_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_29_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_29_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_29_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_29_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_29_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_29_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_29_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_29_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_29_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_29_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_29_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_29_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_29_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_29_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_29_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_29_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_29_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_29_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_29_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_29_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_29_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_29_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_29_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_29_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_29_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_29_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_29_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_29_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_29_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_29_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_29_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_29_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_29_io_o_age),
    .io_i_ROB_first_entry(reservation_station_29_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_30 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_30_clock),
    .reset(reservation_station_30_reset),
    .io_o_valid(reservation_station_30_io_o_valid),
    .io_o_ready_to_issue(reservation_station_30_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_30_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_30_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_30_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_30_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_30_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_30_io_i_exception),
    .io_i_write_slot(reservation_station_30_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_30_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_30_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_30_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_30_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_30_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_30_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_30_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_30_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_30_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_30_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_30_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_30_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_30_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_30_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_30_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_30_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_30_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_30_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_30_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_30_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_30_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_30_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_30_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_30_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_30_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_30_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_30_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_30_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_30_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_30_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_30_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_30_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_30_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_30_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_30_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_30_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_30_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_30_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_30_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_30_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_30_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_30_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_30_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_30_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_30_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_30_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_30_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_30_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_30_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_30_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_30_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_30_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_30_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_30_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_30_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_30_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_30_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_30_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_30_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_30_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_30_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_30_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_30_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_30_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_30_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_30_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_30_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_30_io_o_age),
    .io_i_ROB_first_entry(reservation_station_30_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_31 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_31_clock),
    .reset(reservation_station_31_reset),
    .io_o_valid(reservation_station_31_io_o_valid),
    .io_o_ready_to_issue(reservation_station_31_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_31_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_31_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_31_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_31_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_31_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_31_io_i_exception),
    .io_i_write_slot(reservation_station_31_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_31_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_31_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_31_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_31_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_31_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_31_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_31_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_31_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_31_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_31_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_31_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_31_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_31_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_31_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_31_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_31_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_31_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_31_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_31_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_31_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_31_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_31_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_31_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_31_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_31_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_31_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_31_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_31_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_31_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_31_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_31_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_31_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_31_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_31_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_31_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_31_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_31_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_31_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_31_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_31_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_31_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_31_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_31_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_31_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_31_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_31_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_31_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_31_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_31_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_31_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_31_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_31_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_31_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_31_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_31_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_31_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_31_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_31_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_31_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_31_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_31_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_31_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_31_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_31_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_31_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_31_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_31_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_31_io_o_age),
    .io_i_ROB_first_entry(reservation_station_31_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_32 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_32_clock),
    .reset(reservation_station_32_reset),
    .io_o_valid(reservation_station_32_io_o_valid),
    .io_o_ready_to_issue(reservation_station_32_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_32_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_32_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_32_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_32_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_32_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_32_io_i_exception),
    .io_i_write_slot(reservation_station_32_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_32_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_32_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_32_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_32_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_32_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_32_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_32_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_32_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_32_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_32_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_32_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_32_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_32_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_32_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_32_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_32_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_32_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_32_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_32_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_32_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_32_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_32_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_32_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_32_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_32_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_32_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_32_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_32_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_32_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_32_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_32_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_32_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_32_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_32_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_32_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_32_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_32_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_32_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_32_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_32_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_32_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_32_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_32_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_32_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_32_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_32_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_32_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_32_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_32_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_32_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_32_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_32_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_32_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_32_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_32_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_32_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_32_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_32_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_32_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_32_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_32_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_32_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_32_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_32_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_32_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_32_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_32_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_32_io_o_age),
    .io_i_ROB_first_entry(reservation_station_32_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_33 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_33_clock),
    .reset(reservation_station_33_reset),
    .io_o_valid(reservation_station_33_io_o_valid),
    .io_o_ready_to_issue(reservation_station_33_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_33_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_33_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_33_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_33_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_33_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_33_io_i_exception),
    .io_i_write_slot(reservation_station_33_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_33_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_33_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_33_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_33_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_33_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_33_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_33_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_33_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_33_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_33_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_33_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_33_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_33_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_33_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_33_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_33_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_33_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_33_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_33_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_33_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_33_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_33_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_33_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_33_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_33_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_33_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_33_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_33_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_33_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_33_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_33_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_33_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_33_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_33_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_33_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_33_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_33_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_33_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_33_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_33_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_33_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_33_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_33_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_33_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_33_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_33_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_33_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_33_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_33_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_33_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_33_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_33_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_33_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_33_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_33_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_33_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_33_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_33_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_33_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_33_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_33_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_33_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_33_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_33_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_33_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_33_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_33_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_33_io_o_age),
    .io_i_ROB_first_entry(reservation_station_33_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_34 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_34_clock),
    .reset(reservation_station_34_reset),
    .io_o_valid(reservation_station_34_io_o_valid),
    .io_o_ready_to_issue(reservation_station_34_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_34_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_34_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_34_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_34_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_34_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_34_io_i_exception),
    .io_i_write_slot(reservation_station_34_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_34_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_34_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_34_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_34_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_34_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_34_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_34_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_34_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_34_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_34_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_34_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_34_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_34_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_34_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_34_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_34_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_34_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_34_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_34_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_34_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_34_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_34_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_34_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_34_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_34_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_34_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_34_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_34_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_34_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_34_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_34_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_34_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_34_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_34_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_34_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_34_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_34_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_34_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_34_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_34_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_34_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_34_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_34_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_34_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_34_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_34_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_34_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_34_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_34_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_34_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_34_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_34_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_34_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_34_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_34_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_34_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_34_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_34_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_34_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_34_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_34_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_34_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_34_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_34_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_34_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_34_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_34_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_34_io_o_age),
    .io_i_ROB_first_entry(reservation_station_34_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_35 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_35_clock),
    .reset(reservation_station_35_reset),
    .io_o_valid(reservation_station_35_io_o_valid),
    .io_o_ready_to_issue(reservation_station_35_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_35_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_35_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_35_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_35_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_35_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_35_io_i_exception),
    .io_i_write_slot(reservation_station_35_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_35_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_35_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_35_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_35_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_35_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_35_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_35_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_35_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_35_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_35_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_35_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_35_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_35_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_35_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_35_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_35_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_35_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_35_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_35_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_35_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_35_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_35_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_35_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_35_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_35_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_35_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_35_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_35_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_35_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_35_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_35_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_35_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_35_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_35_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_35_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_35_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_35_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_35_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_35_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_35_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_35_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_35_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_35_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_35_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_35_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_35_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_35_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_35_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_35_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_35_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_35_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_35_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_35_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_35_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_35_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_35_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_35_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_35_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_35_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_35_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_35_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_35_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_35_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_35_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_35_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_35_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_35_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_35_io_o_age),
    .io_i_ROB_first_entry(reservation_station_35_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_36 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_36_clock),
    .reset(reservation_station_36_reset),
    .io_o_valid(reservation_station_36_io_o_valid),
    .io_o_ready_to_issue(reservation_station_36_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_36_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_36_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_36_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_36_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_36_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_36_io_i_exception),
    .io_i_write_slot(reservation_station_36_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_36_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_36_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_36_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_36_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_36_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_36_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_36_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_36_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_36_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_36_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_36_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_36_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_36_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_36_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_36_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_36_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_36_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_36_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_36_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_36_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_36_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_36_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_36_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_36_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_36_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_36_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_36_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_36_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_36_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_36_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_36_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_36_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_36_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_36_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_36_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_36_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_36_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_36_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_36_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_36_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_36_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_36_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_36_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_36_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_36_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_36_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_36_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_36_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_36_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_36_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_36_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_36_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_36_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_36_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_36_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_36_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_36_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_36_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_36_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_36_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_36_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_36_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_36_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_36_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_36_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_36_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_36_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_36_io_o_age),
    .io_i_ROB_first_entry(reservation_station_36_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_37 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_37_clock),
    .reset(reservation_station_37_reset),
    .io_o_valid(reservation_station_37_io_o_valid),
    .io_o_ready_to_issue(reservation_station_37_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_37_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_37_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_37_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_37_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_37_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_37_io_i_exception),
    .io_i_write_slot(reservation_station_37_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_37_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_37_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_37_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_37_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_37_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_37_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_37_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_37_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_37_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_37_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_37_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_37_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_37_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_37_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_37_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_37_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_37_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_37_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_37_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_37_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_37_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_37_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_37_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_37_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_37_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_37_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_37_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_37_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_37_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_37_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_37_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_37_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_37_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_37_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_37_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_37_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_37_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_37_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_37_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_37_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_37_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_37_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_37_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_37_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_37_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_37_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_37_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_37_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_37_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_37_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_37_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_37_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_37_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_37_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_37_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_37_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_37_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_37_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_37_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_37_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_37_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_37_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_37_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_37_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_37_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_37_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_37_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_37_io_o_age),
    .io_i_ROB_first_entry(reservation_station_37_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_38 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_38_clock),
    .reset(reservation_station_38_reset),
    .io_o_valid(reservation_station_38_io_o_valid),
    .io_o_ready_to_issue(reservation_station_38_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_38_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_38_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_38_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_38_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_38_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_38_io_i_exception),
    .io_i_write_slot(reservation_station_38_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_38_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_38_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_38_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_38_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_38_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_38_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_38_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_38_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_38_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_38_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_38_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_38_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_38_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_38_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_38_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_38_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_38_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_38_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_38_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_38_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_38_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_38_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_38_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_38_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_38_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_38_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_38_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_38_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_38_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_38_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_38_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_38_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_38_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_38_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_38_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_38_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_38_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_38_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_38_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_38_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_38_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_38_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_38_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_38_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_38_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_38_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_38_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_38_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_38_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_38_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_38_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_38_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_38_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_38_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_38_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_38_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_38_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_38_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_38_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_38_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_38_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_38_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_38_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_38_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_38_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_38_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_38_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_38_io_o_age),
    .io_i_ROB_first_entry(reservation_station_38_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_39 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_39_clock),
    .reset(reservation_station_39_reset),
    .io_o_valid(reservation_station_39_io_o_valid),
    .io_o_ready_to_issue(reservation_station_39_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_39_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_39_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_39_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_39_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_39_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_39_io_i_exception),
    .io_i_write_slot(reservation_station_39_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_39_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_39_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_39_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_39_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_39_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_39_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_39_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_39_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_39_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_39_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_39_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_39_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_39_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_39_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_39_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_39_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_39_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_39_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_39_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_39_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_39_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_39_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_39_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_39_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_39_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_39_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_39_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_39_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_39_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_39_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_39_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_39_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_39_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_39_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_39_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_39_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_39_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_39_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_39_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_39_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_39_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_39_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_39_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_39_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_39_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_39_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_39_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_39_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_39_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_39_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_39_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_39_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_39_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_39_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_39_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_39_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_39_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_39_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_39_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_39_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_39_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_39_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_39_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_39_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_39_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_39_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_39_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_39_io_o_age),
    .io_i_ROB_first_entry(reservation_station_39_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_40 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_40_clock),
    .reset(reservation_station_40_reset),
    .io_o_valid(reservation_station_40_io_o_valid),
    .io_o_ready_to_issue(reservation_station_40_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_40_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_40_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_40_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_40_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_40_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_40_io_i_exception),
    .io_i_write_slot(reservation_station_40_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_40_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_40_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_40_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_40_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_40_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_40_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_40_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_40_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_40_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_40_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_40_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_40_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_40_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_40_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_40_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_40_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_40_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_40_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_40_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_40_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_40_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_40_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_40_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_40_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_40_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_40_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_40_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_40_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_40_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_40_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_40_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_40_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_40_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_40_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_40_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_40_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_40_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_40_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_40_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_40_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_40_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_40_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_40_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_40_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_40_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_40_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_40_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_40_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_40_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_40_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_40_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_40_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_40_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_40_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_40_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_40_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_40_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_40_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_40_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_40_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_40_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_40_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_40_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_40_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_40_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_40_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_40_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_40_io_o_age),
    .io_i_ROB_first_entry(reservation_station_40_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_41 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_41_clock),
    .reset(reservation_station_41_reset),
    .io_o_valid(reservation_station_41_io_o_valid),
    .io_o_ready_to_issue(reservation_station_41_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_41_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_41_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_41_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_41_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_41_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_41_io_i_exception),
    .io_i_write_slot(reservation_station_41_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_41_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_41_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_41_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_41_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_41_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_41_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_41_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_41_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_41_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_41_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_41_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_41_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_41_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_41_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_41_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_41_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_41_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_41_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_41_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_41_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_41_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_41_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_41_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_41_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_41_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_41_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_41_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_41_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_41_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_41_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_41_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_41_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_41_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_41_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_41_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_41_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_41_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_41_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_41_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_41_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_41_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_41_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_41_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_41_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_41_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_41_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_41_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_41_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_41_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_41_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_41_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_41_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_41_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_41_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_41_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_41_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_41_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_41_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_41_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_41_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_41_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_41_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_41_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_41_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_41_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_41_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_41_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_41_io_o_age),
    .io_i_ROB_first_entry(reservation_station_41_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_42 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_42_clock),
    .reset(reservation_station_42_reset),
    .io_o_valid(reservation_station_42_io_o_valid),
    .io_o_ready_to_issue(reservation_station_42_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_42_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_42_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_42_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_42_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_42_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_42_io_i_exception),
    .io_i_write_slot(reservation_station_42_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_42_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_42_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_42_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_42_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_42_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_42_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_42_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_42_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_42_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_42_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_42_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_42_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_42_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_42_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_42_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_42_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_42_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_42_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_42_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_42_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_42_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_42_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_42_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_42_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_42_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_42_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_42_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_42_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_42_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_42_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_42_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_42_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_42_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_42_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_42_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_42_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_42_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_42_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_42_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_42_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_42_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_42_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_42_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_42_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_42_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_42_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_42_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_42_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_42_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_42_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_42_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_42_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_42_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_42_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_42_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_42_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_42_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_42_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_42_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_42_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_42_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_42_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_42_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_42_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_42_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_42_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_42_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_42_io_o_age),
    .io_i_ROB_first_entry(reservation_station_42_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_43 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_43_clock),
    .reset(reservation_station_43_reset),
    .io_o_valid(reservation_station_43_io_o_valid),
    .io_o_ready_to_issue(reservation_station_43_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_43_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_43_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_43_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_43_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_43_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_43_io_i_exception),
    .io_i_write_slot(reservation_station_43_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_43_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_43_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_43_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_43_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_43_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_43_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_43_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_43_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_43_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_43_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_43_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_43_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_43_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_43_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_43_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_43_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_43_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_43_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_43_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_43_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_43_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_43_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_43_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_43_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_43_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_43_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_43_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_43_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_43_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_43_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_43_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_43_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_43_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_43_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_43_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_43_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_43_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_43_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_43_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_43_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_43_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_43_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_43_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_43_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_43_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_43_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_43_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_43_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_43_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_43_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_43_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_43_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_43_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_43_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_43_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_43_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_43_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_43_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_43_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_43_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_43_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_43_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_43_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_43_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_43_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_43_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_43_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_43_io_o_age),
    .io_i_ROB_first_entry(reservation_station_43_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_44 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_44_clock),
    .reset(reservation_station_44_reset),
    .io_o_valid(reservation_station_44_io_o_valid),
    .io_o_ready_to_issue(reservation_station_44_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_44_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_44_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_44_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_44_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_44_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_44_io_i_exception),
    .io_i_write_slot(reservation_station_44_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_44_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_44_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_44_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_44_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_44_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_44_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_44_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_44_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_44_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_44_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_44_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_44_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_44_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_44_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_44_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_44_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_44_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_44_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_44_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_44_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_44_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_44_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_44_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_44_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_44_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_44_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_44_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_44_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_44_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_44_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_44_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_44_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_44_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_44_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_44_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_44_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_44_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_44_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_44_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_44_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_44_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_44_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_44_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_44_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_44_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_44_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_44_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_44_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_44_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_44_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_44_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_44_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_44_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_44_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_44_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_44_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_44_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_44_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_44_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_44_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_44_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_44_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_44_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_44_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_44_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_44_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_44_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_44_io_o_age),
    .io_i_ROB_first_entry(reservation_station_44_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_45 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_45_clock),
    .reset(reservation_station_45_reset),
    .io_o_valid(reservation_station_45_io_o_valid),
    .io_o_ready_to_issue(reservation_station_45_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_45_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_45_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_45_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_45_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_45_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_45_io_i_exception),
    .io_i_write_slot(reservation_station_45_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_45_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_45_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_45_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_45_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_45_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_45_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_45_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_45_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_45_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_45_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_45_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_45_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_45_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_45_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_45_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_45_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_45_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_45_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_45_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_45_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_45_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_45_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_45_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_45_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_45_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_45_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_45_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_45_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_45_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_45_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_45_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_45_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_45_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_45_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_45_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_45_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_45_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_45_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_45_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_45_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_45_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_45_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_45_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_45_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_45_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_45_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_45_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_45_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_45_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_45_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_45_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_45_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_45_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_45_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_45_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_45_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_45_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_45_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_45_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_45_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_45_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_45_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_45_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_45_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_45_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_45_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_45_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_45_io_o_age),
    .io_i_ROB_first_entry(reservation_station_45_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_46 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_46_clock),
    .reset(reservation_station_46_reset),
    .io_o_valid(reservation_station_46_io_o_valid),
    .io_o_ready_to_issue(reservation_station_46_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_46_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_46_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_46_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_46_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_46_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_46_io_i_exception),
    .io_i_write_slot(reservation_station_46_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_46_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_46_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_46_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_46_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_46_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_46_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_46_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_46_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_46_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_46_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_46_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_46_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_46_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_46_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_46_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_46_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_46_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_46_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_46_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_46_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_46_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_46_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_46_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_46_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_46_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_46_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_46_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_46_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_46_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_46_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_46_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_46_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_46_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_46_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_46_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_46_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_46_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_46_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_46_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_46_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_46_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_46_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_46_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_46_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_46_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_46_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_46_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_46_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_46_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_46_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_46_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_46_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_46_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_46_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_46_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_46_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_46_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_46_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_46_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_46_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_46_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_46_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_46_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_46_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_46_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_46_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_46_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_46_io_o_age),
    .io_i_ROB_first_entry(reservation_station_46_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_47 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_47_clock),
    .reset(reservation_station_47_reset),
    .io_o_valid(reservation_station_47_io_o_valid),
    .io_o_ready_to_issue(reservation_station_47_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_47_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_47_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_47_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_47_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_47_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_47_io_i_exception),
    .io_i_write_slot(reservation_station_47_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_47_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_47_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_47_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_47_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_47_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_47_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_47_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_47_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_47_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_47_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_47_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_47_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_47_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_47_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_47_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_47_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_47_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_47_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_47_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_47_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_47_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_47_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_47_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_47_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_47_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_47_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_47_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_47_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_47_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_47_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_47_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_47_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_47_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_47_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_47_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_47_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_47_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_47_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_47_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_47_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_47_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_47_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_47_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_47_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_47_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_47_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_47_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_47_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_47_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_47_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_47_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_47_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_47_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_47_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_47_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_47_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_47_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_47_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_47_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_47_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_47_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_47_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_47_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_47_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_47_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_47_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_47_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_47_io_o_age),
    .io_i_ROB_first_entry(reservation_station_47_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_48 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_48_clock),
    .reset(reservation_station_48_reset),
    .io_o_valid(reservation_station_48_io_o_valid),
    .io_o_ready_to_issue(reservation_station_48_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_48_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_48_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_48_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_48_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_48_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_48_io_i_exception),
    .io_i_write_slot(reservation_station_48_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_48_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_48_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_48_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_48_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_48_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_48_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_48_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_48_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_48_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_48_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_48_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_48_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_48_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_48_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_48_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_48_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_48_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_48_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_48_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_48_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_48_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_48_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_48_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_48_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_48_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_48_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_48_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_48_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_48_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_48_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_48_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_48_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_48_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_48_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_48_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_48_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_48_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_48_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_48_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_48_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_48_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_48_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_48_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_48_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_48_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_48_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_48_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_48_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_48_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_48_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_48_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_48_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_48_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_48_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_48_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_48_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_48_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_48_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_48_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_48_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_48_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_48_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_48_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_48_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_48_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_48_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_48_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_48_io_o_age),
    .io_i_ROB_first_entry(reservation_station_48_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_49 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_49_clock),
    .reset(reservation_station_49_reset),
    .io_o_valid(reservation_station_49_io_o_valid),
    .io_o_ready_to_issue(reservation_station_49_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_49_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_49_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_49_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_49_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_49_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_49_io_i_exception),
    .io_i_write_slot(reservation_station_49_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_49_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_49_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_49_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_49_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_49_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_49_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_49_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_49_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_49_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_49_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_49_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_49_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_49_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_49_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_49_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_49_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_49_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_49_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_49_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_49_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_49_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_49_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_49_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_49_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_49_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_49_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_49_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_49_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_49_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_49_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_49_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_49_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_49_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_49_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_49_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_49_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_49_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_49_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_49_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_49_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_49_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_49_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_49_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_49_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_49_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_49_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_49_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_49_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_49_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_49_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_49_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_49_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_49_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_49_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_49_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_49_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_49_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_49_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_49_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_49_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_49_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_49_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_49_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_49_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_49_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_49_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_49_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_49_io_o_age),
    .io_i_ROB_first_entry(reservation_station_49_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_50 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_50_clock),
    .reset(reservation_station_50_reset),
    .io_o_valid(reservation_station_50_io_o_valid),
    .io_o_ready_to_issue(reservation_station_50_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_50_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_50_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_50_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_50_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_50_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_50_io_i_exception),
    .io_i_write_slot(reservation_station_50_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_50_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_50_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_50_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_50_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_50_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_50_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_50_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_50_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_50_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_50_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_50_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_50_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_50_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_50_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_50_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_50_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_50_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_50_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_50_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_50_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_50_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_50_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_50_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_50_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_50_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_50_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_50_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_50_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_50_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_50_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_50_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_50_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_50_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_50_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_50_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_50_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_50_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_50_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_50_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_50_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_50_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_50_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_50_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_50_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_50_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_50_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_50_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_50_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_50_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_50_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_50_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_50_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_50_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_50_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_50_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_50_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_50_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_50_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_50_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_50_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_50_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_50_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_50_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_50_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_50_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_50_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_50_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_50_io_o_age),
    .io_i_ROB_first_entry(reservation_station_50_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_51 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_51_clock),
    .reset(reservation_station_51_reset),
    .io_o_valid(reservation_station_51_io_o_valid),
    .io_o_ready_to_issue(reservation_station_51_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_51_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_51_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_51_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_51_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_51_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_51_io_i_exception),
    .io_i_write_slot(reservation_station_51_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_51_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_51_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_51_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_51_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_51_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_51_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_51_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_51_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_51_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_51_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_51_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_51_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_51_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_51_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_51_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_51_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_51_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_51_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_51_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_51_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_51_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_51_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_51_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_51_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_51_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_51_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_51_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_51_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_51_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_51_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_51_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_51_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_51_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_51_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_51_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_51_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_51_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_51_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_51_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_51_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_51_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_51_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_51_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_51_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_51_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_51_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_51_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_51_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_51_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_51_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_51_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_51_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_51_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_51_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_51_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_51_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_51_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_51_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_51_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_51_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_51_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_51_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_51_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_51_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_51_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_51_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_51_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_51_io_o_age),
    .io_i_ROB_first_entry(reservation_station_51_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_52 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_52_clock),
    .reset(reservation_station_52_reset),
    .io_o_valid(reservation_station_52_io_o_valid),
    .io_o_ready_to_issue(reservation_station_52_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_52_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_52_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_52_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_52_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_52_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_52_io_i_exception),
    .io_i_write_slot(reservation_station_52_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_52_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_52_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_52_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_52_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_52_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_52_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_52_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_52_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_52_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_52_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_52_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_52_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_52_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_52_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_52_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_52_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_52_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_52_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_52_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_52_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_52_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_52_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_52_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_52_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_52_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_52_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_52_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_52_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_52_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_52_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_52_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_52_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_52_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_52_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_52_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_52_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_52_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_52_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_52_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_52_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_52_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_52_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_52_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_52_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_52_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_52_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_52_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_52_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_52_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_52_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_52_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_52_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_52_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_52_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_52_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_52_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_52_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_52_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_52_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_52_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_52_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_52_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_52_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_52_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_52_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_52_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_52_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_52_io_o_age),
    .io_i_ROB_first_entry(reservation_station_52_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_53 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_53_clock),
    .reset(reservation_station_53_reset),
    .io_o_valid(reservation_station_53_io_o_valid),
    .io_o_ready_to_issue(reservation_station_53_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_53_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_53_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_53_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_53_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_53_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_53_io_i_exception),
    .io_i_write_slot(reservation_station_53_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_53_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_53_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_53_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_53_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_53_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_53_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_53_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_53_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_53_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_53_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_53_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_53_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_53_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_53_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_53_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_53_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_53_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_53_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_53_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_53_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_53_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_53_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_53_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_53_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_53_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_53_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_53_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_53_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_53_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_53_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_53_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_53_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_53_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_53_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_53_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_53_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_53_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_53_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_53_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_53_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_53_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_53_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_53_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_53_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_53_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_53_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_53_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_53_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_53_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_53_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_53_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_53_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_53_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_53_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_53_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_53_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_53_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_53_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_53_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_53_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_53_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_53_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_53_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_53_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_53_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_53_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_53_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_53_io_o_age),
    .io_i_ROB_first_entry(reservation_station_53_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_54 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_54_clock),
    .reset(reservation_station_54_reset),
    .io_o_valid(reservation_station_54_io_o_valid),
    .io_o_ready_to_issue(reservation_station_54_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_54_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_54_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_54_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_54_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_54_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_54_io_i_exception),
    .io_i_write_slot(reservation_station_54_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_54_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_54_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_54_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_54_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_54_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_54_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_54_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_54_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_54_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_54_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_54_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_54_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_54_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_54_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_54_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_54_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_54_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_54_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_54_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_54_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_54_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_54_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_54_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_54_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_54_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_54_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_54_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_54_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_54_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_54_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_54_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_54_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_54_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_54_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_54_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_54_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_54_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_54_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_54_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_54_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_54_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_54_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_54_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_54_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_54_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_54_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_54_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_54_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_54_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_54_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_54_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_54_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_54_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_54_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_54_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_54_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_54_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_54_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_54_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_54_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_54_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_54_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_54_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_54_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_54_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_54_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_54_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_54_io_o_age),
    .io_i_ROB_first_entry(reservation_station_54_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_55 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_55_clock),
    .reset(reservation_station_55_reset),
    .io_o_valid(reservation_station_55_io_o_valid),
    .io_o_ready_to_issue(reservation_station_55_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_55_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_55_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_55_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_55_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_55_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_55_io_i_exception),
    .io_i_write_slot(reservation_station_55_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_55_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_55_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_55_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_55_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_55_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_55_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_55_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_55_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_55_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_55_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_55_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_55_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_55_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_55_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_55_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_55_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_55_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_55_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_55_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_55_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_55_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_55_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_55_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_55_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_55_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_55_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_55_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_55_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_55_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_55_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_55_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_55_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_55_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_55_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_55_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_55_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_55_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_55_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_55_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_55_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_55_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_55_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_55_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_55_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_55_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_55_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_55_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_55_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_55_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_55_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_55_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_55_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_55_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_55_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_55_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_55_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_55_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_55_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_55_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_55_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_55_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_55_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_55_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_55_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_55_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_55_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_55_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_55_io_o_age),
    .io_i_ROB_first_entry(reservation_station_55_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_56 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_56_clock),
    .reset(reservation_station_56_reset),
    .io_o_valid(reservation_station_56_io_o_valid),
    .io_o_ready_to_issue(reservation_station_56_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_56_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_56_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_56_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_56_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_56_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_56_io_i_exception),
    .io_i_write_slot(reservation_station_56_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_56_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_56_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_56_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_56_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_56_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_56_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_56_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_56_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_56_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_56_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_56_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_56_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_56_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_56_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_56_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_56_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_56_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_56_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_56_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_56_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_56_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_56_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_56_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_56_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_56_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_56_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_56_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_56_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_56_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_56_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_56_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_56_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_56_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_56_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_56_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_56_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_56_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_56_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_56_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_56_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_56_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_56_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_56_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_56_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_56_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_56_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_56_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_56_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_56_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_56_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_56_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_56_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_56_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_56_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_56_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_56_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_56_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_56_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_56_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_56_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_56_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_56_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_56_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_56_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_56_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_56_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_56_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_56_io_o_age),
    .io_i_ROB_first_entry(reservation_station_56_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_57 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_57_clock),
    .reset(reservation_station_57_reset),
    .io_o_valid(reservation_station_57_io_o_valid),
    .io_o_ready_to_issue(reservation_station_57_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_57_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_57_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_57_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_57_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_57_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_57_io_i_exception),
    .io_i_write_slot(reservation_station_57_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_57_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_57_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_57_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_57_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_57_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_57_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_57_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_57_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_57_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_57_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_57_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_57_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_57_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_57_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_57_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_57_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_57_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_57_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_57_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_57_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_57_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_57_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_57_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_57_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_57_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_57_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_57_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_57_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_57_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_57_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_57_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_57_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_57_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_57_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_57_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_57_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_57_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_57_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_57_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_57_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_57_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_57_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_57_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_57_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_57_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_57_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_57_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_57_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_57_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_57_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_57_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_57_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_57_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_57_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_57_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_57_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_57_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_57_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_57_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_57_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_57_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_57_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_57_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_57_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_57_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_57_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_57_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_57_io_o_age),
    .io_i_ROB_first_entry(reservation_station_57_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_58 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_58_clock),
    .reset(reservation_station_58_reset),
    .io_o_valid(reservation_station_58_io_o_valid),
    .io_o_ready_to_issue(reservation_station_58_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_58_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_58_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_58_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_58_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_58_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_58_io_i_exception),
    .io_i_write_slot(reservation_station_58_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_58_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_58_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_58_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_58_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_58_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_58_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_58_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_58_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_58_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_58_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_58_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_58_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_58_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_58_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_58_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_58_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_58_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_58_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_58_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_58_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_58_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_58_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_58_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_58_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_58_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_58_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_58_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_58_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_58_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_58_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_58_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_58_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_58_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_58_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_58_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_58_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_58_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_58_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_58_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_58_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_58_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_58_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_58_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_58_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_58_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_58_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_58_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_58_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_58_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_58_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_58_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_58_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_58_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_58_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_58_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_58_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_58_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_58_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_58_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_58_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_58_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_58_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_58_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_58_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_58_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_58_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_58_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_58_io_o_age),
    .io_i_ROB_first_entry(reservation_station_58_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_59 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_59_clock),
    .reset(reservation_station_59_reset),
    .io_o_valid(reservation_station_59_io_o_valid),
    .io_o_ready_to_issue(reservation_station_59_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_59_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_59_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_59_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_59_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_59_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_59_io_i_exception),
    .io_i_write_slot(reservation_station_59_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_59_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_59_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_59_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_59_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_59_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_59_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_59_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_59_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_59_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_59_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_59_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_59_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_59_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_59_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_59_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_59_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_59_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_59_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_59_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_59_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_59_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_59_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_59_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_59_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_59_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_59_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_59_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_59_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_59_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_59_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_59_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_59_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_59_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_59_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_59_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_59_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_59_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_59_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_59_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_59_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_59_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_59_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_59_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_59_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_59_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_59_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_59_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_59_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_59_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_59_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_59_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_59_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_59_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_59_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_59_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_59_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_59_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_59_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_59_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_59_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_59_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_59_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_59_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_59_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_59_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_59_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_59_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_59_io_o_age),
    .io_i_ROB_first_entry(reservation_station_59_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_60 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_60_clock),
    .reset(reservation_station_60_reset),
    .io_o_valid(reservation_station_60_io_o_valid),
    .io_o_ready_to_issue(reservation_station_60_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_60_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_60_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_60_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_60_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_60_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_60_io_i_exception),
    .io_i_write_slot(reservation_station_60_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_60_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_60_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_60_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_60_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_60_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_60_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_60_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_60_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_60_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_60_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_60_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_60_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_60_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_60_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_60_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_60_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_60_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_60_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_60_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_60_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_60_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_60_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_60_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_60_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_60_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_60_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_60_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_60_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_60_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_60_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_60_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_60_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_60_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_60_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_60_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_60_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_60_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_60_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_60_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_60_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_60_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_60_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_60_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_60_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_60_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_60_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_60_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_60_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_60_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_60_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_60_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_60_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_60_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_60_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_60_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_60_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_60_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_60_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_60_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_60_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_60_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_60_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_60_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_60_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_60_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_60_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_60_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_60_io_o_age),
    .io_i_ROB_first_entry(reservation_station_60_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_61 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_61_clock),
    .reset(reservation_station_61_reset),
    .io_o_valid(reservation_station_61_io_o_valid),
    .io_o_ready_to_issue(reservation_station_61_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_61_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_61_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_61_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_61_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_61_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_61_io_i_exception),
    .io_i_write_slot(reservation_station_61_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_61_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_61_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_61_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_61_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_61_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_61_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_61_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_61_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_61_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_61_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_61_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_61_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_61_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_61_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_61_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_61_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_61_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_61_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_61_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_61_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_61_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_61_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_61_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_61_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_61_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_61_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_61_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_61_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_61_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_61_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_61_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_61_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_61_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_61_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_61_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_61_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_61_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_61_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_61_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_61_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_61_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_61_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_61_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_61_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_61_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_61_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_61_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_61_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_61_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_61_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_61_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_61_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_61_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_61_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_61_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_61_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_61_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_61_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_61_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_61_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_61_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_61_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_61_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_61_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_61_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_61_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_61_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_61_io_o_age),
    .io_i_ROB_first_entry(reservation_station_61_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_62 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_62_clock),
    .reset(reservation_station_62_reset),
    .io_o_valid(reservation_station_62_io_o_valid),
    .io_o_ready_to_issue(reservation_station_62_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_62_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_62_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_62_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_62_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_62_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_62_io_i_exception),
    .io_i_write_slot(reservation_station_62_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_62_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_62_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_62_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_62_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_62_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_62_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_62_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_62_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_62_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_62_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_62_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_62_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_62_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_62_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_62_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_62_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_62_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_62_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_62_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_62_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_62_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_62_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_62_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_62_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_62_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_62_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_62_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_62_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_62_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_62_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_62_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_62_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_62_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_62_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_62_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_62_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_62_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_62_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_62_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_62_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_62_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_62_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_62_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_62_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_62_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_62_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_62_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_62_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_62_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_62_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_62_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_62_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_62_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_62_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_62_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_62_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_62_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_62_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_62_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_62_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_62_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_62_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_62_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_62_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_62_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_62_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_62_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_62_io_o_age),
    .io_i_ROB_first_entry(reservation_station_62_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_63 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_63_clock),
    .reset(reservation_station_63_reset),
    .io_o_valid(reservation_station_63_io_o_valid),
    .io_o_ready_to_issue(reservation_station_63_io_o_ready_to_issue),
    .io_i_allocated_idx(reservation_station_63_io_i_allocated_idx),
    .io_i_issue_granted(reservation_station_63_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_63_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_63_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_63_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_63_io_i_exception),
    .io_i_write_slot(reservation_station_63_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_63_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_63_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_63_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_63_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_63_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_63_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_63_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_63_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_63_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_63_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_63_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_63_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_63_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_63_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_63_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_63_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_63_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_63_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_63_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_63_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_63_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_63_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_63_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_63_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_63_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_63_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_63_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_63_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_63_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_63_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_63_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_63_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_63_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_63_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_63_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_63_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_63_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_63_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_63_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_63_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_63_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_63_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_63_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_63_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_63_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_63_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_63_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_63_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_63_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_63_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_63_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_63_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_63_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_63_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_63_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_63_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_63_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_63_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_63_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_63_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_63_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_63_io_i_exe_value2),
    .io_i_age_pack_issue_valid_0(reservation_station_63_io_i_age_pack_issue_valid_0),
    .io_i_age_pack_issue_valid_1(reservation_station_63_io_i_age_pack_issue_valid_1),
    .io_i_age_pack_max_age(reservation_station_63_io_i_age_pack_max_age),
    .io_i_age_pack_issued_ages_0(reservation_station_63_io_i_age_pack_issued_ages_0),
    .io_i_age_pack_issued_ages_1(reservation_station_63_io_i_age_pack_issued_ages_1),
    .io_o_age(reservation_station_63_io_o_age),
    .io_i_ROB_first_entry(reservation_station_63_io_i_ROB_first_entry)
  );
  assign io_o_issue_packs_0_valid = issue_num == 2'h1 | issue_num == 2'h2; // @[reservation_station.scala 177:38]
  assign io_o_issue_packs_0_pc = _issue1_func_code_T ? reservation_station_0_io_o_uop_pc : _io_o_issue_packs_0_T_126_pc; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_inst = _issue1_func_code_T ? reservation_station_0_io_o_uop_inst :
    _io_o_issue_packs_0_T_126_inst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_func_code = _issue1_func_code_T ? reservation_station_0_io_o_uop_func_code :
    _io_o_issue_packs_0_T_126_func_code; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_valid = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_126_branch_predict_pack_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_target = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_126_branch_predict_pack_target; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_branch_type = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_126_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_select = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_126_branch_predict_pack_select; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_taken = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_126_branch_predict_pack_taken; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_126_phy_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_stale_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_126_stale_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_126_arch_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_inst_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_126_inst_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_regWen = _issue1_func_code_T ? reservation_station_0_io_o_uop_regWen :
    _io_o_issue_packs_0_T_126_regWen; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src1_valid = _issue1_func_code_T ? reservation_station_0_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_126_src1_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_rs1 = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_126_phy_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_rs1 = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_126_arch_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src2_valid = _issue1_func_code_T ? reservation_station_0_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_126_src2_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_rs2 = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_126_phy_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_rs2 = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_126_arch_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_rob_idx = _issue1_func_code_T ? reservation_station_0_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_126_rob_idx; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_imm = _issue1_func_code_T ? reservation_station_0_io_o_uop_imm :
    _io_o_issue_packs_0_T_126_imm; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src1_value = _issue1_func_code_T ? reservation_station_0_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_126_src1_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src2_value = _issue1_func_code_T ? reservation_station_0_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_126_src2_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_op1_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_126_op1_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_op2_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_126_op2_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_alu_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_126_alu_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_branch_type :
    _io_o_issue_packs_0_T_126_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_mem_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_126_mem_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_valid = issue_num == 2'h2; // @[reservation_station.scala 178:31]
  assign io_o_issue_packs_1_pc = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_pc :
    _io_o_issue_packs_1_T_126_pc; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_inst = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_inst :
    _io_o_issue_packs_1_T_126_inst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_func_code = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_func_code :
    _io_o_issue_packs_1_T_126_func_code; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_valid = _issued_age_pack_issued_ages_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_126_branch_predict_pack_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_target = _issued_age_pack_issued_ages_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_126_branch_predict_pack_target; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_branch_type = _issued_age_pack_issued_ages_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_126_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_select = _issued_age_pack_issued_ages_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_126_branch_predict_pack_select; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_taken = _issued_age_pack_issued_ages_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_126_branch_predict_pack_taken; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_dst = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_126_phy_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_stale_dst = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_126_stale_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_dst = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_126_arch_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_inst_type = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_126_inst_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_regWen = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_regWen :
    _io_o_issue_packs_1_T_126_regWen; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src1_valid = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_126_src1_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_rs1 = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_126_phy_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_rs1 = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_126_arch_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src2_valid = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_126_src2_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_rs2 = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_126_phy_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_rs2 = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_126_arch_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_rob_idx = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_126_rob_idx; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_imm = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_imm :
    _io_o_issue_packs_1_T_126_imm; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src1_value = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_src1_value :
    _io_o_issue_packs_1_T_126_src1_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src2_value = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_src2_value :
    _io_o_issue_packs_1_T_126_src2_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_op1_sel = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_126_op1_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_op2_sel = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_126_op2_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_alu_sel = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_126_alu_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_type = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_branch_type
     : _io_o_issue_packs_1_T_126_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_mem_type = _issued_age_pack_issued_ages_1_T ? reservation_station_0_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_126_mem_type; // @[Mux.scala 101:16]
  assign io_o_full = issued_age_pack_max_age > 8'h3c & _write_num_T_2; // @[reservation_station.scala 233:48]
  assign reservation_station_0_clock = clock;
  assign reservation_station_0_reset = reset;
  assign reservation_station_0_io_i_allocated_idx = write_idx2 == 6'h0; // @[reservation_station.scala 246:65]
  assign reservation_station_0_io_i_issue_granted = (_issue1_func_code_T | _issued_age_pack_issued_ages_1_T) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_0_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_0_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_0_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_0_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_0_io_i_write_slot = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_0_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_0_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_0_io_i_uop_valid = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_pc = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_inst = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_func_code = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_target = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_branch_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_select = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_taken = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_phy_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_stale_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_arch_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_inst_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_regWen = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_src1_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_phy_rs1 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_arch_rs1 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_src2_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_phy_rs2 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_arch_rs2 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_rob_idx = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_imm = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_src1_value = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_src2_value = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_op1_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_op2_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_alu_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_branch_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_uop_mem_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_0_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_0_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_0_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_0_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_0_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_0_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_0_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_0_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_0_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_0_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_1_clock = clock;
  assign reservation_station_1_reset = reset;
  assign reservation_station_1_io_i_allocated_idx = write_idx2 == 6'h1; // @[reservation_station.scala 246:65]
  assign reservation_station_1_io_i_issue_granted = (_issue1_func_code_T_1 | _issued_age_pack_issued_ages_1_T_1) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_1_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_1_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_1_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_1_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_1_io_i_write_slot = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_1_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_1_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_1_io_i_uop_valid = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_pc = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_inst = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_func_code = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_target = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_branch_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_select = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_taken = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_phy_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_stale_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_arch_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_inst_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_regWen = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_src1_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_phy_rs1 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_arch_rs1 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_src2_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_phy_rs2 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_arch_rs2 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_rob_idx = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_imm = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_src1_value = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_src2_value = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_op1_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_op2_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_alu_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_branch_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_uop_mem_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_1_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_1_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_1_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_1_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_1_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_1_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_1_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_1_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_1_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_1_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_2_clock = clock;
  assign reservation_station_2_reset = reset;
  assign reservation_station_2_io_i_allocated_idx = write_idx2 == 6'h2; // @[reservation_station.scala 246:65]
  assign reservation_station_2_io_i_issue_granted = (_issue1_func_code_T_2 | _issued_age_pack_issued_ages_1_T_2) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_2_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_2_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_2_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_2_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_2_io_i_write_slot = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_2_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_2_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_2_io_i_uop_valid = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_pc = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_inst = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_func_code = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_target = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_branch_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_select = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_taken = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_phy_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_stale_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_arch_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_inst_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_regWen = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_src1_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_phy_rs1 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_arch_rs1 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_src2_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_phy_rs2 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_arch_rs2 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_rob_idx = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_imm = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_src1_value = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_src2_value = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_op1_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_op2_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_alu_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_branch_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_uop_mem_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_2_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_2_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_2_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_2_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_2_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_2_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_2_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_2_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_2_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_2_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_3_clock = clock;
  assign reservation_station_3_reset = reset;
  assign reservation_station_3_io_i_allocated_idx = write_idx2 == 6'h3; // @[reservation_station.scala 246:65]
  assign reservation_station_3_io_i_issue_granted = (_issue1_func_code_T_3 | _issued_age_pack_issued_ages_1_T_3) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_3_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_3_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_3_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_3_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_3_io_i_write_slot = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_3_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_3_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_3_io_i_uop_valid = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_pc = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_inst = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_func_code = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_target = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_branch_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_select = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_taken = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_phy_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_stale_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_arch_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_inst_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_regWen = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_src1_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_phy_rs1 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_arch_rs1 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_src2_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_phy_rs2 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_arch_rs2 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_rob_idx = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_imm = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_src1_value = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_src2_value = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_op1_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_op2_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_alu_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_branch_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_uop_mem_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_3_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_3_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_3_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_3_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_3_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_3_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_3_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_3_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_3_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_3_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_4_clock = clock;
  assign reservation_station_4_reset = reset;
  assign reservation_station_4_io_i_allocated_idx = write_idx2 == 6'h4; // @[reservation_station.scala 246:65]
  assign reservation_station_4_io_i_issue_granted = (_issue1_func_code_T_4 | _issued_age_pack_issued_ages_1_T_4) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_4_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_4_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_4_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_4_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_4_io_i_write_slot = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_4_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_4_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_4_io_i_uop_valid = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_pc = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_inst = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_func_code = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_target = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_branch_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_select = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_taken = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_phy_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_stale_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_arch_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_inst_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_regWen = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_src1_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_phy_rs1 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_arch_rs1 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_src2_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_phy_rs2 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_arch_rs2 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_rob_idx = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_imm = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_src1_value = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_src2_value = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_op1_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_op2_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_alu_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_branch_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_uop_mem_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_4_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_4_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_4_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_4_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_4_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_4_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_4_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_4_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_4_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_4_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_5_clock = clock;
  assign reservation_station_5_reset = reset;
  assign reservation_station_5_io_i_allocated_idx = write_idx2 == 6'h5; // @[reservation_station.scala 246:65]
  assign reservation_station_5_io_i_issue_granted = (_issue1_func_code_T_5 | _issued_age_pack_issued_ages_1_T_5) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_5_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_5_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_5_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_5_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_5_io_i_write_slot = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_5_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_5_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_5_io_i_uop_valid = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_pc = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_inst = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_func_code = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_target = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_branch_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_select = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_taken = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_phy_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_stale_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_arch_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_inst_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_regWen = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_src1_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_phy_rs1 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_arch_rs1 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_src2_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_phy_rs2 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_arch_rs2 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_rob_idx = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_imm = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_src1_value = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_src2_value = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_op1_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_op2_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_alu_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_branch_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_uop_mem_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_5_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_5_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_5_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_5_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_5_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_5_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_5_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_5_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_5_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_5_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_6_clock = clock;
  assign reservation_station_6_reset = reset;
  assign reservation_station_6_io_i_allocated_idx = write_idx2 == 6'h6; // @[reservation_station.scala 246:65]
  assign reservation_station_6_io_i_issue_granted = (_issue1_func_code_T_6 | _issued_age_pack_issued_ages_1_T_6) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_6_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_6_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_6_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_6_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_6_io_i_write_slot = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_6_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_6_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_6_io_i_uop_valid = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_pc = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_inst = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_func_code = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_target = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_branch_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_select = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_taken = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_phy_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_stale_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_arch_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_inst_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_regWen = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_src1_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_phy_rs1 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_arch_rs1 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_src2_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_phy_rs2 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_arch_rs2 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_rob_idx = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_imm = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_src1_value = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_src2_value = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_op1_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_op2_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_alu_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_branch_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_uop_mem_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_6_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_6_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_6_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_6_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_6_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_6_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_6_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_6_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_6_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_6_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_7_clock = clock;
  assign reservation_station_7_reset = reset;
  assign reservation_station_7_io_i_allocated_idx = write_idx2 == 6'h7; // @[reservation_station.scala 246:65]
  assign reservation_station_7_io_i_issue_granted = (_issue1_func_code_T_7 | _issued_age_pack_issued_ages_1_T_7) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_7_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_7_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_7_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_7_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_7_io_i_write_slot = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_7_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_7_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_7_io_i_uop_valid = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_pc = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_inst = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_func_code = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_target = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_branch_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_select = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_taken = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_phy_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_stale_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_arch_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_inst_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_regWen = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_src1_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_phy_rs1 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_arch_rs1 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_src2_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_phy_rs2 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_arch_rs2 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_rob_idx = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_imm = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_src1_value = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_src2_value = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_op1_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_op2_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_alu_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_branch_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_uop_mem_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_7_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_7_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_7_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_7_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_7_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_7_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_7_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_7_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_7_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_7_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_8_clock = clock;
  assign reservation_station_8_reset = reset;
  assign reservation_station_8_io_i_allocated_idx = write_idx2 == 6'h8; // @[reservation_station.scala 246:65]
  assign reservation_station_8_io_i_issue_granted = (_issue1_func_code_T_8 | _issued_age_pack_issued_ages_1_T_8) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_8_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_8_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_8_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_8_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_8_io_i_write_slot = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_8_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_8_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_8_io_i_uop_valid = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_pc = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_inst = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_func_code = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_target = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_branch_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_select = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_taken = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_phy_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_stale_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_arch_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_inst_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_regWen = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_src1_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_phy_rs1 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_arch_rs1 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_src2_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_phy_rs2 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_arch_rs2 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_rob_idx = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_imm = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_src1_value = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_src2_value = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_op1_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_op2_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_alu_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_branch_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_uop_mem_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_8_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_8_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_8_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_8_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_8_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_8_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_8_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_8_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_8_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_8_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_9_clock = clock;
  assign reservation_station_9_reset = reset;
  assign reservation_station_9_io_i_allocated_idx = write_idx2 == 6'h9; // @[reservation_station.scala 246:65]
  assign reservation_station_9_io_i_issue_granted = (_issue1_func_code_T_9 | _issued_age_pack_issued_ages_1_T_9) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_9_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_9_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_9_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_9_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_9_io_i_write_slot = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : _reservation_station_9_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_9_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_9_io_i_uop_valid = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_pc = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_inst = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_func_code = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_target = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_branch_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_select = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_taken = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_phy_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_stale_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_arch_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_inst_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_regWen = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_src1_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_phy_rs1 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_arch_rs1 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_src2_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_phy_rs2 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_arch_rs2 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_rob_idx = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_imm = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_src1_value = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_src2_value = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_op1_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_op2_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_alu_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_branch_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_uop_mem_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_9_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_9_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_9_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_9_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_9_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_9_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_9_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_9_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_9_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_9_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_10_clock = clock;
  assign reservation_station_10_reset = reset;
  assign reservation_station_10_io_i_allocated_idx = write_idx2 == 6'ha; // @[reservation_station.scala 246:65]
  assign reservation_station_10_io_i_issue_granted = (_issue1_func_code_T_10 | _issued_age_pack_issued_ages_1_T_10) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_10_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_10_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_10_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_10_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_10_io_i_write_slot = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_10_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_10_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_10_io_i_uop_valid = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_pc = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_inst = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_func_code = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_target = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_branch_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_select = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_taken = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_phy_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_stale_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_arch_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_inst_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_regWen = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_src1_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_phy_rs1 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_arch_rs1 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_src2_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_phy_rs2 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_arch_rs2 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_rob_idx = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_imm = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_src1_value = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_src2_value = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_op1_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_op2_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_alu_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_branch_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_uop_mem_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_10_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_10_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_10_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_10_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_10_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_10_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_10_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_10_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_10_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_10_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_11_clock = clock;
  assign reservation_station_11_reset = reset;
  assign reservation_station_11_io_i_allocated_idx = write_idx2 == 6'hb; // @[reservation_station.scala 246:65]
  assign reservation_station_11_io_i_issue_granted = (_issue1_func_code_T_11 | _issued_age_pack_issued_ages_1_T_11) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_11_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_11_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_11_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_11_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_11_io_i_write_slot = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_11_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_11_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_11_io_i_uop_valid = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_pc = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_inst = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_func_code = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_target = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_branch_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_select = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_taken = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_phy_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_stale_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_arch_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_inst_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_regWen = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_src1_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_phy_rs1 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_arch_rs1 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_src2_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_phy_rs2 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_arch_rs2 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_rob_idx = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_imm = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_src1_value = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_src2_value = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_op1_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_op2_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_alu_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_branch_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_uop_mem_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_11_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_11_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_11_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_11_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_11_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_11_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_11_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_11_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_11_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_11_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_12_clock = clock;
  assign reservation_station_12_reset = reset;
  assign reservation_station_12_io_i_allocated_idx = write_idx2 == 6'hc; // @[reservation_station.scala 246:65]
  assign reservation_station_12_io_i_issue_granted = (_issue1_func_code_T_12 | _issued_age_pack_issued_ages_1_T_12) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_12_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_12_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_12_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_12_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_12_io_i_write_slot = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_12_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_12_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_12_io_i_uop_valid = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_pc = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_inst = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_func_code = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_target = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_branch_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_select = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_taken = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_phy_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_stale_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_arch_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_inst_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_regWen = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_src1_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_phy_rs1 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_arch_rs1 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_src2_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_phy_rs2 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_arch_rs2 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_rob_idx = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_imm = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_src1_value = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_src2_value = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_op1_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_op2_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_alu_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_branch_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_uop_mem_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_12_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_12_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_12_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_12_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_12_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_12_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_12_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_12_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_12_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_12_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_13_clock = clock;
  assign reservation_station_13_reset = reset;
  assign reservation_station_13_io_i_allocated_idx = write_idx2 == 6'hd; // @[reservation_station.scala 246:65]
  assign reservation_station_13_io_i_issue_granted = (_issue1_func_code_T_13 | _issued_age_pack_issued_ages_1_T_13) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_13_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_13_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_13_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_13_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_13_io_i_write_slot = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_13_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_13_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_13_io_i_uop_valid = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_pc = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_inst = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_func_code = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_target = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_branch_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_select = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_taken = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_phy_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_stale_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_arch_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_inst_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_regWen = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_src1_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_phy_rs1 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_arch_rs1 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_src2_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_phy_rs2 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_arch_rs2 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_rob_idx = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_imm = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_src1_value = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_src2_value = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_op1_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_op2_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_alu_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_branch_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_uop_mem_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_13_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_13_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_13_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_13_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_13_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_13_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_13_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_13_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_13_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_13_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_14_clock = clock;
  assign reservation_station_14_reset = reset;
  assign reservation_station_14_io_i_allocated_idx = write_idx2 == 6'he; // @[reservation_station.scala 246:65]
  assign reservation_station_14_io_i_issue_granted = (_issue1_func_code_T_14 | _issued_age_pack_issued_ages_1_T_14) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_14_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_14_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_14_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_14_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_14_io_i_write_slot = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_14_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_14_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_14_io_i_uop_valid = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_pc = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_inst = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_func_code = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_target = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_branch_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_select = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_taken = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_phy_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_stale_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_arch_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_inst_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_regWen = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_src1_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_phy_rs1 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_arch_rs1 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_src2_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_phy_rs2 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_arch_rs2 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_rob_idx = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_imm = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_src1_value = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_src2_value = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_op1_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_op2_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_alu_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_branch_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_uop_mem_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_14_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_14_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_14_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_14_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_14_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_14_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_14_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_14_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_14_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_14_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_15_clock = clock;
  assign reservation_station_15_reset = reset;
  assign reservation_station_15_io_i_allocated_idx = write_idx2 == 6'hf; // @[reservation_station.scala 246:65]
  assign reservation_station_15_io_i_issue_granted = (_issue1_func_code_T_15 | _issued_age_pack_issued_ages_1_T_15) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_15_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_15_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_15_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_15_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_15_io_i_write_slot = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_15_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_15_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_15_io_i_uop_valid = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_pc = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_inst = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_func_code = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_target = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_branch_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_select = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_taken = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_phy_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_stale_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_arch_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_inst_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_regWen = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_src1_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_phy_rs1 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_arch_rs1 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_src2_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_phy_rs2 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_arch_rs2 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_rob_idx = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_imm = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_src1_value = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_src2_value = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_op1_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_op2_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_alu_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_branch_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_uop_mem_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_15_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_15_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_15_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_15_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_15_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_15_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_15_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_15_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_15_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_15_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_16_clock = clock;
  assign reservation_station_16_reset = reset;
  assign reservation_station_16_io_i_allocated_idx = write_idx2 == 6'h10; // @[reservation_station.scala 246:65]
  assign reservation_station_16_io_i_issue_granted = (_issue1_func_code_T_16 | _issued_age_pack_issued_ages_1_T_16) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_16_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_16_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_16_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_16_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_16_io_i_write_slot = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_16_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_16_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_16_io_i_uop_valid = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_pc = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_inst = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_func_code = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_target = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_branch_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_select = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_taken = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_phy_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_stale_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_arch_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_inst_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_regWen = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_src1_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_phy_rs1 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_arch_rs1 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_src2_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_phy_rs2 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_arch_rs2 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_rob_idx = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_imm = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_src1_value = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_src2_value = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_op1_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_op2_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_alu_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_branch_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_uop_mem_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_16_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_16_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_16_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_16_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_16_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_16_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_16_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_16_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_16_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_16_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_17_clock = clock;
  assign reservation_station_17_reset = reset;
  assign reservation_station_17_io_i_allocated_idx = write_idx2 == 6'h11; // @[reservation_station.scala 246:65]
  assign reservation_station_17_io_i_issue_granted = (_issue1_func_code_T_17 | _issued_age_pack_issued_ages_1_T_17) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_17_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_17_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_17_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_17_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_17_io_i_write_slot = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_17_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_17_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_17_io_i_uop_valid = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_pc = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_inst = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_func_code = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_target = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_branch_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_select = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_taken = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_phy_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_stale_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_arch_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_inst_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_regWen = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_src1_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_phy_rs1 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_arch_rs1 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_src2_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_phy_rs2 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_arch_rs2 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_rob_idx = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_imm = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_src1_value = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_src2_value = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_op1_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_op2_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_alu_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_branch_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_uop_mem_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_17_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_17_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_17_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_17_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_17_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_17_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_17_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_17_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_17_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_17_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_18_clock = clock;
  assign reservation_station_18_reset = reset;
  assign reservation_station_18_io_i_allocated_idx = write_idx2 == 6'h12; // @[reservation_station.scala 246:65]
  assign reservation_station_18_io_i_issue_granted = (_issue1_func_code_T_18 | _issued_age_pack_issued_ages_1_T_18) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_18_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_18_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_18_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_18_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_18_io_i_write_slot = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_18_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_18_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_18_io_i_uop_valid = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_pc = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_inst = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_func_code = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_target = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_branch_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_select = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_taken = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_phy_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_stale_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_arch_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_inst_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_regWen = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_src1_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_phy_rs1 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_arch_rs1 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_src2_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_phy_rs2 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_arch_rs2 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_rob_idx = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_imm = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_src1_value = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_src2_value = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_op1_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_op2_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_alu_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_branch_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_uop_mem_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_18_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_18_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_18_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_18_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_18_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_18_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_18_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_18_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_18_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_18_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_19_clock = clock;
  assign reservation_station_19_reset = reset;
  assign reservation_station_19_io_i_allocated_idx = write_idx2 == 6'h13; // @[reservation_station.scala 246:65]
  assign reservation_station_19_io_i_issue_granted = (_issue1_func_code_T_19 | _issued_age_pack_issued_ages_1_T_19) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_19_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_19_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_19_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_19_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_19_io_i_write_slot = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_19_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_19_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_19_io_i_uop_valid = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_pc = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_inst = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_func_code = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_target = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_branch_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_select = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_taken = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_phy_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_stale_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_arch_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_inst_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_regWen = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_src1_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_phy_rs1 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_arch_rs1 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_src2_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_phy_rs2 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_arch_rs2 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_rob_idx = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_imm = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_src1_value = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_src2_value = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_op1_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_op2_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_alu_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_branch_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_uop_mem_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_19_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_19_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_19_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_19_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_19_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_19_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_19_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_19_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_19_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_19_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_20_clock = clock;
  assign reservation_station_20_reset = reset;
  assign reservation_station_20_io_i_allocated_idx = write_idx2 == 6'h14; // @[reservation_station.scala 246:65]
  assign reservation_station_20_io_i_issue_granted = (_issue1_func_code_T_20 | _issued_age_pack_issued_ages_1_T_20) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_20_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_20_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_20_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_20_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_20_io_i_write_slot = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_20_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_20_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_20_io_i_uop_valid = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_pc = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_inst = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_func_code = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_target = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_branch_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_select = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_taken = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_phy_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_stale_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_arch_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_inst_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_regWen = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_src1_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_phy_rs1 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_arch_rs1 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_src2_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_phy_rs2 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_arch_rs2 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_rob_idx = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_imm = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_src1_value = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_src2_value = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_op1_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_op2_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_alu_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_branch_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_uop_mem_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_20_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_20_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_20_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_20_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_20_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_20_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_20_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_20_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_20_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_20_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_21_clock = clock;
  assign reservation_station_21_reset = reset;
  assign reservation_station_21_io_i_allocated_idx = write_idx2 == 6'h15; // @[reservation_station.scala 246:65]
  assign reservation_station_21_io_i_issue_granted = (_issue1_func_code_T_21 | _issued_age_pack_issued_ages_1_T_21) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_21_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_21_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_21_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_21_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_21_io_i_write_slot = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_21_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_21_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_21_io_i_uop_valid = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_pc = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_inst = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_func_code = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_target = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_branch_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_select = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_taken = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_phy_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_stale_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_arch_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_inst_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_regWen = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_src1_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_phy_rs1 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_arch_rs1 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_src2_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_phy_rs2 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_arch_rs2 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_rob_idx = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_imm = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_src1_value = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_src2_value = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_op1_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_op2_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_alu_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_branch_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_uop_mem_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_21_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_21_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_21_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_21_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_21_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_21_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_21_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_21_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_21_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_21_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_22_clock = clock;
  assign reservation_station_22_reset = reset;
  assign reservation_station_22_io_i_allocated_idx = write_idx2 == 6'h16; // @[reservation_station.scala 246:65]
  assign reservation_station_22_io_i_issue_granted = (_issue1_func_code_T_22 | _issued_age_pack_issued_ages_1_T_22) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_22_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_22_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_22_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_22_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_22_io_i_write_slot = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_22_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_22_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_22_io_i_uop_valid = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_pc = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_inst = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_func_code = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_target = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_branch_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_select = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_taken = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_phy_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_stale_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_arch_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_inst_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_regWen = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_src1_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_phy_rs1 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_arch_rs1 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_src2_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_phy_rs2 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_arch_rs2 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_rob_idx = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_imm = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_src1_value = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_src2_value = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_op1_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_op2_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_alu_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_branch_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_uop_mem_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_22_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_22_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_22_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_22_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_22_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_22_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_22_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_22_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_22_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_22_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_23_clock = clock;
  assign reservation_station_23_reset = reset;
  assign reservation_station_23_io_i_allocated_idx = write_idx2 == 6'h17; // @[reservation_station.scala 246:65]
  assign reservation_station_23_io_i_issue_granted = (_issue1_func_code_T_23 | _issued_age_pack_issued_ages_1_T_23) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_23_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_23_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_23_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_23_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_23_io_i_write_slot = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_23_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_23_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_23_io_i_uop_valid = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_pc = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_inst = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_func_code = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_target = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_branch_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_select = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_taken = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_phy_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_stale_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_arch_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_inst_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_regWen = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_src1_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_phy_rs1 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_arch_rs1 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_src2_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_phy_rs2 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_arch_rs2 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_rob_idx = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_imm = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_src1_value = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_src2_value = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_op1_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_op2_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_alu_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_branch_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_uop_mem_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_23_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_23_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_23_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_23_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_23_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_23_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_23_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_23_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_23_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_23_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_24_clock = clock;
  assign reservation_station_24_reset = reset;
  assign reservation_station_24_io_i_allocated_idx = write_idx2 == 6'h18; // @[reservation_station.scala 246:65]
  assign reservation_station_24_io_i_issue_granted = (_issue1_func_code_T_24 | _issued_age_pack_issued_ages_1_T_24) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_24_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_24_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_24_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_24_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_24_io_i_write_slot = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_24_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_24_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_24_io_i_uop_valid = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_pc = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_inst = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_func_code = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_target = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_branch_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_select = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_taken = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_phy_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_stale_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_arch_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_inst_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_regWen = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_src1_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_phy_rs1 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_arch_rs1 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_src2_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_phy_rs2 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_arch_rs2 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_rob_idx = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_imm = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_src1_value = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_src2_value = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_op1_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_op2_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_alu_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_branch_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_uop_mem_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_24_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_24_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_24_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_24_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_24_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_24_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_24_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_24_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_24_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_24_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_25_clock = clock;
  assign reservation_station_25_reset = reset;
  assign reservation_station_25_io_i_allocated_idx = write_idx2 == 6'h19; // @[reservation_station.scala 246:65]
  assign reservation_station_25_io_i_issue_granted = (_issue1_func_code_T_25 | _issued_age_pack_issued_ages_1_T_25) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_25_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_25_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_25_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_25_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_25_io_i_write_slot = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_25_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_25_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_25_io_i_uop_valid = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_pc = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_inst = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_func_code = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_target = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_branch_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_select = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_taken = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_phy_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_stale_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_arch_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_inst_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_regWen = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_src1_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_phy_rs1 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_arch_rs1 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_src2_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_phy_rs2 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_arch_rs2 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_rob_idx = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_imm = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_src1_value = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_src2_value = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_op1_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_op2_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_alu_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_branch_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_uop_mem_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_25_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_25_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_25_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_25_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_25_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_25_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_25_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_25_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_25_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_25_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_26_clock = clock;
  assign reservation_station_26_reset = reset;
  assign reservation_station_26_io_i_allocated_idx = write_idx2 == 6'h1a; // @[reservation_station.scala 246:65]
  assign reservation_station_26_io_i_issue_granted = (_issue1_func_code_T_26 | _issued_age_pack_issued_ages_1_T_26) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_26_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_26_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_26_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_26_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_26_io_i_write_slot = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_26_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_26_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_26_io_i_uop_valid = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_pc = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_inst = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_func_code = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_target = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_branch_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_select = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_taken = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_phy_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_stale_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_arch_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_inst_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_regWen = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_src1_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_phy_rs1 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_arch_rs1 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_src2_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_phy_rs2 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_arch_rs2 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_rob_idx = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_imm = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_src1_value = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_src2_value = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_op1_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_op2_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_alu_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_branch_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_uop_mem_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_26_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_26_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_26_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_26_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_26_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_26_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_26_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_26_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_26_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_26_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_27_clock = clock;
  assign reservation_station_27_reset = reset;
  assign reservation_station_27_io_i_allocated_idx = write_idx2 == 6'h1b; // @[reservation_station.scala 246:65]
  assign reservation_station_27_io_i_issue_granted = (_issue1_func_code_T_27 | _issued_age_pack_issued_ages_1_T_27) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_27_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_27_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_27_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_27_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_27_io_i_write_slot = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_27_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_27_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_27_io_i_uop_valid = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_pc = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_inst = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_func_code = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_target = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_branch_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_select = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_taken = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_phy_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_stale_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_arch_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_inst_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_regWen = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_src1_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_phy_rs1 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_arch_rs1 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_src2_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_phy_rs2 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_arch_rs2 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_rob_idx = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_imm = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_src1_value = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_src2_value = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_op1_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_op2_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_alu_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_branch_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_uop_mem_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_27_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_27_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_27_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_27_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_27_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_27_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_27_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_27_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_27_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_27_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_28_clock = clock;
  assign reservation_station_28_reset = reset;
  assign reservation_station_28_io_i_allocated_idx = write_idx2 == 6'h1c; // @[reservation_station.scala 246:65]
  assign reservation_station_28_io_i_issue_granted = (_issue1_func_code_T_28 | _issued_age_pack_issued_ages_1_T_28) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_28_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_28_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_28_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_28_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_28_io_i_write_slot = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_28_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_28_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_28_io_i_uop_valid = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_pc = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_inst = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_func_code = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_target = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_branch_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_select = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_taken = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_phy_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_stale_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_arch_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_inst_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_regWen = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_src1_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_phy_rs1 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_arch_rs1 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_src2_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_phy_rs2 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_arch_rs2 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_rob_idx = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_imm = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_src1_value = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_src2_value = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_op1_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_op2_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_alu_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_branch_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_uop_mem_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_28_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_28_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_28_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_28_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_28_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_28_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_28_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_28_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_28_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_28_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_29_clock = clock;
  assign reservation_station_29_reset = reset;
  assign reservation_station_29_io_i_allocated_idx = write_idx2 == 6'h1d; // @[reservation_station.scala 246:65]
  assign reservation_station_29_io_i_issue_granted = (_issue1_func_code_T_29 | _issued_age_pack_issued_ages_1_T_29) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_29_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_29_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_29_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_29_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_29_io_i_write_slot = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_29_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_29_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_29_io_i_uop_valid = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_pc = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_inst = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_func_code = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_target = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_branch_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_select = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_taken = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_phy_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_stale_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_arch_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_inst_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_regWen = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_src1_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_phy_rs1 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_arch_rs1 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_src2_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_phy_rs2 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_arch_rs2 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_rob_idx = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_imm = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_src1_value = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_src2_value = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_op1_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_op2_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_alu_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_branch_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_uop_mem_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_29_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_29_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_29_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_29_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_29_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_29_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_29_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_29_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_29_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_29_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_30_clock = clock;
  assign reservation_station_30_reset = reset;
  assign reservation_station_30_io_i_allocated_idx = write_idx2 == 6'h1e; // @[reservation_station.scala 246:65]
  assign reservation_station_30_io_i_issue_granted = (_issue1_func_code_T_30 | _issued_age_pack_issued_ages_1_T_30) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_30_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_30_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_30_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_30_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_30_io_i_write_slot = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_30_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_30_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_30_io_i_uop_valid = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_pc = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_inst = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_func_code = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_target = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_branch_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_select = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_taken = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_phy_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_stale_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_arch_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_inst_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_regWen = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_src1_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_phy_rs1 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_arch_rs1 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_src2_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_phy_rs2 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_arch_rs2 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_rob_idx = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_imm = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_src1_value = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_src2_value = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_op1_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_op2_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_alu_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_branch_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_uop_mem_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_30_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_30_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_30_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_30_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_30_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_30_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_30_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_30_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_30_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_30_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_31_clock = clock;
  assign reservation_station_31_reset = reset;
  assign reservation_station_31_io_i_allocated_idx = write_idx2 == 6'h1f; // @[reservation_station.scala 246:65]
  assign reservation_station_31_io_i_issue_granted = (_issue1_func_code_T_31 | _issued_age_pack_issued_ages_1_T_31) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_31_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_31_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_31_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_31_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_31_io_i_write_slot = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_31_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_31_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_31_io_i_uop_valid = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_pc = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_inst = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_func_code = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_target = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_branch_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_select = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_taken = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_phy_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_stale_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_arch_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_inst_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_regWen = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_src1_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_phy_rs1 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_arch_rs1 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_src2_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_phy_rs2 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_arch_rs2 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_rob_idx = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_imm = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_src1_value = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_src2_value = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_op1_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_op2_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_alu_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_branch_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_uop_mem_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_31_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_31_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_31_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_31_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_31_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_31_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_31_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_31_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_31_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_31_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_32_clock = clock;
  assign reservation_station_32_reset = reset;
  assign reservation_station_32_io_i_allocated_idx = write_idx2 == 6'h20; // @[reservation_station.scala 246:65]
  assign reservation_station_32_io_i_issue_granted = (_issue1_func_code_T_32 | _issued_age_pack_issued_ages_1_T_32) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_32_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_32_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_32_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_32_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_32_io_i_write_slot = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_32_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_32_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_32_io_i_uop_valid = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_pc = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_inst = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_func_code = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_valid = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_target = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_branch_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_select = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_taken = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_phy_dst = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_stale_dst = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_arch_dst = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_inst_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_regWen = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_src1_valid = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_phy_rs1 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_arch_rs1 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_src2_valid = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_phy_rs2 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_arch_rs2 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_rob_idx = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_imm = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_src1_value = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_src2_value = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_op1_sel = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_op2_sel = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_alu_sel = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_branch_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_uop_mem_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_32_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_32_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_32_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_32_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_32_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_32_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_32_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_32_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_32_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_32_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_33_clock = clock;
  assign reservation_station_33_reset = reset;
  assign reservation_station_33_io_i_allocated_idx = write_idx2 == 6'h21; // @[reservation_station.scala 246:65]
  assign reservation_station_33_io_i_issue_granted = (_issue1_func_code_T_33 | _issued_age_pack_issued_ages_1_T_33) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_33_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_33_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_33_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_33_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_33_io_i_write_slot = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_33_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_33_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_33_io_i_uop_valid = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_pc = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_inst = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_func_code = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_valid = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_target = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_branch_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_select = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_taken = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_phy_dst = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_stale_dst = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_arch_dst = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_inst_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_regWen = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_src1_valid = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_phy_rs1 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_arch_rs1 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_src2_valid = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_phy_rs2 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_arch_rs2 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_rob_idx = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_imm = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_src1_value = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_src2_value = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_op1_sel = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_op2_sel = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_alu_sel = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_branch_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_uop_mem_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_33_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_33_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_33_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_33_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_33_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_33_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_33_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_33_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_33_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_33_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_34_clock = clock;
  assign reservation_station_34_reset = reset;
  assign reservation_station_34_io_i_allocated_idx = write_idx2 == 6'h22; // @[reservation_station.scala 246:65]
  assign reservation_station_34_io_i_issue_granted = (_issue1_func_code_T_34 | _issued_age_pack_issued_ages_1_T_34) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_34_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_34_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_34_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_34_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_34_io_i_write_slot = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_34_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_34_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_34_io_i_uop_valid = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_pc = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_inst = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_func_code = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_valid = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_target = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_branch_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_select = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_taken = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_phy_dst = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_stale_dst = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_arch_dst = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_inst_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_regWen = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_src1_valid = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_phy_rs1 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_arch_rs1 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_src2_valid = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_phy_rs2 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_arch_rs2 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_rob_idx = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_imm = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_src1_value = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_src2_value = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_op1_sel = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_op2_sel = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_alu_sel = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_branch_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_uop_mem_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_34_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_34_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_34_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_34_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_34_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_34_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_34_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_34_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_34_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_34_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_35_clock = clock;
  assign reservation_station_35_reset = reset;
  assign reservation_station_35_io_i_allocated_idx = write_idx2 == 6'h23; // @[reservation_station.scala 246:65]
  assign reservation_station_35_io_i_issue_granted = (_issue1_func_code_T_35 | _issued_age_pack_issued_ages_1_T_35) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_35_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_35_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_35_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_35_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_35_io_i_write_slot = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_35_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_35_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_35_io_i_uop_valid = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_pc = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_inst = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_func_code = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_valid = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_target = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_branch_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_select = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_taken = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_phy_dst = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_stale_dst = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_arch_dst = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_inst_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_regWen = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_src1_valid = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_phy_rs1 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_arch_rs1 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_src2_valid = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_phy_rs2 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_arch_rs2 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_rob_idx = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_imm = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_src1_value = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_src2_value = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_op1_sel = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_op2_sel = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_alu_sel = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_branch_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_uop_mem_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_35_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_35_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_35_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_35_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_35_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_35_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_35_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_35_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_35_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_35_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_36_clock = clock;
  assign reservation_station_36_reset = reset;
  assign reservation_station_36_io_i_allocated_idx = write_idx2 == 6'h24; // @[reservation_station.scala 246:65]
  assign reservation_station_36_io_i_issue_granted = (_issue1_func_code_T_36 | _issued_age_pack_issued_ages_1_T_36) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_36_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_36_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_36_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_36_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_36_io_i_write_slot = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_36_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_36_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_36_io_i_uop_valid = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_pc = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_inst = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_func_code = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_valid = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_target = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_branch_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_select = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_taken = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_phy_dst = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_stale_dst = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_arch_dst = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_inst_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_regWen = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_src1_valid = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_phy_rs1 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_arch_rs1 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_src2_valid = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_phy_rs2 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_arch_rs2 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_rob_idx = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_imm = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_src1_value = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_src2_value = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_op1_sel = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_op2_sel = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_alu_sel = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_branch_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_uop_mem_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_36_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_36_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_36_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_36_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_36_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_36_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_36_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_36_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_36_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_36_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_37_clock = clock;
  assign reservation_station_37_reset = reset;
  assign reservation_station_37_io_i_allocated_idx = write_idx2 == 6'h25; // @[reservation_station.scala 246:65]
  assign reservation_station_37_io_i_issue_granted = (_issue1_func_code_T_37 | _issued_age_pack_issued_ages_1_T_37) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_37_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_37_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_37_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_37_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_37_io_i_write_slot = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_37_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_37_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_37_io_i_uop_valid = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_pc = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_inst = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_func_code = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_valid = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_target = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_branch_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_select = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_taken = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_phy_dst = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_stale_dst = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_arch_dst = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_inst_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_regWen = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_src1_valid = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_phy_rs1 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_arch_rs1 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_src2_valid = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_phy_rs2 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_arch_rs2 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_rob_idx = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_imm = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_src1_value = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_src2_value = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_op1_sel = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_op2_sel = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_alu_sel = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_branch_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_uop_mem_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_37_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_37_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_37_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_37_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_37_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_37_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_37_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_37_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_37_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_37_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_38_clock = clock;
  assign reservation_station_38_reset = reset;
  assign reservation_station_38_io_i_allocated_idx = write_idx2 == 6'h26; // @[reservation_station.scala 246:65]
  assign reservation_station_38_io_i_issue_granted = (_issue1_func_code_T_38 | _issued_age_pack_issued_ages_1_T_38) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_38_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_38_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_38_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_38_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_38_io_i_write_slot = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_38_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_38_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_38_io_i_uop_valid = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_pc = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_inst = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_func_code = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_valid = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_target = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_branch_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_select = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_taken = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_phy_dst = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_stale_dst = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_arch_dst = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_inst_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_regWen = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_src1_valid = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_phy_rs1 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_arch_rs1 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_src2_valid = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_phy_rs2 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_arch_rs2 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_rob_idx = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_imm = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_src1_value = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_src2_value = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_op1_sel = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_op2_sel = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_alu_sel = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_branch_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_uop_mem_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_38_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_38_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_38_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_38_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_38_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_38_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_38_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_38_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_38_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_38_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_39_clock = clock;
  assign reservation_station_39_reset = reset;
  assign reservation_station_39_io_i_allocated_idx = write_idx2 == 6'h27; // @[reservation_station.scala 246:65]
  assign reservation_station_39_io_i_issue_granted = (_issue1_func_code_T_39 | _issued_age_pack_issued_ages_1_T_39) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_39_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_39_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_39_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_39_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_39_io_i_write_slot = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_39_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_39_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_39_io_i_uop_valid = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_pc = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_inst = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_func_code = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_valid = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_target = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_branch_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_select = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_taken = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_phy_dst = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_stale_dst = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_arch_dst = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_inst_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_regWen = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_src1_valid = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_phy_rs1 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_arch_rs1 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_src2_valid = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_phy_rs2 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_arch_rs2 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_rob_idx = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_imm = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_src1_value = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_src2_value = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_op1_sel = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_op2_sel = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_alu_sel = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_branch_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_uop_mem_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_39_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_39_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_39_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_39_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_39_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_39_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_39_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_39_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_39_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_39_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_40_clock = clock;
  assign reservation_station_40_reset = reset;
  assign reservation_station_40_io_i_allocated_idx = write_idx2 == 6'h28; // @[reservation_station.scala 246:65]
  assign reservation_station_40_io_i_issue_granted = (_issue1_func_code_T_40 | _issued_age_pack_issued_ages_1_T_40) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_40_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_40_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_40_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_40_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_40_io_i_write_slot = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_40_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_40_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_40_io_i_uop_valid = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_pc = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_inst = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_func_code = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_valid = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_target = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_branch_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_select = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_taken = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_phy_dst = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_stale_dst = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_arch_dst = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_inst_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_regWen = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_src1_valid = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_phy_rs1 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_arch_rs1 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_src2_valid = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_phy_rs2 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_arch_rs2 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_rob_idx = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_imm = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_src1_value = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_src2_value = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_op1_sel = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_op2_sel = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_alu_sel = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_branch_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_uop_mem_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_40_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_40_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_40_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_40_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_40_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_40_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_40_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_40_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_40_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_40_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_41_clock = clock;
  assign reservation_station_41_reset = reset;
  assign reservation_station_41_io_i_allocated_idx = write_idx2 == 6'h29; // @[reservation_station.scala 246:65]
  assign reservation_station_41_io_i_issue_granted = (_issue1_func_code_T_41 | _issued_age_pack_issued_ages_1_T_41) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_41_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_41_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_41_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_41_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_41_io_i_write_slot = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_41_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_41_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_41_io_i_uop_valid = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_pc = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_inst = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_func_code = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_valid = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_target = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_branch_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_select = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_taken = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_phy_dst = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_stale_dst = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_arch_dst = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_inst_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_regWen = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_src1_valid = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_phy_rs1 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_arch_rs1 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_src2_valid = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_phy_rs2 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_arch_rs2 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_rob_idx = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_imm = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_src1_value = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_src2_value = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_op1_sel = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_op2_sel = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_alu_sel = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_branch_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_uop_mem_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_41_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_41_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_41_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_41_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_41_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_41_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_41_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_41_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_41_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_41_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_42_clock = clock;
  assign reservation_station_42_reset = reset;
  assign reservation_station_42_io_i_allocated_idx = write_idx2 == 6'h2a; // @[reservation_station.scala 246:65]
  assign reservation_station_42_io_i_issue_granted = (_issue1_func_code_T_42 | _issued_age_pack_issued_ages_1_T_42) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_42_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_42_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_42_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_42_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_42_io_i_write_slot = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_42_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_42_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_42_io_i_uop_valid = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_pc = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_inst = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_func_code = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_valid = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_target = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_branch_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_select = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_taken = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_phy_dst = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_stale_dst = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_arch_dst = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_inst_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_regWen = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_src1_valid = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_phy_rs1 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_arch_rs1 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_src2_valid = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_phy_rs2 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_arch_rs2 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_rob_idx = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_imm = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_src1_value = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_src2_value = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_op1_sel = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_op2_sel = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_alu_sel = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_branch_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_uop_mem_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_42_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_42_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_42_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_42_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_42_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_42_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_42_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_42_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_42_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_42_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_43_clock = clock;
  assign reservation_station_43_reset = reset;
  assign reservation_station_43_io_i_allocated_idx = write_idx2 == 6'h2b; // @[reservation_station.scala 246:65]
  assign reservation_station_43_io_i_issue_granted = (_issue1_func_code_T_43 | _issued_age_pack_issued_ages_1_T_43) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_43_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_43_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_43_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_43_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_43_io_i_write_slot = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_43_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_43_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_43_io_i_uop_valid = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_pc = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_inst = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_func_code = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_valid = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_target = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_branch_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_select = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_taken = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_phy_dst = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_stale_dst = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_arch_dst = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_inst_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_regWen = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_src1_valid = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_phy_rs1 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_arch_rs1 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_src2_valid = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_phy_rs2 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_arch_rs2 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_rob_idx = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_imm = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_src1_value = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_src2_value = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_op1_sel = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_op2_sel = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_alu_sel = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_branch_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_uop_mem_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_43_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_43_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_43_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_43_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_43_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_43_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_43_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_43_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_43_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_43_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_44_clock = clock;
  assign reservation_station_44_reset = reset;
  assign reservation_station_44_io_i_allocated_idx = write_idx2 == 6'h2c; // @[reservation_station.scala 246:65]
  assign reservation_station_44_io_i_issue_granted = (_issue1_func_code_T_44 | _issued_age_pack_issued_ages_1_T_44) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_44_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_44_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_44_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_44_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_44_io_i_write_slot = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_44_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_44_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_44_io_i_uop_valid = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_pc = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_inst = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_func_code = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_valid = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_target = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_branch_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_select = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_taken = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_phy_dst = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_stale_dst = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_arch_dst = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_inst_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_regWen = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_src1_valid = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_phy_rs1 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_arch_rs1 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_src2_valid = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_phy_rs2 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_arch_rs2 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_rob_idx = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_imm = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_src1_value = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_src2_value = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_op1_sel = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_op2_sel = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_alu_sel = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_branch_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_uop_mem_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_44_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_44_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_44_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_44_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_44_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_44_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_44_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_44_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_44_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_44_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_45_clock = clock;
  assign reservation_station_45_reset = reset;
  assign reservation_station_45_io_i_allocated_idx = write_idx2 == 6'h2d; // @[reservation_station.scala 246:65]
  assign reservation_station_45_io_i_issue_granted = (_issue1_func_code_T_45 | _issued_age_pack_issued_ages_1_T_45) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_45_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_45_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_45_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_45_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_45_io_i_write_slot = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_45_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_45_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_45_io_i_uop_valid = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_pc = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_inst = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_func_code = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_valid = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_target = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_branch_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_select = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_taken = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_phy_dst = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_stale_dst = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_arch_dst = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_inst_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_regWen = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_src1_valid = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_phy_rs1 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_arch_rs1 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_src2_valid = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_phy_rs2 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_arch_rs2 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_rob_idx = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_imm = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_src1_value = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_src2_value = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_op1_sel = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_op2_sel = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_alu_sel = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_branch_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_uop_mem_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_45_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_45_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_45_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_45_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_45_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_45_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_45_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_45_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_45_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_45_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_46_clock = clock;
  assign reservation_station_46_reset = reset;
  assign reservation_station_46_io_i_allocated_idx = write_idx2 == 6'h2e; // @[reservation_station.scala 246:65]
  assign reservation_station_46_io_i_issue_granted = (_issue1_func_code_T_46 | _issued_age_pack_issued_ages_1_T_46) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_46_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_46_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_46_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_46_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_46_io_i_write_slot = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_46_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_46_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_46_io_i_uop_valid = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_pc = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_inst = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_func_code = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_valid = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_target = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_branch_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_select = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_taken = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_phy_dst = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_stale_dst = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_arch_dst = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_inst_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_regWen = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_src1_valid = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_phy_rs1 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_arch_rs1 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_src2_valid = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_phy_rs2 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_arch_rs2 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_rob_idx = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_imm = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_src1_value = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_src2_value = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_op1_sel = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_op2_sel = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_alu_sel = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_branch_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_uop_mem_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_46_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_46_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_46_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_46_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_46_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_46_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_46_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_46_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_46_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_46_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_47_clock = clock;
  assign reservation_station_47_reset = reset;
  assign reservation_station_47_io_i_allocated_idx = write_idx2 == 6'h2f; // @[reservation_station.scala 246:65]
  assign reservation_station_47_io_i_issue_granted = (_issue1_func_code_T_47 | _issued_age_pack_issued_ages_1_T_47) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_47_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_47_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_47_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_47_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_47_io_i_write_slot = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_47_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_47_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_47_io_i_uop_valid = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_pc = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_inst = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_func_code = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_valid = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_target = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_branch_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_select = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_taken = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_phy_dst = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_stale_dst = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_arch_dst = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_inst_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_regWen = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_src1_valid = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_phy_rs1 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_arch_rs1 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_src2_valid = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_phy_rs2 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_arch_rs2 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_rob_idx = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_imm = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_src1_value = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_src2_value = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_op1_sel = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_op2_sel = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_alu_sel = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_branch_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_uop_mem_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_47_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_47_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_47_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_47_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_47_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_47_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_47_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_47_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_47_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_47_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_48_clock = clock;
  assign reservation_station_48_reset = reset;
  assign reservation_station_48_io_i_allocated_idx = write_idx2 == 6'h30; // @[reservation_station.scala 246:65]
  assign reservation_station_48_io_i_issue_granted = (_issue1_func_code_T_48 | _issued_age_pack_issued_ages_1_T_48) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_48_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_48_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_48_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_48_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_48_io_i_write_slot = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_48_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_48_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_48_io_i_uop_valid = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_pc = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_inst = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_func_code = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_valid = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_target = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_branch_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_select = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_taken = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_phy_dst = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_stale_dst = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_arch_dst = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_inst_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_regWen = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_src1_valid = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_phy_rs1 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_arch_rs1 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_src2_valid = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_phy_rs2 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_arch_rs2 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_rob_idx = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_imm = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_src1_value = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_src2_value = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_op1_sel = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_op2_sel = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_alu_sel = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_branch_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_uop_mem_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_48_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_48_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_48_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_48_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_48_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_48_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_48_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_48_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_48_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_48_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_49_clock = clock;
  assign reservation_station_49_reset = reset;
  assign reservation_station_49_io_i_allocated_idx = write_idx2 == 6'h31; // @[reservation_station.scala 246:65]
  assign reservation_station_49_io_i_issue_granted = (_issue1_func_code_T_49 | _issued_age_pack_issued_ages_1_T_49) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_49_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_49_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_49_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_49_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_49_io_i_write_slot = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_49_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_49_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_49_io_i_uop_valid = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_pc = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_inst = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_func_code = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_valid = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_target = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_branch_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_select = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_taken = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_phy_dst = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_stale_dst = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_arch_dst = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_inst_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_regWen = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_src1_valid = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_phy_rs1 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_arch_rs1 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_src2_valid = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_phy_rs2 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_arch_rs2 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_rob_idx = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_imm = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_src1_value = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_src2_value = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_op1_sel = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_op2_sel = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_alu_sel = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_branch_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_uop_mem_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_49_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_49_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_49_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_49_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_49_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_49_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_49_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_49_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_49_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_49_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_50_clock = clock;
  assign reservation_station_50_reset = reset;
  assign reservation_station_50_io_i_allocated_idx = write_idx2 == 6'h32; // @[reservation_station.scala 246:65]
  assign reservation_station_50_io_i_issue_granted = (_issue1_func_code_T_50 | _issued_age_pack_issued_ages_1_T_50) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_50_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_50_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_50_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_50_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_50_io_i_write_slot = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_50_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_50_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_50_io_i_uop_valid = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_pc = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_inst = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_func_code = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_valid = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_target = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_branch_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_select = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_taken = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_phy_dst = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_stale_dst = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_arch_dst = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_inst_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_regWen = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_src1_valid = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_phy_rs1 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_arch_rs1 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_src2_valid = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_phy_rs2 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_arch_rs2 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_rob_idx = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_imm = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_src1_value = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_src2_value = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_op1_sel = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_op2_sel = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_alu_sel = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_branch_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_uop_mem_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_50_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_50_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_50_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_50_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_50_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_50_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_50_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_50_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_50_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_50_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_51_clock = clock;
  assign reservation_station_51_reset = reset;
  assign reservation_station_51_io_i_allocated_idx = write_idx2 == 6'h33; // @[reservation_station.scala 246:65]
  assign reservation_station_51_io_i_issue_granted = (_issue1_func_code_T_51 | _issued_age_pack_issued_ages_1_T_51) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_51_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_51_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_51_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_51_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_51_io_i_write_slot = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_51_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_51_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_51_io_i_uop_valid = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_pc = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_inst = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_func_code = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_valid = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_target = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_branch_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_select = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_taken = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_phy_dst = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_stale_dst = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_arch_dst = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_inst_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_regWen = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_src1_valid = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_phy_rs1 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_arch_rs1 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_src2_valid = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_phy_rs2 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_arch_rs2 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_rob_idx = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_imm = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_src1_value = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_src2_value = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_op1_sel = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_op2_sel = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_alu_sel = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_branch_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_uop_mem_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_51_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_51_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_51_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_51_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_51_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_51_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_51_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_51_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_51_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_51_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_52_clock = clock;
  assign reservation_station_52_reset = reset;
  assign reservation_station_52_io_i_allocated_idx = write_idx2 == 6'h34; // @[reservation_station.scala 246:65]
  assign reservation_station_52_io_i_issue_granted = (_issue1_func_code_T_52 | _issued_age_pack_issued_ages_1_T_52) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_52_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_52_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_52_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_52_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_52_io_i_write_slot = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_52_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_52_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_52_io_i_uop_valid = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_pc = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_inst = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_func_code = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_valid = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_target = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_branch_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_select = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_taken = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_phy_dst = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_stale_dst = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_arch_dst = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_inst_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_regWen = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_src1_valid = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_phy_rs1 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_arch_rs1 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_src2_valid = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_phy_rs2 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_arch_rs2 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_rob_idx = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_imm = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_src1_value = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_src2_value = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_op1_sel = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_op2_sel = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_alu_sel = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_branch_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_uop_mem_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_52_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_52_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_52_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_52_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_52_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_52_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_52_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_52_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_52_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_52_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_53_clock = clock;
  assign reservation_station_53_reset = reset;
  assign reservation_station_53_io_i_allocated_idx = write_idx2 == 6'h35; // @[reservation_station.scala 246:65]
  assign reservation_station_53_io_i_issue_granted = (_issue1_func_code_T_53 | _issued_age_pack_issued_ages_1_T_53) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_53_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_53_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_53_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_53_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_53_io_i_write_slot = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_53_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_53_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_53_io_i_uop_valid = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_pc = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_inst = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_func_code = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_valid = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_target = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_branch_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_select = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_taken = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_phy_dst = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_stale_dst = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_arch_dst = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_inst_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_regWen = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_src1_valid = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_phy_rs1 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_arch_rs1 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_src2_valid = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_phy_rs2 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_arch_rs2 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_rob_idx = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_imm = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_src1_value = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_src2_value = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_op1_sel = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_op2_sel = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_alu_sel = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_branch_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_uop_mem_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_53_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_53_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_53_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_53_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_53_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_53_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_53_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_53_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_53_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_53_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_54_clock = clock;
  assign reservation_station_54_reset = reset;
  assign reservation_station_54_io_i_allocated_idx = write_idx2 == 6'h36; // @[reservation_station.scala 246:65]
  assign reservation_station_54_io_i_issue_granted = (_issue1_func_code_T_54 | _issued_age_pack_issued_ages_1_T_54) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_54_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_54_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_54_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_54_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_54_io_i_write_slot = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_54_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_54_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_54_io_i_uop_valid = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_pc = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_inst = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_func_code = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_valid = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_target = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_branch_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_select = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_taken = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_phy_dst = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_stale_dst = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_arch_dst = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_inst_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_regWen = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_src1_valid = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_phy_rs1 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_arch_rs1 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_src2_valid = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_phy_rs2 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_arch_rs2 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_rob_idx = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_imm = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_src1_value = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_src2_value = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_op1_sel = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_op2_sel = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_alu_sel = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_branch_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_uop_mem_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_54_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_54_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_54_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_54_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_54_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_54_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_54_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_54_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_54_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_54_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_55_clock = clock;
  assign reservation_station_55_reset = reset;
  assign reservation_station_55_io_i_allocated_idx = write_idx2 == 6'h37; // @[reservation_station.scala 246:65]
  assign reservation_station_55_io_i_issue_granted = (_issue1_func_code_T_55 | _issued_age_pack_issued_ages_1_T_55) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_55_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_55_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_55_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_55_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_55_io_i_write_slot = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_55_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_55_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_55_io_i_uop_valid = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_pc = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_inst = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_func_code = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_valid = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_target = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_branch_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_select = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_taken = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_phy_dst = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_stale_dst = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_arch_dst = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_inst_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_regWen = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_src1_valid = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_phy_rs1 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_arch_rs1 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_src2_valid = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_phy_rs2 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_arch_rs2 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_rob_idx = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_imm = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_src1_value = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_src2_value = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_op1_sel = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_op2_sel = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_alu_sel = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_branch_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_uop_mem_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_55_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_55_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_55_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_55_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_55_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_55_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_55_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_55_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_55_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_55_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_56_clock = clock;
  assign reservation_station_56_reset = reset;
  assign reservation_station_56_io_i_allocated_idx = write_idx2 == 6'h38; // @[reservation_station.scala 246:65]
  assign reservation_station_56_io_i_issue_granted = (_issue1_func_code_T_56 | _issued_age_pack_issued_ages_1_T_56) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_56_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_56_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_56_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_56_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_56_io_i_write_slot = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_56_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_56_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_56_io_i_uop_valid = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_pc = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_inst = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_func_code = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_valid = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_target = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_branch_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_select = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_taken = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_phy_dst = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_stale_dst = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_arch_dst = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_inst_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_regWen = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_src1_valid = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_phy_rs1 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_arch_rs1 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_src2_valid = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_phy_rs2 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_arch_rs2 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_rob_idx = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_imm = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_src1_value = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_src2_value = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_op1_sel = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_op2_sel = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_alu_sel = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_branch_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_uop_mem_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_56_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_56_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_56_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_56_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_56_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_56_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_56_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_56_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_56_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_56_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_57_clock = clock;
  assign reservation_station_57_reset = reset;
  assign reservation_station_57_io_i_allocated_idx = write_idx2 == 6'h39; // @[reservation_station.scala 246:65]
  assign reservation_station_57_io_i_issue_granted = (_issue1_func_code_T_57 | _issued_age_pack_issued_ages_1_T_57) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_57_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_57_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_57_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_57_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_57_io_i_write_slot = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_57_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_57_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_57_io_i_uop_valid = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_pc = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_inst = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_func_code = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_valid = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_target = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_branch_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_select = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_taken = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_phy_dst = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_stale_dst = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_arch_dst = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_inst_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_regWen = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_src1_valid = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_phy_rs1 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_arch_rs1 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_src2_valid = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_phy_rs2 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_arch_rs2 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_rob_idx = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_imm = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_src1_value = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_src2_value = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_op1_sel = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_op2_sel = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_alu_sel = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_branch_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_uop_mem_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_57_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_57_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_57_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_57_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_57_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_57_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_57_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_57_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_57_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_57_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_58_clock = clock;
  assign reservation_station_58_reset = reset;
  assign reservation_station_58_io_i_allocated_idx = write_idx2 == 6'h3a; // @[reservation_station.scala 246:65]
  assign reservation_station_58_io_i_issue_granted = (_issue1_func_code_T_58 | _issued_age_pack_issued_ages_1_T_58) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_58_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_58_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_58_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_58_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_58_io_i_write_slot = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_58_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_58_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_58_io_i_uop_valid = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_pc = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_inst = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_func_code = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_valid = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_target = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_branch_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_select = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_taken = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_phy_dst = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_stale_dst = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_arch_dst = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_inst_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_regWen = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_src1_valid = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_phy_rs1 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_arch_rs1 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_src2_valid = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_phy_rs2 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_arch_rs2 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_rob_idx = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_imm = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_src1_value = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_src2_value = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_op1_sel = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_op2_sel = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_alu_sel = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_branch_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_uop_mem_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_58_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_58_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_58_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_58_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_58_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_58_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_58_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_58_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_58_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_58_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_59_clock = clock;
  assign reservation_station_59_reset = reset;
  assign reservation_station_59_io_i_allocated_idx = write_idx2 == 6'h3b; // @[reservation_station.scala 246:65]
  assign reservation_station_59_io_i_issue_granted = (_issue1_func_code_T_59 | _issued_age_pack_issued_ages_1_T_59) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_59_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_59_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_59_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_59_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_59_io_i_write_slot = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_59_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_59_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_59_io_i_uop_valid = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_pc = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_inst = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_func_code = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_valid = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_target = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_branch_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_select = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_taken = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_phy_dst = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_stale_dst = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_arch_dst = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_inst_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_regWen = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_src1_valid = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_phy_rs1 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_arch_rs1 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_src2_valid = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_phy_rs2 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_arch_rs2 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_rob_idx = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_imm = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_src1_value = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_src2_value = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_op1_sel = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_op2_sel = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_alu_sel = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_branch_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_uop_mem_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_59_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_59_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_59_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_59_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_59_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_59_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_59_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_59_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_59_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_59_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_60_clock = clock;
  assign reservation_station_60_reset = reset;
  assign reservation_station_60_io_i_allocated_idx = write_idx2 == 6'h3c; // @[reservation_station.scala 246:65]
  assign reservation_station_60_io_i_issue_granted = (_issue1_func_code_T_60 | _issued_age_pack_issued_ages_1_T_60) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_60_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_60_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_60_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_60_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_60_io_i_write_slot = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_60_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_60_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_60_io_i_uop_valid = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_pc = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_inst = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_func_code = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_valid = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_target = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_branch_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_select = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_taken = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_phy_dst = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_stale_dst = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_arch_dst = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_inst_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_regWen = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_src1_valid = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_phy_rs1 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_arch_rs1 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_src2_valid = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_phy_rs2 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_arch_rs2 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_rob_idx = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_imm = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_src1_value = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_src2_value = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_op1_sel = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_op2_sel = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_alu_sel = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_branch_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_uop_mem_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_60_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_60_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_60_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_60_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_60_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_60_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_60_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_60_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_60_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_60_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_61_clock = clock;
  assign reservation_station_61_reset = reset;
  assign reservation_station_61_io_i_allocated_idx = write_idx2 == 6'h3d; // @[reservation_station.scala 246:65]
  assign reservation_station_61_io_i_issue_granted = (_issue1_func_code_T_61 | _issued_age_pack_issued_ages_1_T_61) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_61_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_61_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_61_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_61_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_61_io_i_write_slot = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_61_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_61_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_61_io_i_uop_valid = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_pc = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_inst = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_func_code = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_valid = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_target = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_branch_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_select = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_taken = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_phy_dst = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_stale_dst = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_arch_dst = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_inst_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_regWen = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_src1_valid = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_phy_rs1 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_arch_rs1 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_src2_valid = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_phy_rs2 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_arch_rs2 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_rob_idx = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_imm = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_src1_value = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_src2_value = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_op1_sel = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_op2_sel = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_alu_sel = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_branch_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_uop_mem_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_61_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_61_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_61_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_61_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_61_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_61_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_61_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_61_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_61_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_61_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_62_clock = clock;
  assign reservation_station_62_reset = reset;
  assign reservation_station_62_io_i_allocated_idx = write_idx2 == 6'h3e; // @[reservation_station.scala 246:65]
  assign reservation_station_62_io_i_issue_granted = (_issue1_func_code_T_62 | _issued_age_pack_issued_ages_1_T_62) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_62_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_62_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_62_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_62_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_62_io_i_write_slot = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_62_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_62_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_62_io_i_uop_valid = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_pc = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_inst = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_func_code = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_valid = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_target = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_branch_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_select = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_taken = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_phy_dst = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_stale_dst = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_arch_dst = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_inst_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_regWen = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_src1_valid = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_phy_rs1 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_arch_rs1 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_src2_valid = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_phy_rs2 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_arch_rs2 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_rob_idx = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_imm = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_src1_value = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_src2_value = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_op1_sel = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_op2_sel = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_alu_sel = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_branch_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_uop_mem_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_62_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_62_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_62_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_62_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_62_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_62_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_62_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_62_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_62_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_62_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  assign reservation_station_63_clock = clock;
  assign reservation_station_63_reset = reset;
  assign reservation_station_63_io_i_allocated_idx = write_idx2 == 6'h3f; // @[reservation_station.scala 246:65]
  assign reservation_station_63_io_i_issue_granted = (_issue1_func_code_T_63 | _issued_age_pack_issued_ages_1_T_63) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 241:94]
  assign reservation_station_63_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 242:54]
  assign reservation_station_63_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 242:54]
  assign reservation_station_63_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 242:54]
  assign reservation_station_63_io_i_exception = io_i_exception; // @[reservation_station.scala 243:44]
  assign reservation_station_63_io_i_write_slot = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_valid : _reservation_station_63_io_i_write_slot_T_1 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_63_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 244:46]
  assign reservation_station_63_io_i_uop_valid = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_pc = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_inst = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_func_code = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_valid = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_target = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_branch_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_select = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_taken = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_phy_dst = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_stale_dst = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_arch_dst = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_inst_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_regWen = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_src1_valid = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_phy_rs1 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_arch_rs1 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_src2_valid = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_phy_rs2 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_arch_rs2 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_rob_idx = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_imm = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_src1_value = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_src2_value = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_op1_sel = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_op2_sel = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_alu_sel = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_branch_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_uop_mem_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 253:44]
  assign reservation_station_63_io_i_exe_dst1 = io_i_ex_res_packs_0_valid ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 255:49]
  assign reservation_station_63_io_i_exe_dst2 = io_i_ex_res_packs_1_valid ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 256:49]
  assign reservation_station_63_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 258:45]
  assign reservation_station_63_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 259:45]
  assign reservation_station_63_io_i_age_pack_issue_valid_0 = issued_age_pack_issue_valid_0; // @[reservation_station.scala 245:42]
  assign reservation_station_63_io_i_age_pack_issue_valid_1 = issued_age_pack_issue_valid_1; // @[reservation_station.scala 245:42]
  assign reservation_station_63_io_i_age_pack_max_age = issued_age_pack_max_age; // @[reservation_station.scala 245:42]
  assign reservation_station_63_io_i_age_pack_issued_ages_0 = issued_age_pack_issued_ages_0; // @[reservation_station.scala 245:42]
  assign reservation_station_63_io_i_age_pack_issued_ages_1 = issued_age_pack_issued_ages_1; // @[reservation_station.scala 245:42]
  assign reservation_station_63_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 261:50]
  always @(posedge clock) begin
    if (reset) begin // @[reservation_station.scala 173:35]
      issued_age_pack_issue_valid_0 <= 1'h0; // @[reservation_station.scala 173:35]
    end else if (io_i_exception) begin // @[reservation_station.scala 229:26]
      issued_age_pack_issue_valid_0 <= 1'h0; // @[reservation_station.scala 230:25]
    end else begin
      issued_age_pack_issue_valid_0 <= issue0_valid; // @[reservation_station.scala 224:37]
    end
    if (reset) begin // @[reservation_station.scala 173:35]
      issued_age_pack_issue_valid_1 <= 1'h0; // @[reservation_station.scala 173:35]
    end else if (io_i_exception) begin // @[reservation_station.scala 229:26]
      issued_age_pack_issue_valid_1 <= 1'h0; // @[reservation_station.scala 230:25]
    end else begin
      issued_age_pack_issue_valid_1 <= _issue0_valid_T_1; // @[reservation_station.scala 225:37]
    end
    if (reset) begin // @[reservation_station.scala 173:35]
      issued_age_pack_max_age <= 8'h0; // @[reservation_station.scala 173:35]
    end else if (io_i_exception) begin // @[reservation_station.scala 229:26]
      issued_age_pack_max_age <= 8'h0; // @[reservation_station.scala 230:25]
    end else if (io_o_full) begin // @[reservation_station.scala 222:25]
      issued_age_pack_max_age <= max_age_temp;
    end else begin
      issued_age_pack_max_age <= 8'h3b;
    end
    if (reset) begin // @[reservation_station.scala 173:35]
      issued_age_pack_issued_ages_0 <= 8'h0; // @[reservation_station.scala 173:35]
    end else if (io_i_exception) begin // @[reservation_station.scala 229:26]
      issued_age_pack_issued_ages_0 <= 8'h0; // @[reservation_station.scala 230:25]
    end else if (_issue1_func_code_T) begin // @[Mux.scala 101:16]
      issued_age_pack_issued_ages_0 <= reservation_station_0_io_o_age;
    end else if (_issue1_func_code_T_1) begin // @[Mux.scala 101:16]
      issued_age_pack_issued_ages_0 <= reservation_station_1_io_o_age;
    end else begin
      issued_age_pack_issued_ages_0 <= _issued_age_pack_issued_ages_0_T_125;
    end
    if (reset) begin // @[reservation_station.scala 173:35]
      issued_age_pack_issued_ages_1 <= 8'h0; // @[reservation_station.scala 173:35]
    end else if (io_i_exception) begin // @[reservation_station.scala 229:26]
      issued_age_pack_issued_ages_1 <= 8'h0; // @[reservation_station.scala 230:25]
    end else if (_issued_age_pack_issued_ages_1_T) begin // @[Mux.scala 101:16]
      issued_age_pack_issued_ages_1 <= reservation_station_0_io_o_age;
    end else if (_issued_age_pack_issued_ages_1_T_1) begin // @[Mux.scala 101:16]
      issued_age_pack_issued_ages_1 <= reservation_station_1_io_o_age;
    end else begin
      issued_age_pack_issued_ages_1 <= _issued_age_pack_issued_ages_1_T_125;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  issued_age_pack_issue_valid_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  issued_age_pack_issue_valid_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  issued_age_pack_max_age = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  issued_age_pack_issued_ages_0 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  issued_age_pack_issued_ages_1 = _RAND_4[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

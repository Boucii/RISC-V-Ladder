module RegFile(
  input         clock,
  input         reset,
  input  [6:0]  io_i_raddr1,
  input  [6:0]  io_i_raddr2,
  input  [6:0]  io_i_raddr3,
  input  [6:0]  io_i_raddr4,
  output [63:0] io_o_rdata1,
  output [63:0] io_o_rdata2,
  output [63:0] io_o_rdata3,
  output [63:0] io_o_rdata4,
  input  [6:0]  io_i_waddr1,
  input  [6:0]  io_i_waddr2,
  input  [63:0] io_i_wdata1,
  input  [63:0] io_i_wdata2,
  input         io_i_wenable1,
  input         io_i_wenable2,
  output [63:0] io_o_pregs_0,
  output [63:0] io_o_pregs_1,
  output [63:0] io_o_pregs_2,
  output [63:0] io_o_pregs_3,
  output [63:0] io_o_pregs_4,
  output [63:0] io_o_pregs_5,
  output [63:0] io_o_pregs_6,
  output [63:0] io_o_pregs_7,
  output [63:0] io_o_pregs_8,
  output [63:0] io_o_pregs_9,
  output [63:0] io_o_pregs_10,
  output [63:0] io_o_pregs_11,
  output [63:0] io_o_pregs_12,
  output [63:0] io_o_pregs_13,
  output [63:0] io_o_pregs_14,
  output [63:0] io_o_pregs_15,
  output [63:0] io_o_pregs_16,
  output [63:0] io_o_pregs_17,
  output [63:0] io_o_pregs_18,
  output [63:0] io_o_pregs_19,
  output [63:0] io_o_pregs_20,
  output [63:0] io_o_pregs_21,
  output [63:0] io_o_pregs_22,
  output [63:0] io_o_pregs_23,
  output [63:0] io_o_pregs_24,
  output [63:0] io_o_pregs_25,
  output [63:0] io_o_pregs_26,
  output [63:0] io_o_pregs_27,
  output [63:0] io_o_pregs_28,
  output [63:0] io_o_pregs_29,
  output [63:0] io_o_pregs_30,
  output [63:0] io_o_pregs_31,
  output [63:0] io_o_pregs_32,
  output [63:0] io_o_pregs_33,
  output [63:0] io_o_pregs_34,
  output [63:0] io_o_pregs_35,
  output [63:0] io_o_pregs_36,
  output [63:0] io_o_pregs_37,
  output [63:0] io_o_pregs_38,
  output [63:0] io_o_pregs_39,
  output [63:0] io_o_pregs_40,
  output [63:0] io_o_pregs_41,
  output [63:0] io_o_pregs_42,
  output [63:0] io_o_pregs_43,
  output [63:0] io_o_pregs_44,
  output [63:0] io_o_pregs_45,
  output [63:0] io_o_pregs_46,
  output [63:0] io_o_pregs_47,
  output [63:0] io_o_pregs_48,
  output [63:0] io_o_pregs_49,
  output [63:0] io_o_pregs_50,
  output [63:0] io_o_pregs_51,
  output [63:0] io_o_pregs_52,
  output [63:0] io_o_pregs_53,
  output [63:0] io_o_pregs_54,
  output [63:0] io_o_pregs_55,
  output [63:0] io_o_pregs_56,
  output [63:0] io_o_pregs_57,
  output [63:0] io_o_pregs_58,
  output [63:0] io_o_pregs_59,
  output [63:0] io_o_pregs_60,
  output [63:0] io_o_pregs_61,
  output [63:0] io_o_pregs_62,
  output [63:0] io_o_pregs_63,
  output [63:0] io_o_pregs_64,
  output [63:0] io_o_pregs_65,
  output [63:0] io_o_pregs_66,
  output [63:0] io_o_pregs_67,
  output [63:0] io_o_pregs_68,
  output [63:0] io_o_pregs_69,
  output [63:0] io_o_pregs_70,
  output [63:0] io_o_pregs_71,
  output [63:0] io_o_pregs_72,
  output [63:0] io_o_pregs_73,
  output [63:0] io_o_pregs_74,
  output [63:0] io_o_pregs_75,
  output [63:0] io_o_pregs_76,
  output [63:0] io_o_pregs_77,
  output [63:0] io_o_pregs_78,
  output [63:0] io_o_pregs_79,
  output [63:0] io_o_pregs_80,
  output [63:0] io_o_pregs_81,
  output [63:0] io_o_pregs_82,
  output [63:0] io_o_pregs_83,
  output [63:0] io_o_pregs_84,
  output [63:0] io_o_pregs_85,
  output [63:0] io_o_pregs_86,
  output [63:0] io_o_pregs_87,
  output [63:0] io_o_pregs_88,
  output [63:0] io_o_pregs_89,
  output [63:0] io_o_pregs_90,
  output [63:0] io_o_pregs_91,
  output [63:0] io_o_pregs_92,
  output [63:0] io_o_pregs_93,
  output [63:0] io_o_pregs_94,
  output [63:0] io_o_pregs_95,
  output [63:0] io_o_pregs_96,
  output [63:0] io_o_pregs_97,
  output [63:0] io_o_pregs_98,
  output [63:0] io_o_pregs_99,
  output [63:0] io_o_pregs_100,
  output [63:0] io_o_pregs_101,
  output [63:0] io_o_pregs_102,
  output [63:0] io_o_pregs_103,
  output [63:0] io_o_pregs_104,
  output [63:0] io_o_pregs_105,
  output [63:0] io_o_pregs_106,
  output [63:0] io_o_pregs_107,
  output [63:0] io_o_pregs_108,
  output [63:0] io_o_pregs_109,
  output [63:0] io_o_pregs_110,
  output [63:0] io_o_pregs_111,
  output [63:0] io_o_pregs_112,
  output [63:0] io_o_pregs_113,
  output [63:0] io_o_pregs_114,
  output [63:0] io_o_pregs_115,
  output [63:0] io_o_pregs_116,
  output [63:0] io_o_pregs_117,
  output [63:0] io_o_pregs_118,
  output [63:0] io_o_pregs_119,
  output [63:0] io_o_pregs_120,
  output [63:0] io_o_pregs_121,
  output [63:0] io_o_pregs_122,
  output [63:0] io_o_pregs_123,
  output [63:0] io_o_pregs_124,
  output [63:0] io_o_pregs_125,
  output [63:0] io_o_pregs_126,
  output [63:0] io_o_pregs_127
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regfile_0; // @[regfile.scala 36:24]
  reg [63:0] regfile_1; // @[regfile.scala 36:24]
  reg [63:0] regfile_2; // @[regfile.scala 36:24]
  reg [63:0] regfile_3; // @[regfile.scala 36:24]
  reg [63:0] regfile_4; // @[regfile.scala 36:24]
  reg [63:0] regfile_5; // @[regfile.scala 36:24]
  reg [63:0] regfile_6; // @[regfile.scala 36:24]
  reg [63:0] regfile_7; // @[regfile.scala 36:24]
  reg [63:0] regfile_8; // @[regfile.scala 36:24]
  reg [63:0] regfile_9; // @[regfile.scala 36:24]
  reg [63:0] regfile_10; // @[regfile.scala 36:24]
  reg [63:0] regfile_11; // @[regfile.scala 36:24]
  reg [63:0] regfile_12; // @[regfile.scala 36:24]
  reg [63:0] regfile_13; // @[regfile.scala 36:24]
  reg [63:0] regfile_14; // @[regfile.scala 36:24]
  reg [63:0] regfile_15; // @[regfile.scala 36:24]
  reg [63:0] regfile_16; // @[regfile.scala 36:24]
  reg [63:0] regfile_17; // @[regfile.scala 36:24]
  reg [63:0] regfile_18; // @[regfile.scala 36:24]
  reg [63:0] regfile_19; // @[regfile.scala 36:24]
  reg [63:0] regfile_20; // @[regfile.scala 36:24]
  reg [63:0] regfile_21; // @[regfile.scala 36:24]
  reg [63:0] regfile_22; // @[regfile.scala 36:24]
  reg [63:0] regfile_23; // @[regfile.scala 36:24]
  reg [63:0] regfile_24; // @[regfile.scala 36:24]
  reg [63:0] regfile_25; // @[regfile.scala 36:24]
  reg [63:0] regfile_26; // @[regfile.scala 36:24]
  reg [63:0] regfile_27; // @[regfile.scala 36:24]
  reg [63:0] regfile_28; // @[regfile.scala 36:24]
  reg [63:0] regfile_29; // @[regfile.scala 36:24]
  reg [63:0] regfile_30; // @[regfile.scala 36:24]
  reg [63:0] regfile_31; // @[regfile.scala 36:24]
  reg [63:0] regfile_32; // @[regfile.scala 36:24]
  reg [63:0] regfile_33; // @[regfile.scala 36:24]
  reg [63:0] regfile_34; // @[regfile.scala 36:24]
  reg [63:0] regfile_35; // @[regfile.scala 36:24]
  reg [63:0] regfile_36; // @[regfile.scala 36:24]
  reg [63:0] regfile_37; // @[regfile.scala 36:24]
  reg [63:0] regfile_38; // @[regfile.scala 36:24]
  reg [63:0] regfile_39; // @[regfile.scala 36:24]
  reg [63:0] regfile_40; // @[regfile.scala 36:24]
  reg [63:0] regfile_41; // @[regfile.scala 36:24]
  reg [63:0] regfile_42; // @[regfile.scala 36:24]
  reg [63:0] regfile_43; // @[regfile.scala 36:24]
  reg [63:0] regfile_44; // @[regfile.scala 36:24]
  reg [63:0] regfile_45; // @[regfile.scala 36:24]
  reg [63:0] regfile_46; // @[regfile.scala 36:24]
  reg [63:0] regfile_47; // @[regfile.scala 36:24]
  reg [63:0] regfile_48; // @[regfile.scala 36:24]
  reg [63:0] regfile_49; // @[regfile.scala 36:24]
  reg [63:0] regfile_50; // @[regfile.scala 36:24]
  reg [63:0] regfile_51; // @[regfile.scala 36:24]
  reg [63:0] regfile_52; // @[regfile.scala 36:24]
  reg [63:0] regfile_53; // @[regfile.scala 36:24]
  reg [63:0] regfile_54; // @[regfile.scala 36:24]
  reg [63:0] regfile_55; // @[regfile.scala 36:24]
  reg [63:0] regfile_56; // @[regfile.scala 36:24]
  reg [63:0] regfile_57; // @[regfile.scala 36:24]
  reg [63:0] regfile_58; // @[regfile.scala 36:24]
  reg [63:0] regfile_59; // @[regfile.scala 36:24]
  reg [63:0] regfile_60; // @[regfile.scala 36:24]
  reg [63:0] regfile_61; // @[regfile.scala 36:24]
  reg [63:0] regfile_62; // @[regfile.scala 36:24]
  reg [63:0] regfile_63; // @[regfile.scala 36:24]
  reg [63:0] regfile_64; // @[regfile.scala 36:24]
  reg [63:0] regfile_65; // @[regfile.scala 36:24]
  reg [63:0] regfile_66; // @[regfile.scala 36:24]
  reg [63:0] regfile_67; // @[regfile.scala 36:24]
  reg [63:0] regfile_68; // @[regfile.scala 36:24]
  reg [63:0] regfile_69; // @[regfile.scala 36:24]
  reg [63:0] regfile_70; // @[regfile.scala 36:24]
  reg [63:0] regfile_71; // @[regfile.scala 36:24]
  reg [63:0] regfile_72; // @[regfile.scala 36:24]
  reg [63:0] regfile_73; // @[regfile.scala 36:24]
  reg [63:0] regfile_74; // @[regfile.scala 36:24]
  reg [63:0] regfile_75; // @[regfile.scala 36:24]
  reg [63:0] regfile_76; // @[regfile.scala 36:24]
  reg [63:0] regfile_77; // @[regfile.scala 36:24]
  reg [63:0] regfile_78; // @[regfile.scala 36:24]
  reg [63:0] regfile_79; // @[regfile.scala 36:24]
  reg [63:0] regfile_80; // @[regfile.scala 36:24]
  reg [63:0] regfile_81; // @[regfile.scala 36:24]
  reg [63:0] regfile_82; // @[regfile.scala 36:24]
  reg [63:0] regfile_83; // @[regfile.scala 36:24]
  reg [63:0] regfile_84; // @[regfile.scala 36:24]
  reg [63:0] regfile_85; // @[regfile.scala 36:24]
  reg [63:0] regfile_86; // @[regfile.scala 36:24]
  reg [63:0] regfile_87; // @[regfile.scala 36:24]
  reg [63:0] regfile_88; // @[regfile.scala 36:24]
  reg [63:0] regfile_89; // @[regfile.scala 36:24]
  reg [63:0] regfile_90; // @[regfile.scala 36:24]
  reg [63:0] regfile_91; // @[regfile.scala 36:24]
  reg [63:0] regfile_92; // @[regfile.scala 36:24]
  reg [63:0] regfile_93; // @[regfile.scala 36:24]
  reg [63:0] regfile_94; // @[regfile.scala 36:24]
  reg [63:0] regfile_95; // @[regfile.scala 36:24]
  reg [63:0] regfile_96; // @[regfile.scala 36:24]
  reg [63:0] regfile_97; // @[regfile.scala 36:24]
  reg [63:0] regfile_98; // @[regfile.scala 36:24]
  reg [63:0] regfile_99; // @[regfile.scala 36:24]
  reg [63:0] regfile_100; // @[regfile.scala 36:24]
  reg [63:0] regfile_101; // @[regfile.scala 36:24]
  reg [63:0] regfile_102; // @[regfile.scala 36:24]
  reg [63:0] regfile_103; // @[regfile.scala 36:24]
  reg [63:0] regfile_104; // @[regfile.scala 36:24]
  reg [63:0] regfile_105; // @[regfile.scala 36:24]
  reg [63:0] regfile_106; // @[regfile.scala 36:24]
  reg [63:0] regfile_107; // @[regfile.scala 36:24]
  reg [63:0] regfile_108; // @[regfile.scala 36:24]
  reg [63:0] regfile_109; // @[regfile.scala 36:24]
  reg [63:0] regfile_110; // @[regfile.scala 36:24]
  reg [63:0] regfile_111; // @[regfile.scala 36:24]
  reg [63:0] regfile_112; // @[regfile.scala 36:24]
  reg [63:0] regfile_113; // @[regfile.scala 36:24]
  reg [63:0] regfile_114; // @[regfile.scala 36:24]
  reg [63:0] regfile_115; // @[regfile.scala 36:24]
  reg [63:0] regfile_116; // @[regfile.scala 36:24]
  reg [63:0] regfile_117; // @[regfile.scala 36:24]
  reg [63:0] regfile_118; // @[regfile.scala 36:24]
  reg [63:0] regfile_119; // @[regfile.scala 36:24]
  reg [63:0] regfile_120; // @[regfile.scala 36:24]
  reg [63:0] regfile_121; // @[regfile.scala 36:24]
  reg [63:0] regfile_122; // @[regfile.scala 36:24]
  reg [63:0] regfile_123; // @[regfile.scala 36:24]
  reg [63:0] regfile_124; // @[regfile.scala 36:24]
  reg [63:0] regfile_125; // @[regfile.scala 36:24]
  reg [63:0] regfile_126; // @[regfile.scala 36:24]
  reg [63:0] regfile_127; // @[regfile.scala 36:24]
  wire [63:0] _GEN_0 = 7'h0 == io_i_waddr1 ? io_i_wdata1 : regfile_0; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_1 = 7'h1 == io_i_waddr1 ? io_i_wdata1 : regfile_1; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_2 = 7'h2 == io_i_waddr1 ? io_i_wdata1 : regfile_2; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_3 = 7'h3 == io_i_waddr1 ? io_i_wdata1 : regfile_3; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_4 = 7'h4 == io_i_waddr1 ? io_i_wdata1 : regfile_4; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_5 = 7'h5 == io_i_waddr1 ? io_i_wdata1 : regfile_5; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_6 = 7'h6 == io_i_waddr1 ? io_i_wdata1 : regfile_6; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_7 = 7'h7 == io_i_waddr1 ? io_i_wdata1 : regfile_7; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_8 = 7'h8 == io_i_waddr1 ? io_i_wdata1 : regfile_8; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_9 = 7'h9 == io_i_waddr1 ? io_i_wdata1 : regfile_9; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_10 = 7'ha == io_i_waddr1 ? io_i_wdata1 : regfile_10; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_11 = 7'hb == io_i_waddr1 ? io_i_wdata1 : regfile_11; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_12 = 7'hc == io_i_waddr1 ? io_i_wdata1 : regfile_12; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_13 = 7'hd == io_i_waddr1 ? io_i_wdata1 : regfile_13; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_14 = 7'he == io_i_waddr1 ? io_i_wdata1 : regfile_14; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_15 = 7'hf == io_i_waddr1 ? io_i_wdata1 : regfile_15; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_16 = 7'h10 == io_i_waddr1 ? io_i_wdata1 : regfile_16; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_17 = 7'h11 == io_i_waddr1 ? io_i_wdata1 : regfile_17; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_18 = 7'h12 == io_i_waddr1 ? io_i_wdata1 : regfile_18; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_19 = 7'h13 == io_i_waddr1 ? io_i_wdata1 : regfile_19; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_20 = 7'h14 == io_i_waddr1 ? io_i_wdata1 : regfile_20; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_21 = 7'h15 == io_i_waddr1 ? io_i_wdata1 : regfile_21; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_22 = 7'h16 == io_i_waddr1 ? io_i_wdata1 : regfile_22; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_23 = 7'h17 == io_i_waddr1 ? io_i_wdata1 : regfile_23; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_24 = 7'h18 == io_i_waddr1 ? io_i_wdata1 : regfile_24; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_25 = 7'h19 == io_i_waddr1 ? io_i_wdata1 : regfile_25; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_26 = 7'h1a == io_i_waddr1 ? io_i_wdata1 : regfile_26; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_27 = 7'h1b == io_i_waddr1 ? io_i_wdata1 : regfile_27; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_28 = 7'h1c == io_i_waddr1 ? io_i_wdata1 : regfile_28; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_29 = 7'h1d == io_i_waddr1 ? io_i_wdata1 : regfile_29; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_30 = 7'h1e == io_i_waddr1 ? io_i_wdata1 : regfile_30; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_31 = 7'h1f == io_i_waddr1 ? io_i_wdata1 : regfile_31; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_32 = 7'h20 == io_i_waddr1 ? io_i_wdata1 : regfile_32; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_33 = 7'h21 == io_i_waddr1 ? io_i_wdata1 : regfile_33; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_34 = 7'h22 == io_i_waddr1 ? io_i_wdata1 : regfile_34; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_35 = 7'h23 == io_i_waddr1 ? io_i_wdata1 : regfile_35; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_36 = 7'h24 == io_i_waddr1 ? io_i_wdata1 : regfile_36; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_37 = 7'h25 == io_i_waddr1 ? io_i_wdata1 : regfile_37; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_38 = 7'h26 == io_i_waddr1 ? io_i_wdata1 : regfile_38; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_39 = 7'h27 == io_i_waddr1 ? io_i_wdata1 : regfile_39; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_40 = 7'h28 == io_i_waddr1 ? io_i_wdata1 : regfile_40; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_41 = 7'h29 == io_i_waddr1 ? io_i_wdata1 : regfile_41; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_42 = 7'h2a == io_i_waddr1 ? io_i_wdata1 : regfile_42; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_43 = 7'h2b == io_i_waddr1 ? io_i_wdata1 : regfile_43; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_44 = 7'h2c == io_i_waddr1 ? io_i_wdata1 : regfile_44; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_45 = 7'h2d == io_i_waddr1 ? io_i_wdata1 : regfile_45; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_46 = 7'h2e == io_i_waddr1 ? io_i_wdata1 : regfile_46; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_47 = 7'h2f == io_i_waddr1 ? io_i_wdata1 : regfile_47; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_48 = 7'h30 == io_i_waddr1 ? io_i_wdata1 : regfile_48; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_49 = 7'h31 == io_i_waddr1 ? io_i_wdata1 : regfile_49; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_50 = 7'h32 == io_i_waddr1 ? io_i_wdata1 : regfile_50; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_51 = 7'h33 == io_i_waddr1 ? io_i_wdata1 : regfile_51; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_52 = 7'h34 == io_i_waddr1 ? io_i_wdata1 : regfile_52; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_53 = 7'h35 == io_i_waddr1 ? io_i_wdata1 : regfile_53; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_54 = 7'h36 == io_i_waddr1 ? io_i_wdata1 : regfile_54; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_55 = 7'h37 == io_i_waddr1 ? io_i_wdata1 : regfile_55; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_56 = 7'h38 == io_i_waddr1 ? io_i_wdata1 : regfile_56; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_57 = 7'h39 == io_i_waddr1 ? io_i_wdata1 : regfile_57; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_58 = 7'h3a == io_i_waddr1 ? io_i_wdata1 : regfile_58; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_59 = 7'h3b == io_i_waddr1 ? io_i_wdata1 : regfile_59; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_60 = 7'h3c == io_i_waddr1 ? io_i_wdata1 : regfile_60; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_61 = 7'h3d == io_i_waddr1 ? io_i_wdata1 : regfile_61; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_62 = 7'h3e == io_i_waddr1 ? io_i_wdata1 : regfile_62; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_63 = 7'h3f == io_i_waddr1 ? io_i_wdata1 : regfile_63; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_64 = 7'h40 == io_i_waddr1 ? io_i_wdata1 : regfile_64; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_65 = 7'h41 == io_i_waddr1 ? io_i_wdata1 : regfile_65; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_66 = 7'h42 == io_i_waddr1 ? io_i_wdata1 : regfile_66; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_67 = 7'h43 == io_i_waddr1 ? io_i_wdata1 : regfile_67; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_68 = 7'h44 == io_i_waddr1 ? io_i_wdata1 : regfile_68; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_69 = 7'h45 == io_i_waddr1 ? io_i_wdata1 : regfile_69; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_70 = 7'h46 == io_i_waddr1 ? io_i_wdata1 : regfile_70; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_71 = 7'h47 == io_i_waddr1 ? io_i_wdata1 : regfile_71; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_72 = 7'h48 == io_i_waddr1 ? io_i_wdata1 : regfile_72; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_73 = 7'h49 == io_i_waddr1 ? io_i_wdata1 : regfile_73; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_74 = 7'h4a == io_i_waddr1 ? io_i_wdata1 : regfile_74; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_75 = 7'h4b == io_i_waddr1 ? io_i_wdata1 : regfile_75; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_76 = 7'h4c == io_i_waddr1 ? io_i_wdata1 : regfile_76; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_77 = 7'h4d == io_i_waddr1 ? io_i_wdata1 : regfile_77; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_78 = 7'h4e == io_i_waddr1 ? io_i_wdata1 : regfile_78; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_79 = 7'h4f == io_i_waddr1 ? io_i_wdata1 : regfile_79; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_80 = 7'h50 == io_i_waddr1 ? io_i_wdata1 : regfile_80; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_81 = 7'h51 == io_i_waddr1 ? io_i_wdata1 : regfile_81; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_82 = 7'h52 == io_i_waddr1 ? io_i_wdata1 : regfile_82; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_83 = 7'h53 == io_i_waddr1 ? io_i_wdata1 : regfile_83; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_84 = 7'h54 == io_i_waddr1 ? io_i_wdata1 : regfile_84; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_85 = 7'h55 == io_i_waddr1 ? io_i_wdata1 : regfile_85; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_86 = 7'h56 == io_i_waddr1 ? io_i_wdata1 : regfile_86; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_87 = 7'h57 == io_i_waddr1 ? io_i_wdata1 : regfile_87; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_88 = 7'h58 == io_i_waddr1 ? io_i_wdata1 : regfile_88; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_89 = 7'h59 == io_i_waddr1 ? io_i_wdata1 : regfile_89; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_90 = 7'h5a == io_i_waddr1 ? io_i_wdata1 : regfile_90; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_91 = 7'h5b == io_i_waddr1 ? io_i_wdata1 : regfile_91; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_92 = 7'h5c == io_i_waddr1 ? io_i_wdata1 : regfile_92; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_93 = 7'h5d == io_i_waddr1 ? io_i_wdata1 : regfile_93; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_94 = 7'h5e == io_i_waddr1 ? io_i_wdata1 : regfile_94; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_95 = 7'h5f == io_i_waddr1 ? io_i_wdata1 : regfile_95; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_96 = 7'h60 == io_i_waddr1 ? io_i_wdata1 : regfile_96; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_97 = 7'h61 == io_i_waddr1 ? io_i_wdata1 : regfile_97; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_98 = 7'h62 == io_i_waddr1 ? io_i_wdata1 : regfile_98; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_99 = 7'h63 == io_i_waddr1 ? io_i_wdata1 : regfile_99; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_100 = 7'h64 == io_i_waddr1 ? io_i_wdata1 : regfile_100; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_101 = 7'h65 == io_i_waddr1 ? io_i_wdata1 : regfile_101; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_102 = 7'h66 == io_i_waddr1 ? io_i_wdata1 : regfile_102; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_103 = 7'h67 == io_i_waddr1 ? io_i_wdata1 : regfile_103; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_104 = 7'h68 == io_i_waddr1 ? io_i_wdata1 : regfile_104; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_105 = 7'h69 == io_i_waddr1 ? io_i_wdata1 : regfile_105; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_106 = 7'h6a == io_i_waddr1 ? io_i_wdata1 : regfile_106; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_107 = 7'h6b == io_i_waddr1 ? io_i_wdata1 : regfile_107; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_108 = 7'h6c == io_i_waddr1 ? io_i_wdata1 : regfile_108; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_109 = 7'h6d == io_i_waddr1 ? io_i_wdata1 : regfile_109; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_110 = 7'h6e == io_i_waddr1 ? io_i_wdata1 : regfile_110; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_111 = 7'h6f == io_i_waddr1 ? io_i_wdata1 : regfile_111; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_112 = 7'h70 == io_i_waddr1 ? io_i_wdata1 : regfile_112; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_113 = 7'h71 == io_i_waddr1 ? io_i_wdata1 : regfile_113; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_114 = 7'h72 == io_i_waddr1 ? io_i_wdata1 : regfile_114; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_115 = 7'h73 == io_i_waddr1 ? io_i_wdata1 : regfile_115; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_116 = 7'h74 == io_i_waddr1 ? io_i_wdata1 : regfile_116; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_117 = 7'h75 == io_i_waddr1 ? io_i_wdata1 : regfile_117; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_118 = 7'h76 == io_i_waddr1 ? io_i_wdata1 : regfile_118; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_119 = 7'h77 == io_i_waddr1 ? io_i_wdata1 : regfile_119; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_120 = 7'h78 == io_i_waddr1 ? io_i_wdata1 : regfile_120; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_121 = 7'h79 == io_i_waddr1 ? io_i_wdata1 : regfile_121; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_122 = 7'h7a == io_i_waddr1 ? io_i_wdata1 : regfile_122; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_123 = 7'h7b == io_i_waddr1 ? io_i_wdata1 : regfile_123; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_124 = 7'h7c == io_i_waddr1 ? io_i_wdata1 : regfile_124; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_125 = 7'h7d == io_i_waddr1 ? io_i_wdata1 : regfile_125; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_126 = 7'h7e == io_i_waddr1 ? io_i_wdata1 : regfile_126; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_127 = 7'h7f == io_i_waddr1 ? io_i_wdata1 : regfile_127; // @[regfile.scala 36:24 44:{26,26}]
  wire [63:0] _GEN_128 = io_i_wenable1 ? _GEN_0 : regfile_0; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_129 = io_i_wenable1 ? _GEN_1 : regfile_1; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_130 = io_i_wenable1 ? _GEN_2 : regfile_2; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_131 = io_i_wenable1 ? _GEN_3 : regfile_3; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_132 = io_i_wenable1 ? _GEN_4 : regfile_4; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_133 = io_i_wenable1 ? _GEN_5 : regfile_5; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_134 = io_i_wenable1 ? _GEN_6 : regfile_6; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_135 = io_i_wenable1 ? _GEN_7 : regfile_7; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_136 = io_i_wenable1 ? _GEN_8 : regfile_8; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_137 = io_i_wenable1 ? _GEN_9 : regfile_9; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_138 = io_i_wenable1 ? _GEN_10 : regfile_10; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_139 = io_i_wenable1 ? _GEN_11 : regfile_11; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_140 = io_i_wenable1 ? _GEN_12 : regfile_12; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_141 = io_i_wenable1 ? _GEN_13 : regfile_13; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_142 = io_i_wenable1 ? _GEN_14 : regfile_14; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_143 = io_i_wenable1 ? _GEN_15 : regfile_15; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_144 = io_i_wenable1 ? _GEN_16 : regfile_16; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_145 = io_i_wenable1 ? _GEN_17 : regfile_17; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_146 = io_i_wenable1 ? _GEN_18 : regfile_18; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_147 = io_i_wenable1 ? _GEN_19 : regfile_19; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_148 = io_i_wenable1 ? _GEN_20 : regfile_20; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_149 = io_i_wenable1 ? _GEN_21 : regfile_21; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_150 = io_i_wenable1 ? _GEN_22 : regfile_22; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_151 = io_i_wenable1 ? _GEN_23 : regfile_23; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_152 = io_i_wenable1 ? _GEN_24 : regfile_24; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_153 = io_i_wenable1 ? _GEN_25 : regfile_25; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_154 = io_i_wenable1 ? _GEN_26 : regfile_26; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_155 = io_i_wenable1 ? _GEN_27 : regfile_27; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_156 = io_i_wenable1 ? _GEN_28 : regfile_28; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_157 = io_i_wenable1 ? _GEN_29 : regfile_29; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_158 = io_i_wenable1 ? _GEN_30 : regfile_30; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_159 = io_i_wenable1 ? _GEN_31 : regfile_31; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_160 = io_i_wenable1 ? _GEN_32 : regfile_32; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_161 = io_i_wenable1 ? _GEN_33 : regfile_33; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_162 = io_i_wenable1 ? _GEN_34 : regfile_34; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_163 = io_i_wenable1 ? _GEN_35 : regfile_35; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_164 = io_i_wenable1 ? _GEN_36 : regfile_36; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_165 = io_i_wenable1 ? _GEN_37 : regfile_37; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_166 = io_i_wenable1 ? _GEN_38 : regfile_38; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_167 = io_i_wenable1 ? _GEN_39 : regfile_39; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_168 = io_i_wenable1 ? _GEN_40 : regfile_40; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_169 = io_i_wenable1 ? _GEN_41 : regfile_41; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_170 = io_i_wenable1 ? _GEN_42 : regfile_42; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_171 = io_i_wenable1 ? _GEN_43 : regfile_43; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_172 = io_i_wenable1 ? _GEN_44 : regfile_44; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_173 = io_i_wenable1 ? _GEN_45 : regfile_45; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_174 = io_i_wenable1 ? _GEN_46 : regfile_46; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_175 = io_i_wenable1 ? _GEN_47 : regfile_47; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_176 = io_i_wenable1 ? _GEN_48 : regfile_48; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_177 = io_i_wenable1 ? _GEN_49 : regfile_49; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_178 = io_i_wenable1 ? _GEN_50 : regfile_50; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_179 = io_i_wenable1 ? _GEN_51 : regfile_51; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_180 = io_i_wenable1 ? _GEN_52 : regfile_52; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_181 = io_i_wenable1 ? _GEN_53 : regfile_53; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_182 = io_i_wenable1 ? _GEN_54 : regfile_54; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_183 = io_i_wenable1 ? _GEN_55 : regfile_55; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_184 = io_i_wenable1 ? _GEN_56 : regfile_56; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_185 = io_i_wenable1 ? _GEN_57 : regfile_57; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_186 = io_i_wenable1 ? _GEN_58 : regfile_58; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_187 = io_i_wenable1 ? _GEN_59 : regfile_59; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_188 = io_i_wenable1 ? _GEN_60 : regfile_60; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_189 = io_i_wenable1 ? _GEN_61 : regfile_61; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_190 = io_i_wenable1 ? _GEN_62 : regfile_62; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_191 = io_i_wenable1 ? _GEN_63 : regfile_63; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_192 = io_i_wenable1 ? _GEN_64 : regfile_64; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_193 = io_i_wenable1 ? _GEN_65 : regfile_65; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_194 = io_i_wenable1 ? _GEN_66 : regfile_66; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_195 = io_i_wenable1 ? _GEN_67 : regfile_67; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_196 = io_i_wenable1 ? _GEN_68 : regfile_68; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_197 = io_i_wenable1 ? _GEN_69 : regfile_69; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_198 = io_i_wenable1 ? _GEN_70 : regfile_70; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_199 = io_i_wenable1 ? _GEN_71 : regfile_71; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_200 = io_i_wenable1 ? _GEN_72 : regfile_72; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_201 = io_i_wenable1 ? _GEN_73 : regfile_73; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_202 = io_i_wenable1 ? _GEN_74 : regfile_74; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_203 = io_i_wenable1 ? _GEN_75 : regfile_75; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_204 = io_i_wenable1 ? _GEN_76 : regfile_76; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_205 = io_i_wenable1 ? _GEN_77 : regfile_77; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_206 = io_i_wenable1 ? _GEN_78 : regfile_78; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_207 = io_i_wenable1 ? _GEN_79 : regfile_79; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_208 = io_i_wenable1 ? _GEN_80 : regfile_80; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_209 = io_i_wenable1 ? _GEN_81 : regfile_81; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_210 = io_i_wenable1 ? _GEN_82 : regfile_82; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_211 = io_i_wenable1 ? _GEN_83 : regfile_83; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_212 = io_i_wenable1 ? _GEN_84 : regfile_84; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_213 = io_i_wenable1 ? _GEN_85 : regfile_85; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_214 = io_i_wenable1 ? _GEN_86 : regfile_86; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_215 = io_i_wenable1 ? _GEN_87 : regfile_87; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_216 = io_i_wenable1 ? _GEN_88 : regfile_88; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_217 = io_i_wenable1 ? _GEN_89 : regfile_89; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_218 = io_i_wenable1 ? _GEN_90 : regfile_90; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_219 = io_i_wenable1 ? _GEN_91 : regfile_91; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_220 = io_i_wenable1 ? _GEN_92 : regfile_92; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_221 = io_i_wenable1 ? _GEN_93 : regfile_93; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_222 = io_i_wenable1 ? _GEN_94 : regfile_94; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_223 = io_i_wenable1 ? _GEN_95 : regfile_95; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_224 = io_i_wenable1 ? _GEN_96 : regfile_96; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_225 = io_i_wenable1 ? _GEN_97 : regfile_97; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_226 = io_i_wenable1 ? _GEN_98 : regfile_98; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_227 = io_i_wenable1 ? _GEN_99 : regfile_99; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_228 = io_i_wenable1 ? _GEN_100 : regfile_100; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_229 = io_i_wenable1 ? _GEN_101 : regfile_101; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_230 = io_i_wenable1 ? _GEN_102 : regfile_102; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_231 = io_i_wenable1 ? _GEN_103 : regfile_103; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_232 = io_i_wenable1 ? _GEN_104 : regfile_104; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_233 = io_i_wenable1 ? _GEN_105 : regfile_105; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_234 = io_i_wenable1 ? _GEN_106 : regfile_106; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_235 = io_i_wenable1 ? _GEN_107 : regfile_107; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_236 = io_i_wenable1 ? _GEN_108 : regfile_108; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_237 = io_i_wenable1 ? _GEN_109 : regfile_109; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_238 = io_i_wenable1 ? _GEN_110 : regfile_110; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_239 = io_i_wenable1 ? _GEN_111 : regfile_111; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_240 = io_i_wenable1 ? _GEN_112 : regfile_112; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_241 = io_i_wenable1 ? _GEN_113 : regfile_113; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_242 = io_i_wenable1 ? _GEN_114 : regfile_114; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_243 = io_i_wenable1 ? _GEN_115 : regfile_115; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_244 = io_i_wenable1 ? _GEN_116 : regfile_116; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_245 = io_i_wenable1 ? _GEN_117 : regfile_117; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_246 = io_i_wenable1 ? _GEN_118 : regfile_118; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_247 = io_i_wenable1 ? _GEN_119 : regfile_119; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_248 = io_i_wenable1 ? _GEN_120 : regfile_120; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_249 = io_i_wenable1 ? _GEN_121 : regfile_121; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_250 = io_i_wenable1 ? _GEN_122 : regfile_122; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_251 = io_i_wenable1 ? _GEN_123 : regfile_123; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_252 = io_i_wenable1 ? _GEN_124 : regfile_124; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_253 = io_i_wenable1 ? _GEN_125 : regfile_125; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_254 = io_i_wenable1 ? _GEN_126 : regfile_126; // @[regfile.scala 43:23 36:24]
  wire [63:0] _GEN_255 = io_i_wenable1 ? _GEN_127 : regfile_127; // @[regfile.scala 43:23 36:24]
  wire  _io_o_rdata1_T_1 = io_i_wenable1 & io_i_waddr1 == io_i_raddr1; // @[regfile.scala 52:20]
  wire  _io_o_rdata1_T_3 = io_i_wenable2 & io_i_waddr2 == io_i_raddr1; // @[regfile.scala 53:20]
  wire [63:0] _GEN_513 = 7'h1 == io_i_raddr1 ? regfile_1 : regfile_0; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_514 = 7'h2 == io_i_raddr1 ? regfile_2 : _GEN_513; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_515 = 7'h3 == io_i_raddr1 ? regfile_3 : _GEN_514; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_516 = 7'h4 == io_i_raddr1 ? regfile_4 : _GEN_515; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_517 = 7'h5 == io_i_raddr1 ? regfile_5 : _GEN_516; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_518 = 7'h6 == io_i_raddr1 ? regfile_6 : _GEN_517; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_519 = 7'h7 == io_i_raddr1 ? regfile_7 : _GEN_518; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_520 = 7'h8 == io_i_raddr1 ? regfile_8 : _GEN_519; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_521 = 7'h9 == io_i_raddr1 ? regfile_9 : _GEN_520; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_522 = 7'ha == io_i_raddr1 ? regfile_10 : _GEN_521; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_523 = 7'hb == io_i_raddr1 ? regfile_11 : _GEN_522; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_524 = 7'hc == io_i_raddr1 ? regfile_12 : _GEN_523; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_525 = 7'hd == io_i_raddr1 ? regfile_13 : _GEN_524; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_526 = 7'he == io_i_raddr1 ? regfile_14 : _GEN_525; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_527 = 7'hf == io_i_raddr1 ? regfile_15 : _GEN_526; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_528 = 7'h10 == io_i_raddr1 ? regfile_16 : _GEN_527; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_529 = 7'h11 == io_i_raddr1 ? regfile_17 : _GEN_528; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_530 = 7'h12 == io_i_raddr1 ? regfile_18 : _GEN_529; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_531 = 7'h13 == io_i_raddr1 ? regfile_19 : _GEN_530; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_532 = 7'h14 == io_i_raddr1 ? regfile_20 : _GEN_531; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_533 = 7'h15 == io_i_raddr1 ? regfile_21 : _GEN_532; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_534 = 7'h16 == io_i_raddr1 ? regfile_22 : _GEN_533; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_535 = 7'h17 == io_i_raddr1 ? regfile_23 : _GEN_534; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_536 = 7'h18 == io_i_raddr1 ? regfile_24 : _GEN_535; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_537 = 7'h19 == io_i_raddr1 ? regfile_25 : _GEN_536; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_538 = 7'h1a == io_i_raddr1 ? regfile_26 : _GEN_537; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_539 = 7'h1b == io_i_raddr1 ? regfile_27 : _GEN_538; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_540 = 7'h1c == io_i_raddr1 ? regfile_28 : _GEN_539; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_541 = 7'h1d == io_i_raddr1 ? regfile_29 : _GEN_540; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_542 = 7'h1e == io_i_raddr1 ? regfile_30 : _GEN_541; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_543 = 7'h1f == io_i_raddr1 ? regfile_31 : _GEN_542; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_544 = 7'h20 == io_i_raddr1 ? regfile_32 : _GEN_543; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_545 = 7'h21 == io_i_raddr1 ? regfile_33 : _GEN_544; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_546 = 7'h22 == io_i_raddr1 ? regfile_34 : _GEN_545; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_547 = 7'h23 == io_i_raddr1 ? regfile_35 : _GEN_546; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_548 = 7'h24 == io_i_raddr1 ? regfile_36 : _GEN_547; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_549 = 7'h25 == io_i_raddr1 ? regfile_37 : _GEN_548; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_550 = 7'h26 == io_i_raddr1 ? regfile_38 : _GEN_549; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_551 = 7'h27 == io_i_raddr1 ? regfile_39 : _GEN_550; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_552 = 7'h28 == io_i_raddr1 ? regfile_40 : _GEN_551; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_553 = 7'h29 == io_i_raddr1 ? regfile_41 : _GEN_552; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_554 = 7'h2a == io_i_raddr1 ? regfile_42 : _GEN_553; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_555 = 7'h2b == io_i_raddr1 ? regfile_43 : _GEN_554; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_556 = 7'h2c == io_i_raddr1 ? regfile_44 : _GEN_555; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_557 = 7'h2d == io_i_raddr1 ? regfile_45 : _GEN_556; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_558 = 7'h2e == io_i_raddr1 ? regfile_46 : _GEN_557; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_559 = 7'h2f == io_i_raddr1 ? regfile_47 : _GEN_558; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_560 = 7'h30 == io_i_raddr1 ? regfile_48 : _GEN_559; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_561 = 7'h31 == io_i_raddr1 ? regfile_49 : _GEN_560; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_562 = 7'h32 == io_i_raddr1 ? regfile_50 : _GEN_561; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_563 = 7'h33 == io_i_raddr1 ? regfile_51 : _GEN_562; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_564 = 7'h34 == io_i_raddr1 ? regfile_52 : _GEN_563; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_565 = 7'h35 == io_i_raddr1 ? regfile_53 : _GEN_564; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_566 = 7'h36 == io_i_raddr1 ? regfile_54 : _GEN_565; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_567 = 7'h37 == io_i_raddr1 ? regfile_55 : _GEN_566; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_568 = 7'h38 == io_i_raddr1 ? regfile_56 : _GEN_567; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_569 = 7'h39 == io_i_raddr1 ? regfile_57 : _GEN_568; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_570 = 7'h3a == io_i_raddr1 ? regfile_58 : _GEN_569; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_571 = 7'h3b == io_i_raddr1 ? regfile_59 : _GEN_570; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_572 = 7'h3c == io_i_raddr1 ? regfile_60 : _GEN_571; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_573 = 7'h3d == io_i_raddr1 ? regfile_61 : _GEN_572; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_574 = 7'h3e == io_i_raddr1 ? regfile_62 : _GEN_573; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_575 = 7'h3f == io_i_raddr1 ? regfile_63 : _GEN_574; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_576 = 7'h40 == io_i_raddr1 ? regfile_64 : _GEN_575; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_577 = 7'h41 == io_i_raddr1 ? regfile_65 : _GEN_576; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_578 = 7'h42 == io_i_raddr1 ? regfile_66 : _GEN_577; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_579 = 7'h43 == io_i_raddr1 ? regfile_67 : _GEN_578; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_580 = 7'h44 == io_i_raddr1 ? regfile_68 : _GEN_579; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_581 = 7'h45 == io_i_raddr1 ? regfile_69 : _GEN_580; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_582 = 7'h46 == io_i_raddr1 ? regfile_70 : _GEN_581; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_583 = 7'h47 == io_i_raddr1 ? regfile_71 : _GEN_582; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_584 = 7'h48 == io_i_raddr1 ? regfile_72 : _GEN_583; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_585 = 7'h49 == io_i_raddr1 ? regfile_73 : _GEN_584; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_586 = 7'h4a == io_i_raddr1 ? regfile_74 : _GEN_585; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_587 = 7'h4b == io_i_raddr1 ? regfile_75 : _GEN_586; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_588 = 7'h4c == io_i_raddr1 ? regfile_76 : _GEN_587; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_589 = 7'h4d == io_i_raddr1 ? regfile_77 : _GEN_588; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_590 = 7'h4e == io_i_raddr1 ? regfile_78 : _GEN_589; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_591 = 7'h4f == io_i_raddr1 ? regfile_79 : _GEN_590; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_592 = 7'h50 == io_i_raddr1 ? regfile_80 : _GEN_591; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_593 = 7'h51 == io_i_raddr1 ? regfile_81 : _GEN_592; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_594 = 7'h52 == io_i_raddr1 ? regfile_82 : _GEN_593; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_595 = 7'h53 == io_i_raddr1 ? regfile_83 : _GEN_594; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_596 = 7'h54 == io_i_raddr1 ? regfile_84 : _GEN_595; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_597 = 7'h55 == io_i_raddr1 ? regfile_85 : _GEN_596; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_598 = 7'h56 == io_i_raddr1 ? regfile_86 : _GEN_597; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_599 = 7'h57 == io_i_raddr1 ? regfile_87 : _GEN_598; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_600 = 7'h58 == io_i_raddr1 ? regfile_88 : _GEN_599; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_601 = 7'h59 == io_i_raddr1 ? regfile_89 : _GEN_600; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_602 = 7'h5a == io_i_raddr1 ? regfile_90 : _GEN_601; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_603 = 7'h5b == io_i_raddr1 ? regfile_91 : _GEN_602; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_604 = 7'h5c == io_i_raddr1 ? regfile_92 : _GEN_603; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_605 = 7'h5d == io_i_raddr1 ? regfile_93 : _GEN_604; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_606 = 7'h5e == io_i_raddr1 ? regfile_94 : _GEN_605; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_607 = 7'h5f == io_i_raddr1 ? regfile_95 : _GEN_606; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_608 = 7'h60 == io_i_raddr1 ? regfile_96 : _GEN_607; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_609 = 7'h61 == io_i_raddr1 ? regfile_97 : _GEN_608; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_610 = 7'h62 == io_i_raddr1 ? regfile_98 : _GEN_609; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_611 = 7'h63 == io_i_raddr1 ? regfile_99 : _GEN_610; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_612 = 7'h64 == io_i_raddr1 ? regfile_100 : _GEN_611; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_613 = 7'h65 == io_i_raddr1 ? regfile_101 : _GEN_612; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_614 = 7'h66 == io_i_raddr1 ? regfile_102 : _GEN_613; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_615 = 7'h67 == io_i_raddr1 ? regfile_103 : _GEN_614; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_616 = 7'h68 == io_i_raddr1 ? regfile_104 : _GEN_615; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_617 = 7'h69 == io_i_raddr1 ? regfile_105 : _GEN_616; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_618 = 7'h6a == io_i_raddr1 ? regfile_106 : _GEN_617; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_619 = 7'h6b == io_i_raddr1 ? regfile_107 : _GEN_618; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_620 = 7'h6c == io_i_raddr1 ? regfile_108 : _GEN_619; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_621 = 7'h6d == io_i_raddr1 ? regfile_109 : _GEN_620; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_622 = 7'h6e == io_i_raddr1 ? regfile_110 : _GEN_621; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_623 = 7'h6f == io_i_raddr1 ? regfile_111 : _GEN_622; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_624 = 7'h70 == io_i_raddr1 ? regfile_112 : _GEN_623; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_625 = 7'h71 == io_i_raddr1 ? regfile_113 : _GEN_624; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_626 = 7'h72 == io_i_raddr1 ? regfile_114 : _GEN_625; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_627 = 7'h73 == io_i_raddr1 ? regfile_115 : _GEN_626; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_628 = 7'h74 == io_i_raddr1 ? regfile_116 : _GEN_627; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_629 = 7'h75 == io_i_raddr1 ? regfile_117 : _GEN_628; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_630 = 7'h76 == io_i_raddr1 ? regfile_118 : _GEN_629; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_631 = 7'h77 == io_i_raddr1 ? regfile_119 : _GEN_630; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_632 = 7'h78 == io_i_raddr1 ? regfile_120 : _GEN_631; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_633 = 7'h79 == io_i_raddr1 ? regfile_121 : _GEN_632; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_634 = 7'h7a == io_i_raddr1 ? regfile_122 : _GEN_633; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_635 = 7'h7b == io_i_raddr1 ? regfile_123 : _GEN_634; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_636 = 7'h7c == io_i_raddr1 ? regfile_124 : _GEN_635; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_637 = 7'h7d == io_i_raddr1 ? regfile_125 : _GEN_636; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_638 = 7'h7e == io_i_raddr1 ? regfile_126 : _GEN_637; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_639 = 7'h7f == io_i_raddr1 ? regfile_127 : _GEN_638; // @[Mux.scala 101:{16,16}]
  wire [63:0] _io_o_rdata1_T_4 = _io_o_rdata1_T_3 ? io_i_wdata2 : _GEN_639; // @[Mux.scala 101:16]
  wire  _io_o_rdata2_T_1 = io_i_wenable1 & io_i_waddr1 == io_i_raddr2; // @[regfile.scala 56:20]
  wire  _io_o_rdata2_T_3 = io_i_wenable2 & io_i_waddr2 == io_i_raddr2; // @[regfile.scala 57:20]
  wire [63:0] _GEN_641 = 7'h1 == io_i_raddr2 ? regfile_1 : regfile_0; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_642 = 7'h2 == io_i_raddr2 ? regfile_2 : _GEN_641; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_643 = 7'h3 == io_i_raddr2 ? regfile_3 : _GEN_642; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_644 = 7'h4 == io_i_raddr2 ? regfile_4 : _GEN_643; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_645 = 7'h5 == io_i_raddr2 ? regfile_5 : _GEN_644; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_646 = 7'h6 == io_i_raddr2 ? regfile_6 : _GEN_645; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_647 = 7'h7 == io_i_raddr2 ? regfile_7 : _GEN_646; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_648 = 7'h8 == io_i_raddr2 ? regfile_8 : _GEN_647; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_649 = 7'h9 == io_i_raddr2 ? regfile_9 : _GEN_648; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_650 = 7'ha == io_i_raddr2 ? regfile_10 : _GEN_649; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_651 = 7'hb == io_i_raddr2 ? regfile_11 : _GEN_650; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_652 = 7'hc == io_i_raddr2 ? regfile_12 : _GEN_651; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_653 = 7'hd == io_i_raddr2 ? regfile_13 : _GEN_652; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_654 = 7'he == io_i_raddr2 ? regfile_14 : _GEN_653; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_655 = 7'hf == io_i_raddr2 ? regfile_15 : _GEN_654; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_656 = 7'h10 == io_i_raddr2 ? regfile_16 : _GEN_655; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_657 = 7'h11 == io_i_raddr2 ? regfile_17 : _GEN_656; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_658 = 7'h12 == io_i_raddr2 ? regfile_18 : _GEN_657; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_659 = 7'h13 == io_i_raddr2 ? regfile_19 : _GEN_658; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_660 = 7'h14 == io_i_raddr2 ? regfile_20 : _GEN_659; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_661 = 7'h15 == io_i_raddr2 ? regfile_21 : _GEN_660; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_662 = 7'h16 == io_i_raddr2 ? regfile_22 : _GEN_661; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_663 = 7'h17 == io_i_raddr2 ? regfile_23 : _GEN_662; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_664 = 7'h18 == io_i_raddr2 ? regfile_24 : _GEN_663; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_665 = 7'h19 == io_i_raddr2 ? regfile_25 : _GEN_664; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_666 = 7'h1a == io_i_raddr2 ? regfile_26 : _GEN_665; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_667 = 7'h1b == io_i_raddr2 ? regfile_27 : _GEN_666; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_668 = 7'h1c == io_i_raddr2 ? regfile_28 : _GEN_667; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_669 = 7'h1d == io_i_raddr2 ? regfile_29 : _GEN_668; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_670 = 7'h1e == io_i_raddr2 ? regfile_30 : _GEN_669; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_671 = 7'h1f == io_i_raddr2 ? regfile_31 : _GEN_670; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_672 = 7'h20 == io_i_raddr2 ? regfile_32 : _GEN_671; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_673 = 7'h21 == io_i_raddr2 ? regfile_33 : _GEN_672; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_674 = 7'h22 == io_i_raddr2 ? regfile_34 : _GEN_673; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_675 = 7'h23 == io_i_raddr2 ? regfile_35 : _GEN_674; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_676 = 7'h24 == io_i_raddr2 ? regfile_36 : _GEN_675; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_677 = 7'h25 == io_i_raddr2 ? regfile_37 : _GEN_676; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_678 = 7'h26 == io_i_raddr2 ? regfile_38 : _GEN_677; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_679 = 7'h27 == io_i_raddr2 ? regfile_39 : _GEN_678; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_680 = 7'h28 == io_i_raddr2 ? regfile_40 : _GEN_679; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_681 = 7'h29 == io_i_raddr2 ? regfile_41 : _GEN_680; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_682 = 7'h2a == io_i_raddr2 ? regfile_42 : _GEN_681; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_683 = 7'h2b == io_i_raddr2 ? regfile_43 : _GEN_682; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_684 = 7'h2c == io_i_raddr2 ? regfile_44 : _GEN_683; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_685 = 7'h2d == io_i_raddr2 ? regfile_45 : _GEN_684; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_686 = 7'h2e == io_i_raddr2 ? regfile_46 : _GEN_685; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_687 = 7'h2f == io_i_raddr2 ? regfile_47 : _GEN_686; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_688 = 7'h30 == io_i_raddr2 ? regfile_48 : _GEN_687; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_689 = 7'h31 == io_i_raddr2 ? regfile_49 : _GEN_688; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_690 = 7'h32 == io_i_raddr2 ? regfile_50 : _GEN_689; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_691 = 7'h33 == io_i_raddr2 ? regfile_51 : _GEN_690; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_692 = 7'h34 == io_i_raddr2 ? regfile_52 : _GEN_691; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_693 = 7'h35 == io_i_raddr2 ? regfile_53 : _GEN_692; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_694 = 7'h36 == io_i_raddr2 ? regfile_54 : _GEN_693; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_695 = 7'h37 == io_i_raddr2 ? regfile_55 : _GEN_694; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_696 = 7'h38 == io_i_raddr2 ? regfile_56 : _GEN_695; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_697 = 7'h39 == io_i_raddr2 ? regfile_57 : _GEN_696; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_698 = 7'h3a == io_i_raddr2 ? regfile_58 : _GEN_697; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_699 = 7'h3b == io_i_raddr2 ? regfile_59 : _GEN_698; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_700 = 7'h3c == io_i_raddr2 ? regfile_60 : _GEN_699; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_701 = 7'h3d == io_i_raddr2 ? regfile_61 : _GEN_700; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_702 = 7'h3e == io_i_raddr2 ? regfile_62 : _GEN_701; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_703 = 7'h3f == io_i_raddr2 ? regfile_63 : _GEN_702; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_704 = 7'h40 == io_i_raddr2 ? regfile_64 : _GEN_703; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_705 = 7'h41 == io_i_raddr2 ? regfile_65 : _GEN_704; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_706 = 7'h42 == io_i_raddr2 ? regfile_66 : _GEN_705; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_707 = 7'h43 == io_i_raddr2 ? regfile_67 : _GEN_706; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_708 = 7'h44 == io_i_raddr2 ? regfile_68 : _GEN_707; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_709 = 7'h45 == io_i_raddr2 ? regfile_69 : _GEN_708; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_710 = 7'h46 == io_i_raddr2 ? regfile_70 : _GEN_709; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_711 = 7'h47 == io_i_raddr2 ? regfile_71 : _GEN_710; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_712 = 7'h48 == io_i_raddr2 ? regfile_72 : _GEN_711; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_713 = 7'h49 == io_i_raddr2 ? regfile_73 : _GEN_712; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_714 = 7'h4a == io_i_raddr2 ? regfile_74 : _GEN_713; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_715 = 7'h4b == io_i_raddr2 ? regfile_75 : _GEN_714; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_716 = 7'h4c == io_i_raddr2 ? regfile_76 : _GEN_715; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_717 = 7'h4d == io_i_raddr2 ? regfile_77 : _GEN_716; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_718 = 7'h4e == io_i_raddr2 ? regfile_78 : _GEN_717; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_719 = 7'h4f == io_i_raddr2 ? regfile_79 : _GEN_718; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_720 = 7'h50 == io_i_raddr2 ? regfile_80 : _GEN_719; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_721 = 7'h51 == io_i_raddr2 ? regfile_81 : _GEN_720; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_722 = 7'h52 == io_i_raddr2 ? regfile_82 : _GEN_721; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_723 = 7'h53 == io_i_raddr2 ? regfile_83 : _GEN_722; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_724 = 7'h54 == io_i_raddr2 ? regfile_84 : _GEN_723; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_725 = 7'h55 == io_i_raddr2 ? regfile_85 : _GEN_724; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_726 = 7'h56 == io_i_raddr2 ? regfile_86 : _GEN_725; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_727 = 7'h57 == io_i_raddr2 ? regfile_87 : _GEN_726; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_728 = 7'h58 == io_i_raddr2 ? regfile_88 : _GEN_727; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_729 = 7'h59 == io_i_raddr2 ? regfile_89 : _GEN_728; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_730 = 7'h5a == io_i_raddr2 ? regfile_90 : _GEN_729; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_731 = 7'h5b == io_i_raddr2 ? regfile_91 : _GEN_730; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_732 = 7'h5c == io_i_raddr2 ? regfile_92 : _GEN_731; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_733 = 7'h5d == io_i_raddr2 ? regfile_93 : _GEN_732; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_734 = 7'h5e == io_i_raddr2 ? regfile_94 : _GEN_733; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_735 = 7'h5f == io_i_raddr2 ? regfile_95 : _GEN_734; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_736 = 7'h60 == io_i_raddr2 ? regfile_96 : _GEN_735; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_737 = 7'h61 == io_i_raddr2 ? regfile_97 : _GEN_736; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_738 = 7'h62 == io_i_raddr2 ? regfile_98 : _GEN_737; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_739 = 7'h63 == io_i_raddr2 ? regfile_99 : _GEN_738; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_740 = 7'h64 == io_i_raddr2 ? regfile_100 : _GEN_739; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_741 = 7'h65 == io_i_raddr2 ? regfile_101 : _GEN_740; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_742 = 7'h66 == io_i_raddr2 ? regfile_102 : _GEN_741; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_743 = 7'h67 == io_i_raddr2 ? regfile_103 : _GEN_742; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_744 = 7'h68 == io_i_raddr2 ? regfile_104 : _GEN_743; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_745 = 7'h69 == io_i_raddr2 ? regfile_105 : _GEN_744; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_746 = 7'h6a == io_i_raddr2 ? regfile_106 : _GEN_745; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_747 = 7'h6b == io_i_raddr2 ? regfile_107 : _GEN_746; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_748 = 7'h6c == io_i_raddr2 ? regfile_108 : _GEN_747; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_749 = 7'h6d == io_i_raddr2 ? regfile_109 : _GEN_748; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_750 = 7'h6e == io_i_raddr2 ? regfile_110 : _GEN_749; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_751 = 7'h6f == io_i_raddr2 ? regfile_111 : _GEN_750; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_752 = 7'h70 == io_i_raddr2 ? regfile_112 : _GEN_751; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_753 = 7'h71 == io_i_raddr2 ? regfile_113 : _GEN_752; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_754 = 7'h72 == io_i_raddr2 ? regfile_114 : _GEN_753; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_755 = 7'h73 == io_i_raddr2 ? regfile_115 : _GEN_754; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_756 = 7'h74 == io_i_raddr2 ? regfile_116 : _GEN_755; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_757 = 7'h75 == io_i_raddr2 ? regfile_117 : _GEN_756; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_758 = 7'h76 == io_i_raddr2 ? regfile_118 : _GEN_757; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_759 = 7'h77 == io_i_raddr2 ? regfile_119 : _GEN_758; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_760 = 7'h78 == io_i_raddr2 ? regfile_120 : _GEN_759; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_761 = 7'h79 == io_i_raddr2 ? regfile_121 : _GEN_760; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_762 = 7'h7a == io_i_raddr2 ? regfile_122 : _GEN_761; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_763 = 7'h7b == io_i_raddr2 ? regfile_123 : _GEN_762; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_764 = 7'h7c == io_i_raddr2 ? regfile_124 : _GEN_763; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_765 = 7'h7d == io_i_raddr2 ? regfile_125 : _GEN_764; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_766 = 7'h7e == io_i_raddr2 ? regfile_126 : _GEN_765; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_767 = 7'h7f == io_i_raddr2 ? regfile_127 : _GEN_766; // @[Mux.scala 101:{16,16}]
  wire [63:0] _io_o_rdata2_T_4 = _io_o_rdata2_T_3 ? io_i_wdata2 : _GEN_767; // @[Mux.scala 101:16]
  wire  _io_o_rdata3_T_1 = io_i_wenable1 & io_i_waddr1 == io_i_raddr3; // @[regfile.scala 60:20]
  wire  _io_o_rdata3_T_3 = io_i_wenable2 & io_i_waddr2 == io_i_raddr3; // @[regfile.scala 61:20]
  wire [63:0] _GEN_769 = 7'h1 == io_i_raddr3 ? regfile_1 : regfile_0; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_770 = 7'h2 == io_i_raddr3 ? regfile_2 : _GEN_769; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_771 = 7'h3 == io_i_raddr3 ? regfile_3 : _GEN_770; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_772 = 7'h4 == io_i_raddr3 ? regfile_4 : _GEN_771; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_773 = 7'h5 == io_i_raddr3 ? regfile_5 : _GEN_772; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_774 = 7'h6 == io_i_raddr3 ? regfile_6 : _GEN_773; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_775 = 7'h7 == io_i_raddr3 ? regfile_7 : _GEN_774; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_776 = 7'h8 == io_i_raddr3 ? regfile_8 : _GEN_775; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_777 = 7'h9 == io_i_raddr3 ? regfile_9 : _GEN_776; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_778 = 7'ha == io_i_raddr3 ? regfile_10 : _GEN_777; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_779 = 7'hb == io_i_raddr3 ? regfile_11 : _GEN_778; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_780 = 7'hc == io_i_raddr3 ? regfile_12 : _GEN_779; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_781 = 7'hd == io_i_raddr3 ? regfile_13 : _GEN_780; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_782 = 7'he == io_i_raddr3 ? regfile_14 : _GEN_781; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_783 = 7'hf == io_i_raddr3 ? regfile_15 : _GEN_782; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_784 = 7'h10 == io_i_raddr3 ? regfile_16 : _GEN_783; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_785 = 7'h11 == io_i_raddr3 ? regfile_17 : _GEN_784; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_786 = 7'h12 == io_i_raddr3 ? regfile_18 : _GEN_785; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_787 = 7'h13 == io_i_raddr3 ? regfile_19 : _GEN_786; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_788 = 7'h14 == io_i_raddr3 ? regfile_20 : _GEN_787; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_789 = 7'h15 == io_i_raddr3 ? regfile_21 : _GEN_788; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_790 = 7'h16 == io_i_raddr3 ? regfile_22 : _GEN_789; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_791 = 7'h17 == io_i_raddr3 ? regfile_23 : _GEN_790; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_792 = 7'h18 == io_i_raddr3 ? regfile_24 : _GEN_791; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_793 = 7'h19 == io_i_raddr3 ? regfile_25 : _GEN_792; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_794 = 7'h1a == io_i_raddr3 ? regfile_26 : _GEN_793; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_795 = 7'h1b == io_i_raddr3 ? regfile_27 : _GEN_794; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_796 = 7'h1c == io_i_raddr3 ? regfile_28 : _GEN_795; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_797 = 7'h1d == io_i_raddr3 ? regfile_29 : _GEN_796; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_798 = 7'h1e == io_i_raddr3 ? regfile_30 : _GEN_797; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_799 = 7'h1f == io_i_raddr3 ? regfile_31 : _GEN_798; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_800 = 7'h20 == io_i_raddr3 ? regfile_32 : _GEN_799; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_801 = 7'h21 == io_i_raddr3 ? regfile_33 : _GEN_800; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_802 = 7'h22 == io_i_raddr3 ? regfile_34 : _GEN_801; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_803 = 7'h23 == io_i_raddr3 ? regfile_35 : _GEN_802; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_804 = 7'h24 == io_i_raddr3 ? regfile_36 : _GEN_803; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_805 = 7'h25 == io_i_raddr3 ? regfile_37 : _GEN_804; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_806 = 7'h26 == io_i_raddr3 ? regfile_38 : _GEN_805; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_807 = 7'h27 == io_i_raddr3 ? regfile_39 : _GEN_806; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_808 = 7'h28 == io_i_raddr3 ? regfile_40 : _GEN_807; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_809 = 7'h29 == io_i_raddr3 ? regfile_41 : _GEN_808; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_810 = 7'h2a == io_i_raddr3 ? regfile_42 : _GEN_809; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_811 = 7'h2b == io_i_raddr3 ? regfile_43 : _GEN_810; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_812 = 7'h2c == io_i_raddr3 ? regfile_44 : _GEN_811; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_813 = 7'h2d == io_i_raddr3 ? regfile_45 : _GEN_812; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_814 = 7'h2e == io_i_raddr3 ? regfile_46 : _GEN_813; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_815 = 7'h2f == io_i_raddr3 ? regfile_47 : _GEN_814; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_816 = 7'h30 == io_i_raddr3 ? regfile_48 : _GEN_815; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_817 = 7'h31 == io_i_raddr3 ? regfile_49 : _GEN_816; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_818 = 7'h32 == io_i_raddr3 ? regfile_50 : _GEN_817; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_819 = 7'h33 == io_i_raddr3 ? regfile_51 : _GEN_818; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_820 = 7'h34 == io_i_raddr3 ? regfile_52 : _GEN_819; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_821 = 7'h35 == io_i_raddr3 ? regfile_53 : _GEN_820; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_822 = 7'h36 == io_i_raddr3 ? regfile_54 : _GEN_821; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_823 = 7'h37 == io_i_raddr3 ? regfile_55 : _GEN_822; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_824 = 7'h38 == io_i_raddr3 ? regfile_56 : _GEN_823; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_825 = 7'h39 == io_i_raddr3 ? regfile_57 : _GEN_824; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_826 = 7'h3a == io_i_raddr3 ? regfile_58 : _GEN_825; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_827 = 7'h3b == io_i_raddr3 ? regfile_59 : _GEN_826; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_828 = 7'h3c == io_i_raddr3 ? regfile_60 : _GEN_827; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_829 = 7'h3d == io_i_raddr3 ? regfile_61 : _GEN_828; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_830 = 7'h3e == io_i_raddr3 ? regfile_62 : _GEN_829; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_831 = 7'h3f == io_i_raddr3 ? regfile_63 : _GEN_830; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_832 = 7'h40 == io_i_raddr3 ? regfile_64 : _GEN_831; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_833 = 7'h41 == io_i_raddr3 ? regfile_65 : _GEN_832; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_834 = 7'h42 == io_i_raddr3 ? regfile_66 : _GEN_833; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_835 = 7'h43 == io_i_raddr3 ? regfile_67 : _GEN_834; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_836 = 7'h44 == io_i_raddr3 ? regfile_68 : _GEN_835; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_837 = 7'h45 == io_i_raddr3 ? regfile_69 : _GEN_836; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_838 = 7'h46 == io_i_raddr3 ? regfile_70 : _GEN_837; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_839 = 7'h47 == io_i_raddr3 ? regfile_71 : _GEN_838; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_840 = 7'h48 == io_i_raddr3 ? regfile_72 : _GEN_839; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_841 = 7'h49 == io_i_raddr3 ? regfile_73 : _GEN_840; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_842 = 7'h4a == io_i_raddr3 ? regfile_74 : _GEN_841; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_843 = 7'h4b == io_i_raddr3 ? regfile_75 : _GEN_842; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_844 = 7'h4c == io_i_raddr3 ? regfile_76 : _GEN_843; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_845 = 7'h4d == io_i_raddr3 ? regfile_77 : _GEN_844; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_846 = 7'h4e == io_i_raddr3 ? regfile_78 : _GEN_845; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_847 = 7'h4f == io_i_raddr3 ? regfile_79 : _GEN_846; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_848 = 7'h50 == io_i_raddr3 ? regfile_80 : _GEN_847; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_849 = 7'h51 == io_i_raddr3 ? regfile_81 : _GEN_848; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_850 = 7'h52 == io_i_raddr3 ? regfile_82 : _GEN_849; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_851 = 7'h53 == io_i_raddr3 ? regfile_83 : _GEN_850; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_852 = 7'h54 == io_i_raddr3 ? regfile_84 : _GEN_851; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_853 = 7'h55 == io_i_raddr3 ? regfile_85 : _GEN_852; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_854 = 7'h56 == io_i_raddr3 ? regfile_86 : _GEN_853; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_855 = 7'h57 == io_i_raddr3 ? regfile_87 : _GEN_854; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_856 = 7'h58 == io_i_raddr3 ? regfile_88 : _GEN_855; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_857 = 7'h59 == io_i_raddr3 ? regfile_89 : _GEN_856; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_858 = 7'h5a == io_i_raddr3 ? regfile_90 : _GEN_857; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_859 = 7'h5b == io_i_raddr3 ? regfile_91 : _GEN_858; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_860 = 7'h5c == io_i_raddr3 ? regfile_92 : _GEN_859; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_861 = 7'h5d == io_i_raddr3 ? regfile_93 : _GEN_860; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_862 = 7'h5e == io_i_raddr3 ? regfile_94 : _GEN_861; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_863 = 7'h5f == io_i_raddr3 ? regfile_95 : _GEN_862; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_864 = 7'h60 == io_i_raddr3 ? regfile_96 : _GEN_863; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_865 = 7'h61 == io_i_raddr3 ? regfile_97 : _GEN_864; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_866 = 7'h62 == io_i_raddr3 ? regfile_98 : _GEN_865; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_867 = 7'h63 == io_i_raddr3 ? regfile_99 : _GEN_866; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_868 = 7'h64 == io_i_raddr3 ? regfile_100 : _GEN_867; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_869 = 7'h65 == io_i_raddr3 ? regfile_101 : _GEN_868; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_870 = 7'h66 == io_i_raddr3 ? regfile_102 : _GEN_869; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_871 = 7'h67 == io_i_raddr3 ? regfile_103 : _GEN_870; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_872 = 7'h68 == io_i_raddr3 ? regfile_104 : _GEN_871; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_873 = 7'h69 == io_i_raddr3 ? regfile_105 : _GEN_872; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_874 = 7'h6a == io_i_raddr3 ? regfile_106 : _GEN_873; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_875 = 7'h6b == io_i_raddr3 ? regfile_107 : _GEN_874; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_876 = 7'h6c == io_i_raddr3 ? regfile_108 : _GEN_875; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_877 = 7'h6d == io_i_raddr3 ? regfile_109 : _GEN_876; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_878 = 7'h6e == io_i_raddr3 ? regfile_110 : _GEN_877; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_879 = 7'h6f == io_i_raddr3 ? regfile_111 : _GEN_878; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_880 = 7'h70 == io_i_raddr3 ? regfile_112 : _GEN_879; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_881 = 7'h71 == io_i_raddr3 ? regfile_113 : _GEN_880; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_882 = 7'h72 == io_i_raddr3 ? regfile_114 : _GEN_881; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_883 = 7'h73 == io_i_raddr3 ? regfile_115 : _GEN_882; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_884 = 7'h74 == io_i_raddr3 ? regfile_116 : _GEN_883; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_885 = 7'h75 == io_i_raddr3 ? regfile_117 : _GEN_884; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_886 = 7'h76 == io_i_raddr3 ? regfile_118 : _GEN_885; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_887 = 7'h77 == io_i_raddr3 ? regfile_119 : _GEN_886; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_888 = 7'h78 == io_i_raddr3 ? regfile_120 : _GEN_887; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_889 = 7'h79 == io_i_raddr3 ? regfile_121 : _GEN_888; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_890 = 7'h7a == io_i_raddr3 ? regfile_122 : _GEN_889; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_891 = 7'h7b == io_i_raddr3 ? regfile_123 : _GEN_890; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_892 = 7'h7c == io_i_raddr3 ? regfile_124 : _GEN_891; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_893 = 7'h7d == io_i_raddr3 ? regfile_125 : _GEN_892; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_894 = 7'h7e == io_i_raddr3 ? regfile_126 : _GEN_893; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_895 = 7'h7f == io_i_raddr3 ? regfile_127 : _GEN_894; // @[Mux.scala 101:{16,16}]
  wire [63:0] _io_o_rdata3_T_4 = _io_o_rdata3_T_3 ? io_i_wdata2 : _GEN_895; // @[Mux.scala 101:16]
  wire  _io_o_rdata4_T_1 = io_i_wenable1 & io_i_waddr1 == io_i_raddr4; // @[regfile.scala 64:20]
  wire  _io_o_rdata4_T_3 = io_i_wenable2 & io_i_waddr2 == io_i_raddr4; // @[regfile.scala 65:20]
  wire [63:0] _GEN_897 = 7'h1 == io_i_raddr4 ? regfile_1 : regfile_0; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_898 = 7'h2 == io_i_raddr4 ? regfile_2 : _GEN_897; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_899 = 7'h3 == io_i_raddr4 ? regfile_3 : _GEN_898; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_900 = 7'h4 == io_i_raddr4 ? regfile_4 : _GEN_899; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_901 = 7'h5 == io_i_raddr4 ? regfile_5 : _GEN_900; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_902 = 7'h6 == io_i_raddr4 ? regfile_6 : _GEN_901; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_903 = 7'h7 == io_i_raddr4 ? regfile_7 : _GEN_902; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_904 = 7'h8 == io_i_raddr4 ? regfile_8 : _GEN_903; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_905 = 7'h9 == io_i_raddr4 ? regfile_9 : _GEN_904; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_906 = 7'ha == io_i_raddr4 ? regfile_10 : _GEN_905; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_907 = 7'hb == io_i_raddr4 ? regfile_11 : _GEN_906; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_908 = 7'hc == io_i_raddr4 ? regfile_12 : _GEN_907; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_909 = 7'hd == io_i_raddr4 ? regfile_13 : _GEN_908; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_910 = 7'he == io_i_raddr4 ? regfile_14 : _GEN_909; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_911 = 7'hf == io_i_raddr4 ? regfile_15 : _GEN_910; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_912 = 7'h10 == io_i_raddr4 ? regfile_16 : _GEN_911; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_913 = 7'h11 == io_i_raddr4 ? regfile_17 : _GEN_912; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_914 = 7'h12 == io_i_raddr4 ? regfile_18 : _GEN_913; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_915 = 7'h13 == io_i_raddr4 ? regfile_19 : _GEN_914; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_916 = 7'h14 == io_i_raddr4 ? regfile_20 : _GEN_915; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_917 = 7'h15 == io_i_raddr4 ? regfile_21 : _GEN_916; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_918 = 7'h16 == io_i_raddr4 ? regfile_22 : _GEN_917; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_919 = 7'h17 == io_i_raddr4 ? regfile_23 : _GEN_918; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_920 = 7'h18 == io_i_raddr4 ? regfile_24 : _GEN_919; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_921 = 7'h19 == io_i_raddr4 ? regfile_25 : _GEN_920; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_922 = 7'h1a == io_i_raddr4 ? regfile_26 : _GEN_921; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_923 = 7'h1b == io_i_raddr4 ? regfile_27 : _GEN_922; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_924 = 7'h1c == io_i_raddr4 ? regfile_28 : _GEN_923; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_925 = 7'h1d == io_i_raddr4 ? regfile_29 : _GEN_924; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_926 = 7'h1e == io_i_raddr4 ? regfile_30 : _GEN_925; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_927 = 7'h1f == io_i_raddr4 ? regfile_31 : _GEN_926; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_928 = 7'h20 == io_i_raddr4 ? regfile_32 : _GEN_927; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_929 = 7'h21 == io_i_raddr4 ? regfile_33 : _GEN_928; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_930 = 7'h22 == io_i_raddr4 ? regfile_34 : _GEN_929; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_931 = 7'h23 == io_i_raddr4 ? regfile_35 : _GEN_930; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_932 = 7'h24 == io_i_raddr4 ? regfile_36 : _GEN_931; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_933 = 7'h25 == io_i_raddr4 ? regfile_37 : _GEN_932; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_934 = 7'h26 == io_i_raddr4 ? regfile_38 : _GEN_933; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_935 = 7'h27 == io_i_raddr4 ? regfile_39 : _GEN_934; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_936 = 7'h28 == io_i_raddr4 ? regfile_40 : _GEN_935; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_937 = 7'h29 == io_i_raddr4 ? regfile_41 : _GEN_936; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_938 = 7'h2a == io_i_raddr4 ? regfile_42 : _GEN_937; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_939 = 7'h2b == io_i_raddr4 ? regfile_43 : _GEN_938; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_940 = 7'h2c == io_i_raddr4 ? regfile_44 : _GEN_939; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_941 = 7'h2d == io_i_raddr4 ? regfile_45 : _GEN_940; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_942 = 7'h2e == io_i_raddr4 ? regfile_46 : _GEN_941; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_943 = 7'h2f == io_i_raddr4 ? regfile_47 : _GEN_942; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_944 = 7'h30 == io_i_raddr4 ? regfile_48 : _GEN_943; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_945 = 7'h31 == io_i_raddr4 ? regfile_49 : _GEN_944; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_946 = 7'h32 == io_i_raddr4 ? regfile_50 : _GEN_945; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_947 = 7'h33 == io_i_raddr4 ? regfile_51 : _GEN_946; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_948 = 7'h34 == io_i_raddr4 ? regfile_52 : _GEN_947; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_949 = 7'h35 == io_i_raddr4 ? regfile_53 : _GEN_948; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_950 = 7'h36 == io_i_raddr4 ? regfile_54 : _GEN_949; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_951 = 7'h37 == io_i_raddr4 ? regfile_55 : _GEN_950; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_952 = 7'h38 == io_i_raddr4 ? regfile_56 : _GEN_951; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_953 = 7'h39 == io_i_raddr4 ? regfile_57 : _GEN_952; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_954 = 7'h3a == io_i_raddr4 ? regfile_58 : _GEN_953; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_955 = 7'h3b == io_i_raddr4 ? regfile_59 : _GEN_954; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_956 = 7'h3c == io_i_raddr4 ? regfile_60 : _GEN_955; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_957 = 7'h3d == io_i_raddr4 ? regfile_61 : _GEN_956; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_958 = 7'h3e == io_i_raddr4 ? regfile_62 : _GEN_957; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_959 = 7'h3f == io_i_raddr4 ? regfile_63 : _GEN_958; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_960 = 7'h40 == io_i_raddr4 ? regfile_64 : _GEN_959; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_961 = 7'h41 == io_i_raddr4 ? regfile_65 : _GEN_960; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_962 = 7'h42 == io_i_raddr4 ? regfile_66 : _GEN_961; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_963 = 7'h43 == io_i_raddr4 ? regfile_67 : _GEN_962; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_964 = 7'h44 == io_i_raddr4 ? regfile_68 : _GEN_963; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_965 = 7'h45 == io_i_raddr4 ? regfile_69 : _GEN_964; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_966 = 7'h46 == io_i_raddr4 ? regfile_70 : _GEN_965; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_967 = 7'h47 == io_i_raddr4 ? regfile_71 : _GEN_966; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_968 = 7'h48 == io_i_raddr4 ? regfile_72 : _GEN_967; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_969 = 7'h49 == io_i_raddr4 ? regfile_73 : _GEN_968; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_970 = 7'h4a == io_i_raddr4 ? regfile_74 : _GEN_969; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_971 = 7'h4b == io_i_raddr4 ? regfile_75 : _GEN_970; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_972 = 7'h4c == io_i_raddr4 ? regfile_76 : _GEN_971; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_973 = 7'h4d == io_i_raddr4 ? regfile_77 : _GEN_972; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_974 = 7'h4e == io_i_raddr4 ? regfile_78 : _GEN_973; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_975 = 7'h4f == io_i_raddr4 ? regfile_79 : _GEN_974; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_976 = 7'h50 == io_i_raddr4 ? regfile_80 : _GEN_975; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_977 = 7'h51 == io_i_raddr4 ? regfile_81 : _GEN_976; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_978 = 7'h52 == io_i_raddr4 ? regfile_82 : _GEN_977; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_979 = 7'h53 == io_i_raddr4 ? regfile_83 : _GEN_978; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_980 = 7'h54 == io_i_raddr4 ? regfile_84 : _GEN_979; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_981 = 7'h55 == io_i_raddr4 ? regfile_85 : _GEN_980; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_982 = 7'h56 == io_i_raddr4 ? regfile_86 : _GEN_981; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_983 = 7'h57 == io_i_raddr4 ? regfile_87 : _GEN_982; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_984 = 7'h58 == io_i_raddr4 ? regfile_88 : _GEN_983; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_985 = 7'h59 == io_i_raddr4 ? regfile_89 : _GEN_984; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_986 = 7'h5a == io_i_raddr4 ? regfile_90 : _GEN_985; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_987 = 7'h5b == io_i_raddr4 ? regfile_91 : _GEN_986; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_988 = 7'h5c == io_i_raddr4 ? regfile_92 : _GEN_987; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_989 = 7'h5d == io_i_raddr4 ? regfile_93 : _GEN_988; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_990 = 7'h5e == io_i_raddr4 ? regfile_94 : _GEN_989; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_991 = 7'h5f == io_i_raddr4 ? regfile_95 : _GEN_990; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_992 = 7'h60 == io_i_raddr4 ? regfile_96 : _GEN_991; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_993 = 7'h61 == io_i_raddr4 ? regfile_97 : _GEN_992; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_994 = 7'h62 == io_i_raddr4 ? regfile_98 : _GEN_993; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_995 = 7'h63 == io_i_raddr4 ? regfile_99 : _GEN_994; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_996 = 7'h64 == io_i_raddr4 ? regfile_100 : _GEN_995; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_997 = 7'h65 == io_i_raddr4 ? regfile_101 : _GEN_996; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_998 = 7'h66 == io_i_raddr4 ? regfile_102 : _GEN_997; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_999 = 7'h67 == io_i_raddr4 ? regfile_103 : _GEN_998; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1000 = 7'h68 == io_i_raddr4 ? regfile_104 : _GEN_999; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1001 = 7'h69 == io_i_raddr4 ? regfile_105 : _GEN_1000; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1002 = 7'h6a == io_i_raddr4 ? regfile_106 : _GEN_1001; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1003 = 7'h6b == io_i_raddr4 ? regfile_107 : _GEN_1002; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1004 = 7'h6c == io_i_raddr4 ? regfile_108 : _GEN_1003; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1005 = 7'h6d == io_i_raddr4 ? regfile_109 : _GEN_1004; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1006 = 7'h6e == io_i_raddr4 ? regfile_110 : _GEN_1005; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1007 = 7'h6f == io_i_raddr4 ? regfile_111 : _GEN_1006; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1008 = 7'h70 == io_i_raddr4 ? regfile_112 : _GEN_1007; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1009 = 7'h71 == io_i_raddr4 ? regfile_113 : _GEN_1008; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1010 = 7'h72 == io_i_raddr4 ? regfile_114 : _GEN_1009; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1011 = 7'h73 == io_i_raddr4 ? regfile_115 : _GEN_1010; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1012 = 7'h74 == io_i_raddr4 ? regfile_116 : _GEN_1011; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1013 = 7'h75 == io_i_raddr4 ? regfile_117 : _GEN_1012; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1014 = 7'h76 == io_i_raddr4 ? regfile_118 : _GEN_1013; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1015 = 7'h77 == io_i_raddr4 ? regfile_119 : _GEN_1014; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1016 = 7'h78 == io_i_raddr4 ? regfile_120 : _GEN_1015; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1017 = 7'h79 == io_i_raddr4 ? regfile_121 : _GEN_1016; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1018 = 7'h7a == io_i_raddr4 ? regfile_122 : _GEN_1017; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1019 = 7'h7b == io_i_raddr4 ? regfile_123 : _GEN_1018; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1020 = 7'h7c == io_i_raddr4 ? regfile_124 : _GEN_1019; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1021 = 7'h7d == io_i_raddr4 ? regfile_125 : _GEN_1020; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1022 = 7'h7e == io_i_raddr4 ? regfile_126 : _GEN_1021; // @[Mux.scala 101:{16,16}]
  wire [63:0] _GEN_1023 = 7'h7f == io_i_raddr4 ? regfile_127 : _GEN_1022; // @[Mux.scala 101:{16,16}]
  wire [63:0] _io_o_rdata4_T_4 = _io_o_rdata4_T_3 ? io_i_wdata2 : _GEN_1023; // @[Mux.scala 101:16]
  wire [63:0] debug_regs_0 = regfile_0; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_1 = regfile_1; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_2 = regfile_2; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_3 = regfile_3; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_4 = regfile_4; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_5 = regfile_5; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_6 = regfile_6; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_7 = regfile_7; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_8 = regfile_8; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_9 = regfile_9; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_10 = regfile_10; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_11 = regfile_11; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_12 = regfile_12; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_13 = regfile_13; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_14 = regfile_14; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_15 = regfile_15; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_16 = regfile_16; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_17 = regfile_17; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_18 = regfile_18; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_19 = regfile_19; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_20 = regfile_20; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_21 = regfile_21; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_22 = regfile_22; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_23 = regfile_23; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_24 = regfile_24; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_25 = regfile_25; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_26 = regfile_26; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_27 = regfile_27; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_28 = regfile_28; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_29 = regfile_29; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_30 = regfile_30; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_31 = regfile_31; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_32 = regfile_32; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_33 = regfile_33; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_34 = regfile_34; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_35 = regfile_35; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_36 = regfile_36; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_37 = regfile_37; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_38 = regfile_38; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_39 = regfile_39; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_40 = regfile_40; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_41 = regfile_41; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_42 = regfile_42; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_43 = regfile_43; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_44 = regfile_44; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_45 = regfile_45; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_46 = regfile_46; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_47 = regfile_47; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_48 = regfile_48; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_49 = regfile_49; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_50 = regfile_50; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_51 = regfile_51; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_52 = regfile_52; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_53 = regfile_53; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_54 = regfile_54; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_55 = regfile_55; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_56 = regfile_56; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_57 = regfile_57; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_58 = regfile_58; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_59 = regfile_59; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_60 = regfile_60; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_61 = regfile_61; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_62 = regfile_62; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_63 = regfile_63; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_64 = regfile_64; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_65 = regfile_65; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_66 = regfile_66; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_67 = regfile_67; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_68 = regfile_68; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_69 = regfile_69; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_70 = regfile_70; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_71 = regfile_71; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_72 = regfile_72; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_73 = regfile_73; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_74 = regfile_74; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_75 = regfile_75; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_76 = regfile_76; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_77 = regfile_77; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_78 = regfile_78; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_79 = regfile_79; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_80 = regfile_80; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_81 = regfile_81; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_82 = regfile_82; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_83 = regfile_83; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_84 = regfile_84; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_85 = regfile_85; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_86 = regfile_86; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_87 = regfile_87; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_88 = regfile_88; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_89 = regfile_89; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_90 = regfile_90; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_91 = regfile_91; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_92 = regfile_92; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_93 = regfile_93; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_94 = regfile_94; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_95 = regfile_95; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_96 = regfile_96; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_97 = regfile_97; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_98 = regfile_98; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_99 = regfile_99; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_100 = regfile_100; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_101 = regfile_101; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_102 = regfile_102; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_103 = regfile_103; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_104 = regfile_104; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_105 = regfile_105; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_106 = regfile_106; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_107 = regfile_107; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_108 = regfile_108; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_109 = regfile_109; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_110 = regfile_110; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_111 = regfile_111; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_112 = regfile_112; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_113 = regfile_113; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_114 = regfile_114; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_115 = regfile_115; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_116 = regfile_116; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_117 = regfile_117; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_118 = regfile_118; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_119 = regfile_119; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_120 = regfile_120; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_121 = regfile_121; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_122 = regfile_122; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_123 = regfile_123; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_124 = regfile_124; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_125 = regfile_125; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_126 = regfile_126; // @[regfile.scala 37:24 39:14]
  wire [63:0] debug_regs_127 = regfile_127; // @[regfile.scala 37:24 39:14]
  assign io_o_rdata1 = _io_o_rdata1_T_1 ? io_i_wdata1 : _io_o_rdata1_T_4; // @[Mux.scala 101:16]
  assign io_o_rdata2 = _io_o_rdata2_T_1 ? io_i_wdata1 : _io_o_rdata2_T_4; // @[Mux.scala 101:16]
  assign io_o_rdata3 = _io_o_rdata3_T_1 ? io_i_wdata1 : _io_o_rdata3_T_4; // @[Mux.scala 101:16]
  assign io_o_rdata4 = _io_o_rdata4_T_1 ? io_i_wdata1 : _io_o_rdata4_T_4; // @[Mux.scala 101:16]
  assign io_o_pregs_0 = regfile_0; // @[regfile.scala 41:14]
  assign io_o_pregs_1 = regfile_1; // @[regfile.scala 41:14]
  assign io_o_pregs_2 = regfile_2; // @[regfile.scala 41:14]
  assign io_o_pregs_3 = regfile_3; // @[regfile.scala 41:14]
  assign io_o_pregs_4 = regfile_4; // @[regfile.scala 41:14]
  assign io_o_pregs_5 = regfile_5; // @[regfile.scala 41:14]
  assign io_o_pregs_6 = regfile_6; // @[regfile.scala 41:14]
  assign io_o_pregs_7 = regfile_7; // @[regfile.scala 41:14]
  assign io_o_pregs_8 = regfile_8; // @[regfile.scala 41:14]
  assign io_o_pregs_9 = regfile_9; // @[regfile.scala 41:14]
  assign io_o_pregs_10 = regfile_10; // @[regfile.scala 41:14]
  assign io_o_pregs_11 = regfile_11; // @[regfile.scala 41:14]
  assign io_o_pregs_12 = regfile_12; // @[regfile.scala 41:14]
  assign io_o_pregs_13 = regfile_13; // @[regfile.scala 41:14]
  assign io_o_pregs_14 = regfile_14; // @[regfile.scala 41:14]
  assign io_o_pregs_15 = regfile_15; // @[regfile.scala 41:14]
  assign io_o_pregs_16 = regfile_16; // @[regfile.scala 41:14]
  assign io_o_pregs_17 = regfile_17; // @[regfile.scala 41:14]
  assign io_o_pregs_18 = regfile_18; // @[regfile.scala 41:14]
  assign io_o_pregs_19 = regfile_19; // @[regfile.scala 41:14]
  assign io_o_pregs_20 = regfile_20; // @[regfile.scala 41:14]
  assign io_o_pregs_21 = regfile_21; // @[regfile.scala 41:14]
  assign io_o_pregs_22 = regfile_22; // @[regfile.scala 41:14]
  assign io_o_pregs_23 = regfile_23; // @[regfile.scala 41:14]
  assign io_o_pregs_24 = regfile_24; // @[regfile.scala 41:14]
  assign io_o_pregs_25 = regfile_25; // @[regfile.scala 41:14]
  assign io_o_pregs_26 = regfile_26; // @[regfile.scala 41:14]
  assign io_o_pregs_27 = regfile_27; // @[regfile.scala 41:14]
  assign io_o_pregs_28 = regfile_28; // @[regfile.scala 41:14]
  assign io_o_pregs_29 = regfile_29; // @[regfile.scala 41:14]
  assign io_o_pregs_30 = regfile_30; // @[regfile.scala 41:14]
  assign io_o_pregs_31 = regfile_31; // @[regfile.scala 41:14]
  assign io_o_pregs_32 = regfile_32; // @[regfile.scala 41:14]
  assign io_o_pregs_33 = regfile_33; // @[regfile.scala 41:14]
  assign io_o_pregs_34 = regfile_34; // @[regfile.scala 41:14]
  assign io_o_pregs_35 = regfile_35; // @[regfile.scala 41:14]
  assign io_o_pregs_36 = regfile_36; // @[regfile.scala 41:14]
  assign io_o_pregs_37 = regfile_37; // @[regfile.scala 41:14]
  assign io_o_pregs_38 = regfile_38; // @[regfile.scala 41:14]
  assign io_o_pregs_39 = regfile_39; // @[regfile.scala 41:14]
  assign io_o_pregs_40 = regfile_40; // @[regfile.scala 41:14]
  assign io_o_pregs_41 = regfile_41; // @[regfile.scala 41:14]
  assign io_o_pregs_42 = regfile_42; // @[regfile.scala 41:14]
  assign io_o_pregs_43 = regfile_43; // @[regfile.scala 41:14]
  assign io_o_pregs_44 = regfile_44; // @[regfile.scala 41:14]
  assign io_o_pregs_45 = regfile_45; // @[regfile.scala 41:14]
  assign io_o_pregs_46 = regfile_46; // @[regfile.scala 41:14]
  assign io_o_pregs_47 = regfile_47; // @[regfile.scala 41:14]
  assign io_o_pregs_48 = regfile_48; // @[regfile.scala 41:14]
  assign io_o_pregs_49 = regfile_49; // @[regfile.scala 41:14]
  assign io_o_pregs_50 = regfile_50; // @[regfile.scala 41:14]
  assign io_o_pregs_51 = regfile_51; // @[regfile.scala 41:14]
  assign io_o_pregs_52 = regfile_52; // @[regfile.scala 41:14]
  assign io_o_pregs_53 = regfile_53; // @[regfile.scala 41:14]
  assign io_o_pregs_54 = regfile_54; // @[regfile.scala 41:14]
  assign io_o_pregs_55 = regfile_55; // @[regfile.scala 41:14]
  assign io_o_pregs_56 = regfile_56; // @[regfile.scala 41:14]
  assign io_o_pregs_57 = regfile_57; // @[regfile.scala 41:14]
  assign io_o_pregs_58 = regfile_58; // @[regfile.scala 41:14]
  assign io_o_pregs_59 = regfile_59; // @[regfile.scala 41:14]
  assign io_o_pregs_60 = regfile_60; // @[regfile.scala 41:14]
  assign io_o_pregs_61 = regfile_61; // @[regfile.scala 41:14]
  assign io_o_pregs_62 = regfile_62; // @[regfile.scala 41:14]
  assign io_o_pregs_63 = regfile_63; // @[regfile.scala 41:14]
  assign io_o_pregs_64 = regfile_64; // @[regfile.scala 41:14]
  assign io_o_pregs_65 = regfile_65; // @[regfile.scala 41:14]
  assign io_o_pregs_66 = regfile_66; // @[regfile.scala 41:14]
  assign io_o_pregs_67 = regfile_67; // @[regfile.scala 41:14]
  assign io_o_pregs_68 = regfile_68; // @[regfile.scala 41:14]
  assign io_o_pregs_69 = regfile_69; // @[regfile.scala 41:14]
  assign io_o_pregs_70 = regfile_70; // @[regfile.scala 41:14]
  assign io_o_pregs_71 = regfile_71; // @[regfile.scala 41:14]
  assign io_o_pregs_72 = regfile_72; // @[regfile.scala 41:14]
  assign io_o_pregs_73 = regfile_73; // @[regfile.scala 41:14]
  assign io_o_pregs_74 = regfile_74; // @[regfile.scala 41:14]
  assign io_o_pregs_75 = regfile_75; // @[regfile.scala 41:14]
  assign io_o_pregs_76 = regfile_76; // @[regfile.scala 41:14]
  assign io_o_pregs_77 = regfile_77; // @[regfile.scala 41:14]
  assign io_o_pregs_78 = regfile_78; // @[regfile.scala 41:14]
  assign io_o_pregs_79 = regfile_79; // @[regfile.scala 41:14]
  assign io_o_pregs_80 = regfile_80; // @[regfile.scala 41:14]
  assign io_o_pregs_81 = regfile_81; // @[regfile.scala 41:14]
  assign io_o_pregs_82 = regfile_82; // @[regfile.scala 41:14]
  assign io_o_pregs_83 = regfile_83; // @[regfile.scala 41:14]
  assign io_o_pregs_84 = regfile_84; // @[regfile.scala 41:14]
  assign io_o_pregs_85 = regfile_85; // @[regfile.scala 41:14]
  assign io_o_pregs_86 = regfile_86; // @[regfile.scala 41:14]
  assign io_o_pregs_87 = regfile_87; // @[regfile.scala 41:14]
  assign io_o_pregs_88 = regfile_88; // @[regfile.scala 41:14]
  assign io_o_pregs_89 = regfile_89; // @[regfile.scala 41:14]
  assign io_o_pregs_90 = regfile_90; // @[regfile.scala 41:14]
  assign io_o_pregs_91 = regfile_91; // @[regfile.scala 41:14]
  assign io_o_pregs_92 = regfile_92; // @[regfile.scala 41:14]
  assign io_o_pregs_93 = regfile_93; // @[regfile.scala 41:14]
  assign io_o_pregs_94 = regfile_94; // @[regfile.scala 41:14]
  assign io_o_pregs_95 = regfile_95; // @[regfile.scala 41:14]
  assign io_o_pregs_96 = regfile_96; // @[regfile.scala 41:14]
  assign io_o_pregs_97 = regfile_97; // @[regfile.scala 41:14]
  assign io_o_pregs_98 = regfile_98; // @[regfile.scala 41:14]
  assign io_o_pregs_99 = regfile_99; // @[regfile.scala 41:14]
  assign io_o_pregs_100 = regfile_100; // @[regfile.scala 41:14]
  assign io_o_pregs_101 = regfile_101; // @[regfile.scala 41:14]
  assign io_o_pregs_102 = regfile_102; // @[regfile.scala 41:14]
  assign io_o_pregs_103 = regfile_103; // @[regfile.scala 41:14]
  assign io_o_pregs_104 = regfile_104; // @[regfile.scala 41:14]
  assign io_o_pregs_105 = regfile_105; // @[regfile.scala 41:14]
  assign io_o_pregs_106 = regfile_106; // @[regfile.scala 41:14]
  assign io_o_pregs_107 = regfile_107; // @[regfile.scala 41:14]
  assign io_o_pregs_108 = regfile_108; // @[regfile.scala 41:14]
  assign io_o_pregs_109 = regfile_109; // @[regfile.scala 41:14]
  assign io_o_pregs_110 = regfile_110; // @[regfile.scala 41:14]
  assign io_o_pregs_111 = regfile_111; // @[regfile.scala 41:14]
  assign io_o_pregs_112 = regfile_112; // @[regfile.scala 41:14]
  assign io_o_pregs_113 = regfile_113; // @[regfile.scala 41:14]
  assign io_o_pregs_114 = regfile_114; // @[regfile.scala 41:14]
  assign io_o_pregs_115 = regfile_115; // @[regfile.scala 41:14]
  assign io_o_pregs_116 = regfile_116; // @[regfile.scala 41:14]
  assign io_o_pregs_117 = regfile_117; // @[regfile.scala 41:14]
  assign io_o_pregs_118 = regfile_118; // @[regfile.scala 41:14]
  assign io_o_pregs_119 = regfile_119; // @[regfile.scala 41:14]
  assign io_o_pregs_120 = regfile_120; // @[regfile.scala 41:14]
  assign io_o_pregs_121 = regfile_121; // @[regfile.scala 41:14]
  assign io_o_pregs_122 = regfile_122; // @[regfile.scala 41:14]
  assign io_o_pregs_123 = regfile_123; // @[regfile.scala 41:14]
  assign io_o_pregs_124 = regfile_124; // @[regfile.scala 41:14]
  assign io_o_pregs_125 = regfile_125; // @[regfile.scala 41:14]
  assign io_o_pregs_126 = regfile_126; // @[regfile.scala 41:14]
  assign io_o_pregs_127 = regfile_127; // @[regfile.scala 41:14]
  always @(posedge clock) begin
    if (reset) begin // @[regfile.scala 36:24]
      regfile_0 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h0 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_0 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_0 <= _GEN_128;
      end
    end else begin
      regfile_0 <= _GEN_128;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_1 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_1 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_1 <= _GEN_129;
      end
    end else begin
      regfile_1 <= _GEN_129;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_2 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_2 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_2 <= _GEN_130;
      end
    end else begin
      regfile_2 <= _GEN_130;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_3 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_3 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_3 <= _GEN_131;
      end
    end else begin
      regfile_3 <= _GEN_131;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_4 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_4 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_4 <= _GEN_132;
      end
    end else begin
      regfile_4 <= _GEN_132;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_5 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_5 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_5 <= _GEN_133;
      end
    end else begin
      regfile_5 <= _GEN_133;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_6 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_6 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_6 <= _GEN_134;
      end
    end else begin
      regfile_6 <= _GEN_134;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_7 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_7 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_7 <= _GEN_135;
      end
    end else begin
      regfile_7 <= _GEN_135;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_8 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h8 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_8 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_8 <= _GEN_136;
      end
    end else begin
      regfile_8 <= _GEN_136;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_9 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h9 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_9 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_9 <= _GEN_137;
      end
    end else begin
      regfile_9 <= _GEN_137;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_10 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'ha == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_10 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_10 <= _GEN_138;
      end
    end else begin
      regfile_10 <= _GEN_138;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_11 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'hb == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_11 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_11 <= _GEN_139;
      end
    end else begin
      regfile_11 <= _GEN_139;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_12 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'hc == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_12 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_12 <= _GEN_140;
      end
    end else begin
      regfile_12 <= _GEN_140;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_13 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'hd == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_13 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_13 <= _GEN_141;
      end
    end else begin
      regfile_13 <= _GEN_141;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_14 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'he == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_14 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_14 <= _GEN_142;
      end
    end else begin
      regfile_14 <= _GEN_142;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_15 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'hf == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_15 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_15 <= _GEN_143;
      end
    end else begin
      regfile_15 <= _GEN_143;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_16 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h10 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_16 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_16 <= _GEN_144;
      end
    end else begin
      regfile_16 <= _GEN_144;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_17 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h11 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_17 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_17 <= _GEN_145;
      end
    end else begin
      regfile_17 <= _GEN_145;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_18 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h12 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_18 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_18 <= _GEN_146;
      end
    end else begin
      regfile_18 <= _GEN_146;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_19 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h13 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_19 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_19 <= _GEN_147;
      end
    end else begin
      regfile_19 <= _GEN_147;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_20 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h14 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_20 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_20 <= _GEN_148;
      end
    end else begin
      regfile_20 <= _GEN_148;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_21 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h15 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_21 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_21 <= _GEN_149;
      end
    end else begin
      regfile_21 <= _GEN_149;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_22 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h16 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_22 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_22 <= _GEN_150;
      end
    end else begin
      regfile_22 <= _GEN_150;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_23 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h17 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_23 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_23 <= _GEN_151;
      end
    end else begin
      regfile_23 <= _GEN_151;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_24 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h18 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_24 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_24 <= _GEN_152;
      end
    end else begin
      regfile_24 <= _GEN_152;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_25 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h19 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_25 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_25 <= _GEN_153;
      end
    end else begin
      regfile_25 <= _GEN_153;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_26 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_26 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_26 <= _GEN_154;
      end
    end else begin
      regfile_26 <= _GEN_154;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_27 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_27 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_27 <= _GEN_155;
      end
    end else begin
      regfile_27 <= _GEN_155;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_28 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_28 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_28 <= _GEN_156;
      end
    end else begin
      regfile_28 <= _GEN_156;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_29 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_29 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_29 <= _GEN_157;
      end
    end else begin
      regfile_29 <= _GEN_157;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_30 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_30 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_30 <= _GEN_158;
      end
    end else begin
      regfile_30 <= _GEN_158;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_31 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h1f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_31 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_31 <= _GEN_159;
      end
    end else begin
      regfile_31 <= _GEN_159;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_32 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h20 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_32 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_32 <= _GEN_160;
      end
    end else begin
      regfile_32 <= _GEN_160;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_33 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h21 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_33 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_33 <= _GEN_161;
      end
    end else begin
      regfile_33 <= _GEN_161;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_34 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h22 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_34 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_34 <= _GEN_162;
      end
    end else begin
      regfile_34 <= _GEN_162;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_35 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h23 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_35 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_35 <= _GEN_163;
      end
    end else begin
      regfile_35 <= _GEN_163;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_36 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h24 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_36 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_36 <= _GEN_164;
      end
    end else begin
      regfile_36 <= _GEN_164;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_37 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h25 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_37 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_37 <= _GEN_165;
      end
    end else begin
      regfile_37 <= _GEN_165;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_38 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h26 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_38 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_38 <= _GEN_166;
      end
    end else begin
      regfile_38 <= _GEN_166;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_39 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h27 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_39 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_39 <= _GEN_167;
      end
    end else begin
      regfile_39 <= _GEN_167;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_40 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h28 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_40 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_40 <= _GEN_168;
      end
    end else begin
      regfile_40 <= _GEN_168;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_41 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h29 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_41 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_41 <= _GEN_169;
      end
    end else begin
      regfile_41 <= _GEN_169;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_42 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_42 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_42 <= _GEN_170;
      end
    end else begin
      regfile_42 <= _GEN_170;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_43 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_43 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_43 <= _GEN_171;
      end
    end else begin
      regfile_43 <= _GEN_171;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_44 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_44 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_44 <= _GEN_172;
      end
    end else begin
      regfile_44 <= _GEN_172;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_45 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_45 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_45 <= _GEN_173;
      end
    end else begin
      regfile_45 <= _GEN_173;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_46 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_46 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_46 <= _GEN_174;
      end
    end else begin
      regfile_46 <= _GEN_174;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_47 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h2f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_47 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_47 <= _GEN_175;
      end
    end else begin
      regfile_47 <= _GEN_175;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_48 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h30 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_48 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_48 <= _GEN_176;
      end
    end else begin
      regfile_48 <= _GEN_176;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_49 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h31 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_49 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_49 <= _GEN_177;
      end
    end else begin
      regfile_49 <= _GEN_177;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_50 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h32 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_50 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_50 <= _GEN_178;
      end
    end else begin
      regfile_50 <= _GEN_178;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_51 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h33 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_51 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_51 <= _GEN_179;
      end
    end else begin
      regfile_51 <= _GEN_179;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_52 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h34 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_52 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_52 <= _GEN_180;
      end
    end else begin
      regfile_52 <= _GEN_180;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_53 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h35 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_53 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_53 <= _GEN_181;
      end
    end else begin
      regfile_53 <= _GEN_181;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_54 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h36 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_54 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_54 <= _GEN_182;
      end
    end else begin
      regfile_54 <= _GEN_182;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_55 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h37 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_55 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_55 <= _GEN_183;
      end
    end else begin
      regfile_55 <= _GEN_183;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_56 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h38 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_56 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_56 <= _GEN_184;
      end
    end else begin
      regfile_56 <= _GEN_184;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_57 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h39 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_57 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_57 <= _GEN_185;
      end
    end else begin
      regfile_57 <= _GEN_185;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_58 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_58 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_58 <= _GEN_186;
      end
    end else begin
      regfile_58 <= _GEN_186;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_59 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_59 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_59 <= _GEN_187;
      end
    end else begin
      regfile_59 <= _GEN_187;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_60 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_60 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_60 <= _GEN_188;
      end
    end else begin
      regfile_60 <= _GEN_188;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_61 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_61 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_61 <= _GEN_189;
      end
    end else begin
      regfile_61 <= _GEN_189;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_62 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_62 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_62 <= _GEN_190;
      end
    end else begin
      regfile_62 <= _GEN_190;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_63 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h3f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_63 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_63 <= _GEN_191;
      end
    end else begin
      regfile_63 <= _GEN_191;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_64 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h40 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_64 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_64 <= _GEN_192;
      end
    end else begin
      regfile_64 <= _GEN_192;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_65 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h41 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_65 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_65 <= _GEN_193;
      end
    end else begin
      regfile_65 <= _GEN_193;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_66 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h42 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_66 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_66 <= _GEN_194;
      end
    end else begin
      regfile_66 <= _GEN_194;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_67 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h43 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_67 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_67 <= _GEN_195;
      end
    end else begin
      regfile_67 <= _GEN_195;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_68 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h44 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_68 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_68 <= _GEN_196;
      end
    end else begin
      regfile_68 <= _GEN_196;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_69 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h45 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_69 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_69 <= _GEN_197;
      end
    end else begin
      regfile_69 <= _GEN_197;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_70 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h46 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_70 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_70 <= _GEN_198;
      end
    end else begin
      regfile_70 <= _GEN_198;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_71 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h47 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_71 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_71 <= _GEN_199;
      end
    end else begin
      regfile_71 <= _GEN_199;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_72 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h48 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_72 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_72 <= _GEN_200;
      end
    end else begin
      regfile_72 <= _GEN_200;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_73 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h49 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_73 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_73 <= _GEN_201;
      end
    end else begin
      regfile_73 <= _GEN_201;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_74 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_74 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_74 <= _GEN_202;
      end
    end else begin
      regfile_74 <= _GEN_202;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_75 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_75 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_75 <= _GEN_203;
      end
    end else begin
      regfile_75 <= _GEN_203;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_76 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_76 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_76 <= _GEN_204;
      end
    end else begin
      regfile_76 <= _GEN_204;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_77 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_77 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_77 <= _GEN_205;
      end
    end else begin
      regfile_77 <= _GEN_205;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_78 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_78 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_78 <= _GEN_206;
      end
    end else begin
      regfile_78 <= _GEN_206;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_79 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h4f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_79 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_79 <= _GEN_207;
      end
    end else begin
      regfile_79 <= _GEN_207;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_80 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h50 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_80 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_80 <= _GEN_208;
      end
    end else begin
      regfile_80 <= _GEN_208;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_81 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h51 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_81 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_81 <= _GEN_209;
      end
    end else begin
      regfile_81 <= _GEN_209;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_82 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h52 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_82 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_82 <= _GEN_210;
      end
    end else begin
      regfile_82 <= _GEN_210;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_83 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h53 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_83 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_83 <= _GEN_211;
      end
    end else begin
      regfile_83 <= _GEN_211;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_84 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h54 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_84 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_84 <= _GEN_212;
      end
    end else begin
      regfile_84 <= _GEN_212;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_85 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h55 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_85 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_85 <= _GEN_213;
      end
    end else begin
      regfile_85 <= _GEN_213;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_86 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h56 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_86 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_86 <= _GEN_214;
      end
    end else begin
      regfile_86 <= _GEN_214;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_87 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h57 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_87 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_87 <= _GEN_215;
      end
    end else begin
      regfile_87 <= _GEN_215;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_88 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h58 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_88 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_88 <= _GEN_216;
      end
    end else begin
      regfile_88 <= _GEN_216;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_89 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h59 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_89 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_89 <= _GEN_217;
      end
    end else begin
      regfile_89 <= _GEN_217;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_90 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_90 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_90 <= _GEN_218;
      end
    end else begin
      regfile_90 <= _GEN_218;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_91 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_91 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_91 <= _GEN_219;
      end
    end else begin
      regfile_91 <= _GEN_219;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_92 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_92 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_92 <= _GEN_220;
      end
    end else begin
      regfile_92 <= _GEN_220;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_93 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_93 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_93 <= _GEN_221;
      end
    end else begin
      regfile_93 <= _GEN_221;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_94 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_94 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_94 <= _GEN_222;
      end
    end else begin
      regfile_94 <= _GEN_222;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_95 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h5f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_95 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_95 <= _GEN_223;
      end
    end else begin
      regfile_95 <= _GEN_223;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_96 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h60 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_96 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_96 <= _GEN_224;
      end
    end else begin
      regfile_96 <= _GEN_224;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_97 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h61 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_97 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_97 <= _GEN_225;
      end
    end else begin
      regfile_97 <= _GEN_225;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_98 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h62 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_98 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_98 <= _GEN_226;
      end
    end else begin
      regfile_98 <= _GEN_226;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_99 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h63 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_99 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_99 <= _GEN_227;
      end
    end else begin
      regfile_99 <= _GEN_227;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_100 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h64 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_100 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_100 <= _GEN_228;
      end
    end else begin
      regfile_100 <= _GEN_228;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_101 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h65 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_101 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_101 <= _GEN_229;
      end
    end else begin
      regfile_101 <= _GEN_229;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_102 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h66 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_102 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_102 <= _GEN_230;
      end
    end else begin
      regfile_102 <= _GEN_230;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_103 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h67 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_103 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_103 <= _GEN_231;
      end
    end else begin
      regfile_103 <= _GEN_231;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_104 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h68 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_104 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_104 <= _GEN_232;
      end
    end else begin
      regfile_104 <= _GEN_232;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_105 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h69 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_105 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_105 <= _GEN_233;
      end
    end else begin
      regfile_105 <= _GEN_233;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_106 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_106 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_106 <= _GEN_234;
      end
    end else begin
      regfile_106 <= _GEN_234;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_107 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_107 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_107 <= _GEN_235;
      end
    end else begin
      regfile_107 <= _GEN_235;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_108 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_108 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_108 <= _GEN_236;
      end
    end else begin
      regfile_108 <= _GEN_236;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_109 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_109 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_109 <= _GEN_237;
      end
    end else begin
      regfile_109 <= _GEN_237;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_110 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_110 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_110 <= _GEN_238;
      end
    end else begin
      regfile_110 <= _GEN_238;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_111 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h6f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_111 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_111 <= _GEN_239;
      end
    end else begin
      regfile_111 <= _GEN_239;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_112 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h70 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_112 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_112 <= _GEN_240;
      end
    end else begin
      regfile_112 <= _GEN_240;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_113 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h71 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_113 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_113 <= _GEN_241;
      end
    end else begin
      regfile_113 <= _GEN_241;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_114 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h72 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_114 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_114 <= _GEN_242;
      end
    end else begin
      regfile_114 <= _GEN_242;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_115 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h73 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_115 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_115 <= _GEN_243;
      end
    end else begin
      regfile_115 <= _GEN_243;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_116 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h74 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_116 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_116 <= _GEN_244;
      end
    end else begin
      regfile_116 <= _GEN_244;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_117 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h75 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_117 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_117 <= _GEN_245;
      end
    end else begin
      regfile_117 <= _GEN_245;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_118 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h76 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_118 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_118 <= _GEN_246;
      end
    end else begin
      regfile_118 <= _GEN_246;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_119 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h77 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_119 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_119 <= _GEN_247;
      end
    end else begin
      regfile_119 <= _GEN_247;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_120 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h78 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_120 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_120 <= _GEN_248;
      end
    end else begin
      regfile_120 <= _GEN_248;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_121 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h79 == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_121 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_121 <= _GEN_249;
      end
    end else begin
      regfile_121 <= _GEN_249;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_122 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7a == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_122 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_122 <= _GEN_250;
      end
    end else begin
      regfile_122 <= _GEN_250;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_123 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7b == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_123 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_123 <= _GEN_251;
      end
    end else begin
      regfile_123 <= _GEN_251;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_124 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7c == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_124 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_124 <= _GEN_252;
      end
    end else begin
      regfile_124 <= _GEN_252;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_125 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7d == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_125 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_125 <= _GEN_253;
      end
    end else begin
      regfile_125 <= _GEN_253;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_126 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7e == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_126 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_126 <= _GEN_254;
      end
    end else begin
      regfile_126 <= _GEN_254;
    end
    if (reset) begin // @[regfile.scala 36:24]
      regfile_127 <= 64'h0; // @[regfile.scala 36:24]
    end else if (io_i_wenable2) begin // @[regfile.scala 47:23]
      if (7'h7f == io_i_waddr2) begin // @[regfile.scala 48:26]
        regfile_127 <= io_i_wdata2; // @[regfile.scala 48:26]
      end else begin
        regfile_127 <= _GEN_255;
      end
    end else begin
      regfile_127 <= _GEN_255;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regfile_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regfile_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regfile_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regfile_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regfile_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regfile_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regfile_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regfile_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regfile_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regfile_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regfile_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regfile_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regfile_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regfile_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regfile_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regfile_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regfile_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regfile_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regfile_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regfile_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regfile_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regfile_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regfile_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regfile_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regfile_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regfile_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regfile_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regfile_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regfile_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regfile_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regfile_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regfile_31 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  regfile_32 = _RAND_32[63:0];
  _RAND_33 = {2{`RANDOM}};
  regfile_33 = _RAND_33[63:0];
  _RAND_34 = {2{`RANDOM}};
  regfile_34 = _RAND_34[63:0];
  _RAND_35 = {2{`RANDOM}};
  regfile_35 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  regfile_36 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  regfile_37 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  regfile_38 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  regfile_39 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  regfile_40 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  regfile_41 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  regfile_42 = _RAND_42[63:0];
  _RAND_43 = {2{`RANDOM}};
  regfile_43 = _RAND_43[63:0];
  _RAND_44 = {2{`RANDOM}};
  regfile_44 = _RAND_44[63:0];
  _RAND_45 = {2{`RANDOM}};
  regfile_45 = _RAND_45[63:0];
  _RAND_46 = {2{`RANDOM}};
  regfile_46 = _RAND_46[63:0];
  _RAND_47 = {2{`RANDOM}};
  regfile_47 = _RAND_47[63:0];
  _RAND_48 = {2{`RANDOM}};
  regfile_48 = _RAND_48[63:0];
  _RAND_49 = {2{`RANDOM}};
  regfile_49 = _RAND_49[63:0];
  _RAND_50 = {2{`RANDOM}};
  regfile_50 = _RAND_50[63:0];
  _RAND_51 = {2{`RANDOM}};
  regfile_51 = _RAND_51[63:0];
  _RAND_52 = {2{`RANDOM}};
  regfile_52 = _RAND_52[63:0];
  _RAND_53 = {2{`RANDOM}};
  regfile_53 = _RAND_53[63:0];
  _RAND_54 = {2{`RANDOM}};
  regfile_54 = _RAND_54[63:0];
  _RAND_55 = {2{`RANDOM}};
  regfile_55 = _RAND_55[63:0];
  _RAND_56 = {2{`RANDOM}};
  regfile_56 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  regfile_57 = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  regfile_58 = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  regfile_59 = _RAND_59[63:0];
  _RAND_60 = {2{`RANDOM}};
  regfile_60 = _RAND_60[63:0];
  _RAND_61 = {2{`RANDOM}};
  regfile_61 = _RAND_61[63:0];
  _RAND_62 = {2{`RANDOM}};
  regfile_62 = _RAND_62[63:0];
  _RAND_63 = {2{`RANDOM}};
  regfile_63 = _RAND_63[63:0];
  _RAND_64 = {2{`RANDOM}};
  regfile_64 = _RAND_64[63:0];
  _RAND_65 = {2{`RANDOM}};
  regfile_65 = _RAND_65[63:0];
  _RAND_66 = {2{`RANDOM}};
  regfile_66 = _RAND_66[63:0];
  _RAND_67 = {2{`RANDOM}};
  regfile_67 = _RAND_67[63:0];
  _RAND_68 = {2{`RANDOM}};
  regfile_68 = _RAND_68[63:0];
  _RAND_69 = {2{`RANDOM}};
  regfile_69 = _RAND_69[63:0];
  _RAND_70 = {2{`RANDOM}};
  regfile_70 = _RAND_70[63:0];
  _RAND_71 = {2{`RANDOM}};
  regfile_71 = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  regfile_72 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  regfile_73 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  regfile_74 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  regfile_75 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  regfile_76 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  regfile_77 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  regfile_78 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  regfile_79 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  regfile_80 = _RAND_80[63:0];
  _RAND_81 = {2{`RANDOM}};
  regfile_81 = _RAND_81[63:0];
  _RAND_82 = {2{`RANDOM}};
  regfile_82 = _RAND_82[63:0];
  _RAND_83 = {2{`RANDOM}};
  regfile_83 = _RAND_83[63:0];
  _RAND_84 = {2{`RANDOM}};
  regfile_84 = _RAND_84[63:0];
  _RAND_85 = {2{`RANDOM}};
  regfile_85 = _RAND_85[63:0];
  _RAND_86 = {2{`RANDOM}};
  regfile_86 = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  regfile_87 = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  regfile_88 = _RAND_88[63:0];
  _RAND_89 = {2{`RANDOM}};
  regfile_89 = _RAND_89[63:0];
  _RAND_90 = {2{`RANDOM}};
  regfile_90 = _RAND_90[63:0];
  _RAND_91 = {2{`RANDOM}};
  regfile_91 = _RAND_91[63:0];
  _RAND_92 = {2{`RANDOM}};
  regfile_92 = _RAND_92[63:0];
  _RAND_93 = {2{`RANDOM}};
  regfile_93 = _RAND_93[63:0];
  _RAND_94 = {2{`RANDOM}};
  regfile_94 = _RAND_94[63:0];
  _RAND_95 = {2{`RANDOM}};
  regfile_95 = _RAND_95[63:0];
  _RAND_96 = {2{`RANDOM}};
  regfile_96 = _RAND_96[63:0];
  _RAND_97 = {2{`RANDOM}};
  regfile_97 = _RAND_97[63:0];
  _RAND_98 = {2{`RANDOM}};
  regfile_98 = _RAND_98[63:0];
  _RAND_99 = {2{`RANDOM}};
  regfile_99 = _RAND_99[63:0];
  _RAND_100 = {2{`RANDOM}};
  regfile_100 = _RAND_100[63:0];
  _RAND_101 = {2{`RANDOM}};
  regfile_101 = _RAND_101[63:0];
  _RAND_102 = {2{`RANDOM}};
  regfile_102 = _RAND_102[63:0];
  _RAND_103 = {2{`RANDOM}};
  regfile_103 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  regfile_104 = _RAND_104[63:0];
  _RAND_105 = {2{`RANDOM}};
  regfile_105 = _RAND_105[63:0];
  _RAND_106 = {2{`RANDOM}};
  regfile_106 = _RAND_106[63:0];
  _RAND_107 = {2{`RANDOM}};
  regfile_107 = _RAND_107[63:0];
  _RAND_108 = {2{`RANDOM}};
  regfile_108 = _RAND_108[63:0];
  _RAND_109 = {2{`RANDOM}};
  regfile_109 = _RAND_109[63:0];
  _RAND_110 = {2{`RANDOM}};
  regfile_110 = _RAND_110[63:0];
  _RAND_111 = {2{`RANDOM}};
  regfile_111 = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  regfile_112 = _RAND_112[63:0];
  _RAND_113 = {2{`RANDOM}};
  regfile_113 = _RAND_113[63:0];
  _RAND_114 = {2{`RANDOM}};
  regfile_114 = _RAND_114[63:0];
  _RAND_115 = {2{`RANDOM}};
  regfile_115 = _RAND_115[63:0];
  _RAND_116 = {2{`RANDOM}};
  regfile_116 = _RAND_116[63:0];
  _RAND_117 = {2{`RANDOM}};
  regfile_117 = _RAND_117[63:0];
  _RAND_118 = {2{`RANDOM}};
  regfile_118 = _RAND_118[63:0];
  _RAND_119 = {2{`RANDOM}};
  regfile_119 = _RAND_119[63:0];
  _RAND_120 = {2{`RANDOM}};
  regfile_120 = _RAND_120[63:0];
  _RAND_121 = {2{`RANDOM}};
  regfile_121 = _RAND_121[63:0];
  _RAND_122 = {2{`RANDOM}};
  regfile_122 = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  regfile_123 = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  regfile_124 = _RAND_124[63:0];
  _RAND_125 = {2{`RANDOM}};
  regfile_125 = _RAND_125[63:0];
  _RAND_126 = {2{`RANDOM}};
  regfile_126 = _RAND_126[63:0];
  _RAND_127 = {2{`RANDOM}};
  regfile_127 = _RAND_127[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

module Dcache(
  input          clock,
  input          reset,
  output         io_cpu_mem_data_valid,
  output         io_cpu_mem_addr_ready,
  input          io_cpu_mem_Mwout,
  input  [63:0]  io_cpu_mem_Maddr,
  input          io_cpu_mem_Men,
  input  [31:0]  io_cpu_mem_Mlen,
  output [63:0]  io_cpu_mem_MdataIn,
  input  [63:0]  io_cpu_mem_MdataOut,
  output         io_mem_master_readAddr_valid,
  output [63:0]  io_mem_master_readAddr_bits_addr,
  output         io_mem_master_readData_ready,
  input          io_mem_master_readData_valid,
  input  [127:0] io_mem_master_readData_bits_data,
  input          io_mem_master_writeAddr_ready,
  output         io_mem_master_writeAddr_valid,
  output [63:0]  io_mem_master_writeAddr_bits_addr,
  input          io_mem_master_writeData_ready,
  output         io_mem_master_writeData_valid,
  output [127:0] io_mem_master_writeData_bits_data,
  output [15:0]  io_mem_master_writeData_bits_strb,
  output         io_mem_master_writeResp_ready,
  input          io_mem_master_writeResp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_256;
  reg [63:0] _RAND_257;
  reg [63:0] _RAND_258;
  reg [63:0] _RAND_259;
  reg [63:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [63:0] _RAND_263;
  reg [63:0] _RAND_264;
  reg [63:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [127:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
`endif // RANDOMIZE_REG_INIT
  wire  data_array_0_clock; // @[dcache.scala 52:36]
  wire  data_array_0_reset; // @[dcache.scala 52:36]
  wire  data_array_0_io_i_wen; // @[dcache.scala 52:36]
  wire [15:0] data_array_0_io_i_wstrb; // @[dcache.scala 52:36]
  wire [6:0] data_array_0_io_i_addr; // @[dcache.scala 52:36]
  wire [127:0] data_array_0_io_i_wdata; // @[dcache.scala 52:36]
  wire [127:0] data_array_0_io_o_rdata; // @[dcache.scala 52:36]
  wire  data_array_1_clock; // @[dcache.scala 52:36]
  wire  data_array_1_reset; // @[dcache.scala 52:36]
  wire  data_array_1_io_i_wen; // @[dcache.scala 52:36]
  wire [15:0] data_array_1_io_i_wstrb; // @[dcache.scala 52:36]
  wire [6:0] data_array_1_io_i_addr; // @[dcache.scala 52:36]
  wire [127:0] data_array_1_io_i_wdata; // @[dcache.scala 52:36]
  wire [127:0] data_array_1_io_o_rdata; // @[dcache.scala 52:36]
  wire [17:0] _VGA_MEM_BLK_E_T = 9'h190 * 9'h12c; // @[dcache.scala 30:56]
  wire [63:0] _GEN_3335 = {{46'd0}, _VGA_MEM_BLK_E_T}; // @[dcache.scala 30:47]
  wire [63:0] VGA_MEM_BLK_E = 64'ha1000000 + _GEN_3335; // @[dcache.scala 30:47]
  reg  cpu_mem_Mwout; // @[dcache.scala 35:22]
  reg [63:0] cpu_mem_Maddr; // @[dcache.scala 35:22]
  reg  cpu_mem_Men; // @[dcache.scala 35:22]
  reg [31:0] cpu_mem_Mlen; // @[dcache.scala 35:22]
  reg [63:0] cpu_mem_MdataOut; // @[dcache.scala 35:22]
  reg  last_req_Mwout; // @[dcache.scala 36:23]
  reg [63:0] last_req_Maddr; // @[dcache.scala 36:23]
  reg  last_req_Men; // @[dcache.scala 36:23]
  reg [31:0] last_req_Mlen; // @[dcache.scala 36:23]
  reg [63:0] last_req_MdataOut; // @[dcache.scala 36:23]
  wire  _new_req_T_5 = last_req_Mlen == cpu_mem_Mlen; // @[dcache.scala 39:19]
  wire  _new_req_T_6 = last_req_Mwout == cpu_mem_Mwout & last_req_Men == cpu_mem_Men & last_req_Maddr == cpu_mem_Maddr
     & _new_req_T_5; // @[dcache.scala 38:113]
  wire  _new_req_T_8 = _new_req_T_6 & last_req_MdataOut == cpu_mem_MdataOut; // @[dcache.scala 39:35]
  wire  new_req = ~_new_req_T_8; // @[dcache.scala 38:15]
  reg [52:0] tags0_0; // @[dcache.scala 46:20]
  reg [52:0] tags0_1; // @[dcache.scala 46:20]
  reg [52:0] tags0_2; // @[dcache.scala 46:20]
  reg [52:0] tags0_3; // @[dcache.scala 46:20]
  reg [52:0] tags0_4; // @[dcache.scala 46:20]
  reg [52:0] tags0_5; // @[dcache.scala 46:20]
  reg [52:0] tags0_6; // @[dcache.scala 46:20]
  reg [52:0] tags0_7; // @[dcache.scala 46:20]
  reg [52:0] tags0_8; // @[dcache.scala 46:20]
  reg [52:0] tags0_9; // @[dcache.scala 46:20]
  reg [52:0] tags0_10; // @[dcache.scala 46:20]
  reg [52:0] tags0_11; // @[dcache.scala 46:20]
  reg [52:0] tags0_12; // @[dcache.scala 46:20]
  reg [52:0] tags0_13; // @[dcache.scala 46:20]
  reg [52:0] tags0_14; // @[dcache.scala 46:20]
  reg [52:0] tags0_15; // @[dcache.scala 46:20]
  reg [52:0] tags0_16; // @[dcache.scala 46:20]
  reg [52:0] tags0_17; // @[dcache.scala 46:20]
  reg [52:0] tags0_18; // @[dcache.scala 46:20]
  reg [52:0] tags0_19; // @[dcache.scala 46:20]
  reg [52:0] tags0_20; // @[dcache.scala 46:20]
  reg [52:0] tags0_21; // @[dcache.scala 46:20]
  reg [52:0] tags0_22; // @[dcache.scala 46:20]
  reg [52:0] tags0_23; // @[dcache.scala 46:20]
  reg [52:0] tags0_24; // @[dcache.scala 46:20]
  reg [52:0] tags0_25; // @[dcache.scala 46:20]
  reg [52:0] tags0_26; // @[dcache.scala 46:20]
  reg [52:0] tags0_27; // @[dcache.scala 46:20]
  reg [52:0] tags0_28; // @[dcache.scala 46:20]
  reg [52:0] tags0_29; // @[dcache.scala 46:20]
  reg [52:0] tags0_30; // @[dcache.scala 46:20]
  reg [52:0] tags0_31; // @[dcache.scala 46:20]
  reg [52:0] tags0_32; // @[dcache.scala 46:20]
  reg [52:0] tags0_33; // @[dcache.scala 46:20]
  reg [52:0] tags0_34; // @[dcache.scala 46:20]
  reg [52:0] tags0_35; // @[dcache.scala 46:20]
  reg [52:0] tags0_36; // @[dcache.scala 46:20]
  reg [52:0] tags0_37; // @[dcache.scala 46:20]
  reg [52:0] tags0_38; // @[dcache.scala 46:20]
  reg [52:0] tags0_39; // @[dcache.scala 46:20]
  reg [52:0] tags0_40; // @[dcache.scala 46:20]
  reg [52:0] tags0_41; // @[dcache.scala 46:20]
  reg [52:0] tags0_42; // @[dcache.scala 46:20]
  reg [52:0] tags0_43; // @[dcache.scala 46:20]
  reg [52:0] tags0_44; // @[dcache.scala 46:20]
  reg [52:0] tags0_45; // @[dcache.scala 46:20]
  reg [52:0] tags0_46; // @[dcache.scala 46:20]
  reg [52:0] tags0_47; // @[dcache.scala 46:20]
  reg [52:0] tags0_48; // @[dcache.scala 46:20]
  reg [52:0] tags0_49; // @[dcache.scala 46:20]
  reg [52:0] tags0_50; // @[dcache.scala 46:20]
  reg [52:0] tags0_51; // @[dcache.scala 46:20]
  reg [52:0] tags0_52; // @[dcache.scala 46:20]
  reg [52:0] tags0_53; // @[dcache.scala 46:20]
  reg [52:0] tags0_54; // @[dcache.scala 46:20]
  reg [52:0] tags0_55; // @[dcache.scala 46:20]
  reg [52:0] tags0_56; // @[dcache.scala 46:20]
  reg [52:0] tags0_57; // @[dcache.scala 46:20]
  reg [52:0] tags0_58; // @[dcache.scala 46:20]
  reg [52:0] tags0_59; // @[dcache.scala 46:20]
  reg [52:0] tags0_60; // @[dcache.scala 46:20]
  reg [52:0] tags0_61; // @[dcache.scala 46:20]
  reg [52:0] tags0_62; // @[dcache.scala 46:20]
  reg [52:0] tags0_63; // @[dcache.scala 46:20]
  reg [52:0] tags0_64; // @[dcache.scala 46:20]
  reg [52:0] tags0_65; // @[dcache.scala 46:20]
  reg [52:0] tags0_66; // @[dcache.scala 46:20]
  reg [52:0] tags0_67; // @[dcache.scala 46:20]
  reg [52:0] tags0_68; // @[dcache.scala 46:20]
  reg [52:0] tags0_69; // @[dcache.scala 46:20]
  reg [52:0] tags0_70; // @[dcache.scala 46:20]
  reg [52:0] tags0_71; // @[dcache.scala 46:20]
  reg [52:0] tags0_72; // @[dcache.scala 46:20]
  reg [52:0] tags0_73; // @[dcache.scala 46:20]
  reg [52:0] tags0_74; // @[dcache.scala 46:20]
  reg [52:0] tags0_75; // @[dcache.scala 46:20]
  reg [52:0] tags0_76; // @[dcache.scala 46:20]
  reg [52:0] tags0_77; // @[dcache.scala 46:20]
  reg [52:0] tags0_78; // @[dcache.scala 46:20]
  reg [52:0] tags0_79; // @[dcache.scala 46:20]
  reg [52:0] tags0_80; // @[dcache.scala 46:20]
  reg [52:0] tags0_81; // @[dcache.scala 46:20]
  reg [52:0] tags0_82; // @[dcache.scala 46:20]
  reg [52:0] tags0_83; // @[dcache.scala 46:20]
  reg [52:0] tags0_84; // @[dcache.scala 46:20]
  reg [52:0] tags0_85; // @[dcache.scala 46:20]
  reg [52:0] tags0_86; // @[dcache.scala 46:20]
  reg [52:0] tags0_87; // @[dcache.scala 46:20]
  reg [52:0] tags0_88; // @[dcache.scala 46:20]
  reg [52:0] tags0_89; // @[dcache.scala 46:20]
  reg [52:0] tags0_90; // @[dcache.scala 46:20]
  reg [52:0] tags0_91; // @[dcache.scala 46:20]
  reg [52:0] tags0_92; // @[dcache.scala 46:20]
  reg [52:0] tags0_93; // @[dcache.scala 46:20]
  reg [52:0] tags0_94; // @[dcache.scala 46:20]
  reg [52:0] tags0_95; // @[dcache.scala 46:20]
  reg [52:0] tags0_96; // @[dcache.scala 46:20]
  reg [52:0] tags0_97; // @[dcache.scala 46:20]
  reg [52:0] tags0_98; // @[dcache.scala 46:20]
  reg [52:0] tags0_99; // @[dcache.scala 46:20]
  reg [52:0] tags0_100; // @[dcache.scala 46:20]
  reg [52:0] tags0_101; // @[dcache.scala 46:20]
  reg [52:0] tags0_102; // @[dcache.scala 46:20]
  reg [52:0] tags0_103; // @[dcache.scala 46:20]
  reg [52:0] tags0_104; // @[dcache.scala 46:20]
  reg [52:0] tags0_105; // @[dcache.scala 46:20]
  reg [52:0] tags0_106; // @[dcache.scala 46:20]
  reg [52:0] tags0_107; // @[dcache.scala 46:20]
  reg [52:0] tags0_108; // @[dcache.scala 46:20]
  reg [52:0] tags0_109; // @[dcache.scala 46:20]
  reg [52:0] tags0_110; // @[dcache.scala 46:20]
  reg [52:0] tags0_111; // @[dcache.scala 46:20]
  reg [52:0] tags0_112; // @[dcache.scala 46:20]
  reg [52:0] tags0_113; // @[dcache.scala 46:20]
  reg [52:0] tags0_114; // @[dcache.scala 46:20]
  reg [52:0] tags0_115; // @[dcache.scala 46:20]
  reg [52:0] tags0_116; // @[dcache.scala 46:20]
  reg [52:0] tags0_117; // @[dcache.scala 46:20]
  reg [52:0] tags0_118; // @[dcache.scala 46:20]
  reg [52:0] tags0_119; // @[dcache.scala 46:20]
  reg [52:0] tags0_120; // @[dcache.scala 46:20]
  reg [52:0] tags0_121; // @[dcache.scala 46:20]
  reg [52:0] tags0_122; // @[dcache.scala 46:20]
  reg [52:0] tags0_123; // @[dcache.scala 46:20]
  reg [52:0] tags0_124; // @[dcache.scala 46:20]
  reg [52:0] tags0_125; // @[dcache.scala 46:20]
  reg [52:0] tags0_126; // @[dcache.scala 46:20]
  reg [52:0] tags0_127; // @[dcache.scala 46:20]
  reg [52:0] tags1_0; // @[dcache.scala 47:20]
  reg [52:0] tags1_1; // @[dcache.scala 47:20]
  reg [52:0] tags1_2; // @[dcache.scala 47:20]
  reg [52:0] tags1_3; // @[dcache.scala 47:20]
  reg [52:0] tags1_4; // @[dcache.scala 47:20]
  reg [52:0] tags1_5; // @[dcache.scala 47:20]
  reg [52:0] tags1_6; // @[dcache.scala 47:20]
  reg [52:0] tags1_7; // @[dcache.scala 47:20]
  reg [52:0] tags1_8; // @[dcache.scala 47:20]
  reg [52:0] tags1_9; // @[dcache.scala 47:20]
  reg [52:0] tags1_10; // @[dcache.scala 47:20]
  reg [52:0] tags1_11; // @[dcache.scala 47:20]
  reg [52:0] tags1_12; // @[dcache.scala 47:20]
  reg [52:0] tags1_13; // @[dcache.scala 47:20]
  reg [52:0] tags1_14; // @[dcache.scala 47:20]
  reg [52:0] tags1_15; // @[dcache.scala 47:20]
  reg [52:0] tags1_16; // @[dcache.scala 47:20]
  reg [52:0] tags1_17; // @[dcache.scala 47:20]
  reg [52:0] tags1_18; // @[dcache.scala 47:20]
  reg [52:0] tags1_19; // @[dcache.scala 47:20]
  reg [52:0] tags1_20; // @[dcache.scala 47:20]
  reg [52:0] tags1_21; // @[dcache.scala 47:20]
  reg [52:0] tags1_22; // @[dcache.scala 47:20]
  reg [52:0] tags1_23; // @[dcache.scala 47:20]
  reg [52:0] tags1_24; // @[dcache.scala 47:20]
  reg [52:0] tags1_25; // @[dcache.scala 47:20]
  reg [52:0] tags1_26; // @[dcache.scala 47:20]
  reg [52:0] tags1_27; // @[dcache.scala 47:20]
  reg [52:0] tags1_28; // @[dcache.scala 47:20]
  reg [52:0] tags1_29; // @[dcache.scala 47:20]
  reg [52:0] tags1_30; // @[dcache.scala 47:20]
  reg [52:0] tags1_31; // @[dcache.scala 47:20]
  reg [52:0] tags1_32; // @[dcache.scala 47:20]
  reg [52:0] tags1_33; // @[dcache.scala 47:20]
  reg [52:0] tags1_34; // @[dcache.scala 47:20]
  reg [52:0] tags1_35; // @[dcache.scala 47:20]
  reg [52:0] tags1_36; // @[dcache.scala 47:20]
  reg [52:0] tags1_37; // @[dcache.scala 47:20]
  reg [52:0] tags1_38; // @[dcache.scala 47:20]
  reg [52:0] tags1_39; // @[dcache.scala 47:20]
  reg [52:0] tags1_40; // @[dcache.scala 47:20]
  reg [52:0] tags1_41; // @[dcache.scala 47:20]
  reg [52:0] tags1_42; // @[dcache.scala 47:20]
  reg [52:0] tags1_43; // @[dcache.scala 47:20]
  reg [52:0] tags1_44; // @[dcache.scala 47:20]
  reg [52:0] tags1_45; // @[dcache.scala 47:20]
  reg [52:0] tags1_46; // @[dcache.scala 47:20]
  reg [52:0] tags1_47; // @[dcache.scala 47:20]
  reg [52:0] tags1_48; // @[dcache.scala 47:20]
  reg [52:0] tags1_49; // @[dcache.scala 47:20]
  reg [52:0] tags1_50; // @[dcache.scala 47:20]
  reg [52:0] tags1_51; // @[dcache.scala 47:20]
  reg [52:0] tags1_52; // @[dcache.scala 47:20]
  reg [52:0] tags1_53; // @[dcache.scala 47:20]
  reg [52:0] tags1_54; // @[dcache.scala 47:20]
  reg [52:0] tags1_55; // @[dcache.scala 47:20]
  reg [52:0] tags1_56; // @[dcache.scala 47:20]
  reg [52:0] tags1_57; // @[dcache.scala 47:20]
  reg [52:0] tags1_58; // @[dcache.scala 47:20]
  reg [52:0] tags1_59; // @[dcache.scala 47:20]
  reg [52:0] tags1_60; // @[dcache.scala 47:20]
  reg [52:0] tags1_61; // @[dcache.scala 47:20]
  reg [52:0] tags1_62; // @[dcache.scala 47:20]
  reg [52:0] tags1_63; // @[dcache.scala 47:20]
  reg [52:0] tags1_64; // @[dcache.scala 47:20]
  reg [52:0] tags1_65; // @[dcache.scala 47:20]
  reg [52:0] tags1_66; // @[dcache.scala 47:20]
  reg [52:0] tags1_67; // @[dcache.scala 47:20]
  reg [52:0] tags1_68; // @[dcache.scala 47:20]
  reg [52:0] tags1_69; // @[dcache.scala 47:20]
  reg [52:0] tags1_70; // @[dcache.scala 47:20]
  reg [52:0] tags1_71; // @[dcache.scala 47:20]
  reg [52:0] tags1_72; // @[dcache.scala 47:20]
  reg [52:0] tags1_73; // @[dcache.scala 47:20]
  reg [52:0] tags1_74; // @[dcache.scala 47:20]
  reg [52:0] tags1_75; // @[dcache.scala 47:20]
  reg [52:0] tags1_76; // @[dcache.scala 47:20]
  reg [52:0] tags1_77; // @[dcache.scala 47:20]
  reg [52:0] tags1_78; // @[dcache.scala 47:20]
  reg [52:0] tags1_79; // @[dcache.scala 47:20]
  reg [52:0] tags1_80; // @[dcache.scala 47:20]
  reg [52:0] tags1_81; // @[dcache.scala 47:20]
  reg [52:0] tags1_82; // @[dcache.scala 47:20]
  reg [52:0] tags1_83; // @[dcache.scala 47:20]
  reg [52:0] tags1_84; // @[dcache.scala 47:20]
  reg [52:0] tags1_85; // @[dcache.scala 47:20]
  reg [52:0] tags1_86; // @[dcache.scala 47:20]
  reg [52:0] tags1_87; // @[dcache.scala 47:20]
  reg [52:0] tags1_88; // @[dcache.scala 47:20]
  reg [52:0] tags1_89; // @[dcache.scala 47:20]
  reg [52:0] tags1_90; // @[dcache.scala 47:20]
  reg [52:0] tags1_91; // @[dcache.scala 47:20]
  reg [52:0] tags1_92; // @[dcache.scala 47:20]
  reg [52:0] tags1_93; // @[dcache.scala 47:20]
  reg [52:0] tags1_94; // @[dcache.scala 47:20]
  reg [52:0] tags1_95; // @[dcache.scala 47:20]
  reg [52:0] tags1_96; // @[dcache.scala 47:20]
  reg [52:0] tags1_97; // @[dcache.scala 47:20]
  reg [52:0] tags1_98; // @[dcache.scala 47:20]
  reg [52:0] tags1_99; // @[dcache.scala 47:20]
  reg [52:0] tags1_100; // @[dcache.scala 47:20]
  reg [52:0] tags1_101; // @[dcache.scala 47:20]
  reg [52:0] tags1_102; // @[dcache.scala 47:20]
  reg [52:0] tags1_103; // @[dcache.scala 47:20]
  reg [52:0] tags1_104; // @[dcache.scala 47:20]
  reg [52:0] tags1_105; // @[dcache.scala 47:20]
  reg [52:0] tags1_106; // @[dcache.scala 47:20]
  reg [52:0] tags1_107; // @[dcache.scala 47:20]
  reg [52:0] tags1_108; // @[dcache.scala 47:20]
  reg [52:0] tags1_109; // @[dcache.scala 47:20]
  reg [52:0] tags1_110; // @[dcache.scala 47:20]
  reg [52:0] tags1_111; // @[dcache.scala 47:20]
  reg [52:0] tags1_112; // @[dcache.scala 47:20]
  reg [52:0] tags1_113; // @[dcache.scala 47:20]
  reg [52:0] tags1_114; // @[dcache.scala 47:20]
  reg [52:0] tags1_115; // @[dcache.scala 47:20]
  reg [52:0] tags1_116; // @[dcache.scala 47:20]
  reg [52:0] tags1_117; // @[dcache.scala 47:20]
  reg [52:0] tags1_118; // @[dcache.scala 47:20]
  reg [52:0] tags1_119; // @[dcache.scala 47:20]
  reg [52:0] tags1_120; // @[dcache.scala 47:20]
  reg [52:0] tags1_121; // @[dcache.scala 47:20]
  reg [52:0] tags1_122; // @[dcache.scala 47:20]
  reg [52:0] tags1_123; // @[dcache.scala 47:20]
  reg [52:0] tags1_124; // @[dcache.scala 47:20]
  reg [52:0] tags1_125; // @[dcache.scala 47:20]
  reg [52:0] tags1_126; // @[dcache.scala 47:20]
  reg [52:0] tags1_127; // @[dcache.scala 47:20]
  reg  valid0_0; // @[dcache.scala 48:21]
  reg  valid0_1; // @[dcache.scala 48:21]
  reg  valid0_2; // @[dcache.scala 48:21]
  reg  valid0_3; // @[dcache.scala 48:21]
  reg  valid0_4; // @[dcache.scala 48:21]
  reg  valid0_5; // @[dcache.scala 48:21]
  reg  valid0_6; // @[dcache.scala 48:21]
  reg  valid0_7; // @[dcache.scala 48:21]
  reg  valid0_8; // @[dcache.scala 48:21]
  reg  valid0_9; // @[dcache.scala 48:21]
  reg  valid0_10; // @[dcache.scala 48:21]
  reg  valid0_11; // @[dcache.scala 48:21]
  reg  valid0_12; // @[dcache.scala 48:21]
  reg  valid0_13; // @[dcache.scala 48:21]
  reg  valid0_14; // @[dcache.scala 48:21]
  reg  valid0_15; // @[dcache.scala 48:21]
  reg  valid0_16; // @[dcache.scala 48:21]
  reg  valid0_17; // @[dcache.scala 48:21]
  reg  valid0_18; // @[dcache.scala 48:21]
  reg  valid0_19; // @[dcache.scala 48:21]
  reg  valid0_20; // @[dcache.scala 48:21]
  reg  valid0_21; // @[dcache.scala 48:21]
  reg  valid0_22; // @[dcache.scala 48:21]
  reg  valid0_23; // @[dcache.scala 48:21]
  reg  valid0_24; // @[dcache.scala 48:21]
  reg  valid0_25; // @[dcache.scala 48:21]
  reg  valid0_26; // @[dcache.scala 48:21]
  reg  valid0_27; // @[dcache.scala 48:21]
  reg  valid0_28; // @[dcache.scala 48:21]
  reg  valid0_29; // @[dcache.scala 48:21]
  reg  valid0_30; // @[dcache.scala 48:21]
  reg  valid0_31; // @[dcache.scala 48:21]
  reg  valid0_32; // @[dcache.scala 48:21]
  reg  valid0_33; // @[dcache.scala 48:21]
  reg  valid0_34; // @[dcache.scala 48:21]
  reg  valid0_35; // @[dcache.scala 48:21]
  reg  valid0_36; // @[dcache.scala 48:21]
  reg  valid0_37; // @[dcache.scala 48:21]
  reg  valid0_38; // @[dcache.scala 48:21]
  reg  valid0_39; // @[dcache.scala 48:21]
  reg  valid0_40; // @[dcache.scala 48:21]
  reg  valid0_41; // @[dcache.scala 48:21]
  reg  valid0_42; // @[dcache.scala 48:21]
  reg  valid0_43; // @[dcache.scala 48:21]
  reg  valid0_44; // @[dcache.scala 48:21]
  reg  valid0_45; // @[dcache.scala 48:21]
  reg  valid0_46; // @[dcache.scala 48:21]
  reg  valid0_47; // @[dcache.scala 48:21]
  reg  valid0_48; // @[dcache.scala 48:21]
  reg  valid0_49; // @[dcache.scala 48:21]
  reg  valid0_50; // @[dcache.scala 48:21]
  reg  valid0_51; // @[dcache.scala 48:21]
  reg  valid0_52; // @[dcache.scala 48:21]
  reg  valid0_53; // @[dcache.scala 48:21]
  reg  valid0_54; // @[dcache.scala 48:21]
  reg  valid0_55; // @[dcache.scala 48:21]
  reg  valid0_56; // @[dcache.scala 48:21]
  reg  valid0_57; // @[dcache.scala 48:21]
  reg  valid0_58; // @[dcache.scala 48:21]
  reg  valid0_59; // @[dcache.scala 48:21]
  reg  valid0_60; // @[dcache.scala 48:21]
  reg  valid0_61; // @[dcache.scala 48:21]
  reg  valid0_62; // @[dcache.scala 48:21]
  reg  valid0_63; // @[dcache.scala 48:21]
  reg  valid0_64; // @[dcache.scala 48:21]
  reg  valid0_65; // @[dcache.scala 48:21]
  reg  valid0_66; // @[dcache.scala 48:21]
  reg  valid0_67; // @[dcache.scala 48:21]
  reg  valid0_68; // @[dcache.scala 48:21]
  reg  valid0_69; // @[dcache.scala 48:21]
  reg  valid0_70; // @[dcache.scala 48:21]
  reg  valid0_71; // @[dcache.scala 48:21]
  reg  valid0_72; // @[dcache.scala 48:21]
  reg  valid0_73; // @[dcache.scala 48:21]
  reg  valid0_74; // @[dcache.scala 48:21]
  reg  valid0_75; // @[dcache.scala 48:21]
  reg  valid0_76; // @[dcache.scala 48:21]
  reg  valid0_77; // @[dcache.scala 48:21]
  reg  valid0_78; // @[dcache.scala 48:21]
  reg  valid0_79; // @[dcache.scala 48:21]
  reg  valid0_80; // @[dcache.scala 48:21]
  reg  valid0_81; // @[dcache.scala 48:21]
  reg  valid0_82; // @[dcache.scala 48:21]
  reg  valid0_83; // @[dcache.scala 48:21]
  reg  valid0_84; // @[dcache.scala 48:21]
  reg  valid0_85; // @[dcache.scala 48:21]
  reg  valid0_86; // @[dcache.scala 48:21]
  reg  valid0_87; // @[dcache.scala 48:21]
  reg  valid0_88; // @[dcache.scala 48:21]
  reg  valid0_89; // @[dcache.scala 48:21]
  reg  valid0_90; // @[dcache.scala 48:21]
  reg  valid0_91; // @[dcache.scala 48:21]
  reg  valid0_92; // @[dcache.scala 48:21]
  reg  valid0_93; // @[dcache.scala 48:21]
  reg  valid0_94; // @[dcache.scala 48:21]
  reg  valid0_95; // @[dcache.scala 48:21]
  reg  valid0_96; // @[dcache.scala 48:21]
  reg  valid0_97; // @[dcache.scala 48:21]
  reg  valid0_98; // @[dcache.scala 48:21]
  reg  valid0_99; // @[dcache.scala 48:21]
  reg  valid0_100; // @[dcache.scala 48:21]
  reg  valid0_101; // @[dcache.scala 48:21]
  reg  valid0_102; // @[dcache.scala 48:21]
  reg  valid0_103; // @[dcache.scala 48:21]
  reg  valid0_104; // @[dcache.scala 48:21]
  reg  valid0_105; // @[dcache.scala 48:21]
  reg  valid0_106; // @[dcache.scala 48:21]
  reg  valid0_107; // @[dcache.scala 48:21]
  reg  valid0_108; // @[dcache.scala 48:21]
  reg  valid0_109; // @[dcache.scala 48:21]
  reg  valid0_110; // @[dcache.scala 48:21]
  reg  valid0_111; // @[dcache.scala 48:21]
  reg  valid0_112; // @[dcache.scala 48:21]
  reg  valid0_113; // @[dcache.scala 48:21]
  reg  valid0_114; // @[dcache.scala 48:21]
  reg  valid0_115; // @[dcache.scala 48:21]
  reg  valid0_116; // @[dcache.scala 48:21]
  reg  valid0_117; // @[dcache.scala 48:21]
  reg  valid0_118; // @[dcache.scala 48:21]
  reg  valid0_119; // @[dcache.scala 48:21]
  reg  valid0_120; // @[dcache.scala 48:21]
  reg  valid0_121; // @[dcache.scala 48:21]
  reg  valid0_122; // @[dcache.scala 48:21]
  reg  valid0_123; // @[dcache.scala 48:21]
  reg  valid0_124; // @[dcache.scala 48:21]
  reg  valid0_125; // @[dcache.scala 48:21]
  reg  valid0_126; // @[dcache.scala 48:21]
  reg  valid0_127; // @[dcache.scala 48:21]
  reg  valid1_0; // @[dcache.scala 49:21]
  reg  valid1_1; // @[dcache.scala 49:21]
  reg  valid1_2; // @[dcache.scala 49:21]
  reg  valid1_3; // @[dcache.scala 49:21]
  reg  valid1_4; // @[dcache.scala 49:21]
  reg  valid1_5; // @[dcache.scala 49:21]
  reg  valid1_6; // @[dcache.scala 49:21]
  reg  valid1_7; // @[dcache.scala 49:21]
  reg  valid1_8; // @[dcache.scala 49:21]
  reg  valid1_9; // @[dcache.scala 49:21]
  reg  valid1_10; // @[dcache.scala 49:21]
  reg  valid1_11; // @[dcache.scala 49:21]
  reg  valid1_12; // @[dcache.scala 49:21]
  reg  valid1_13; // @[dcache.scala 49:21]
  reg  valid1_14; // @[dcache.scala 49:21]
  reg  valid1_15; // @[dcache.scala 49:21]
  reg  valid1_16; // @[dcache.scala 49:21]
  reg  valid1_17; // @[dcache.scala 49:21]
  reg  valid1_18; // @[dcache.scala 49:21]
  reg  valid1_19; // @[dcache.scala 49:21]
  reg  valid1_20; // @[dcache.scala 49:21]
  reg  valid1_21; // @[dcache.scala 49:21]
  reg  valid1_22; // @[dcache.scala 49:21]
  reg  valid1_23; // @[dcache.scala 49:21]
  reg  valid1_24; // @[dcache.scala 49:21]
  reg  valid1_25; // @[dcache.scala 49:21]
  reg  valid1_26; // @[dcache.scala 49:21]
  reg  valid1_27; // @[dcache.scala 49:21]
  reg  valid1_28; // @[dcache.scala 49:21]
  reg  valid1_29; // @[dcache.scala 49:21]
  reg  valid1_30; // @[dcache.scala 49:21]
  reg  valid1_31; // @[dcache.scala 49:21]
  reg  valid1_32; // @[dcache.scala 49:21]
  reg  valid1_33; // @[dcache.scala 49:21]
  reg  valid1_34; // @[dcache.scala 49:21]
  reg  valid1_35; // @[dcache.scala 49:21]
  reg  valid1_36; // @[dcache.scala 49:21]
  reg  valid1_37; // @[dcache.scala 49:21]
  reg  valid1_38; // @[dcache.scala 49:21]
  reg  valid1_39; // @[dcache.scala 49:21]
  reg  valid1_40; // @[dcache.scala 49:21]
  reg  valid1_41; // @[dcache.scala 49:21]
  reg  valid1_42; // @[dcache.scala 49:21]
  reg  valid1_43; // @[dcache.scala 49:21]
  reg  valid1_44; // @[dcache.scala 49:21]
  reg  valid1_45; // @[dcache.scala 49:21]
  reg  valid1_46; // @[dcache.scala 49:21]
  reg  valid1_47; // @[dcache.scala 49:21]
  reg  valid1_48; // @[dcache.scala 49:21]
  reg  valid1_49; // @[dcache.scala 49:21]
  reg  valid1_50; // @[dcache.scala 49:21]
  reg  valid1_51; // @[dcache.scala 49:21]
  reg  valid1_52; // @[dcache.scala 49:21]
  reg  valid1_53; // @[dcache.scala 49:21]
  reg  valid1_54; // @[dcache.scala 49:21]
  reg  valid1_55; // @[dcache.scala 49:21]
  reg  valid1_56; // @[dcache.scala 49:21]
  reg  valid1_57; // @[dcache.scala 49:21]
  reg  valid1_58; // @[dcache.scala 49:21]
  reg  valid1_59; // @[dcache.scala 49:21]
  reg  valid1_60; // @[dcache.scala 49:21]
  reg  valid1_61; // @[dcache.scala 49:21]
  reg  valid1_62; // @[dcache.scala 49:21]
  reg  valid1_63; // @[dcache.scala 49:21]
  reg  valid1_64; // @[dcache.scala 49:21]
  reg  valid1_65; // @[dcache.scala 49:21]
  reg  valid1_66; // @[dcache.scala 49:21]
  reg  valid1_67; // @[dcache.scala 49:21]
  reg  valid1_68; // @[dcache.scala 49:21]
  reg  valid1_69; // @[dcache.scala 49:21]
  reg  valid1_70; // @[dcache.scala 49:21]
  reg  valid1_71; // @[dcache.scala 49:21]
  reg  valid1_72; // @[dcache.scala 49:21]
  reg  valid1_73; // @[dcache.scala 49:21]
  reg  valid1_74; // @[dcache.scala 49:21]
  reg  valid1_75; // @[dcache.scala 49:21]
  reg  valid1_76; // @[dcache.scala 49:21]
  reg  valid1_77; // @[dcache.scala 49:21]
  reg  valid1_78; // @[dcache.scala 49:21]
  reg  valid1_79; // @[dcache.scala 49:21]
  reg  valid1_80; // @[dcache.scala 49:21]
  reg  valid1_81; // @[dcache.scala 49:21]
  reg  valid1_82; // @[dcache.scala 49:21]
  reg  valid1_83; // @[dcache.scala 49:21]
  reg  valid1_84; // @[dcache.scala 49:21]
  reg  valid1_85; // @[dcache.scala 49:21]
  reg  valid1_86; // @[dcache.scala 49:21]
  reg  valid1_87; // @[dcache.scala 49:21]
  reg  valid1_88; // @[dcache.scala 49:21]
  reg  valid1_89; // @[dcache.scala 49:21]
  reg  valid1_90; // @[dcache.scala 49:21]
  reg  valid1_91; // @[dcache.scala 49:21]
  reg  valid1_92; // @[dcache.scala 49:21]
  reg  valid1_93; // @[dcache.scala 49:21]
  reg  valid1_94; // @[dcache.scala 49:21]
  reg  valid1_95; // @[dcache.scala 49:21]
  reg  valid1_96; // @[dcache.scala 49:21]
  reg  valid1_97; // @[dcache.scala 49:21]
  reg  valid1_98; // @[dcache.scala 49:21]
  reg  valid1_99; // @[dcache.scala 49:21]
  reg  valid1_100; // @[dcache.scala 49:21]
  reg  valid1_101; // @[dcache.scala 49:21]
  reg  valid1_102; // @[dcache.scala 49:21]
  reg  valid1_103; // @[dcache.scala 49:21]
  reg  valid1_104; // @[dcache.scala 49:21]
  reg  valid1_105; // @[dcache.scala 49:21]
  reg  valid1_106; // @[dcache.scala 49:21]
  reg  valid1_107; // @[dcache.scala 49:21]
  reg  valid1_108; // @[dcache.scala 49:21]
  reg  valid1_109; // @[dcache.scala 49:21]
  reg  valid1_110; // @[dcache.scala 49:21]
  reg  valid1_111; // @[dcache.scala 49:21]
  reg  valid1_112; // @[dcache.scala 49:21]
  reg  valid1_113; // @[dcache.scala 49:21]
  reg  valid1_114; // @[dcache.scala 49:21]
  reg  valid1_115; // @[dcache.scala 49:21]
  reg  valid1_116; // @[dcache.scala 49:21]
  reg  valid1_117; // @[dcache.scala 49:21]
  reg  valid1_118; // @[dcache.scala 49:21]
  reg  valid1_119; // @[dcache.scala 49:21]
  reg  valid1_120; // @[dcache.scala 49:21]
  reg  valid1_121; // @[dcache.scala 49:21]
  reg  valid1_122; // @[dcache.scala 49:21]
  reg  valid1_123; // @[dcache.scala 49:21]
  reg  valid1_124; // @[dcache.scala 49:21]
  reg  valid1_125; // @[dcache.scala 49:21]
  reg  valid1_126; // @[dcache.scala 49:21]
  reg  valid1_127; // @[dcache.scala 49:21]
  reg  dirty0_0; // @[dcache.scala 50:21]
  reg  dirty0_1; // @[dcache.scala 50:21]
  reg  dirty0_2; // @[dcache.scala 50:21]
  reg  dirty0_3; // @[dcache.scala 50:21]
  reg  dirty0_4; // @[dcache.scala 50:21]
  reg  dirty0_5; // @[dcache.scala 50:21]
  reg  dirty0_6; // @[dcache.scala 50:21]
  reg  dirty0_7; // @[dcache.scala 50:21]
  reg  dirty0_8; // @[dcache.scala 50:21]
  reg  dirty0_9; // @[dcache.scala 50:21]
  reg  dirty0_10; // @[dcache.scala 50:21]
  reg  dirty0_11; // @[dcache.scala 50:21]
  reg  dirty0_12; // @[dcache.scala 50:21]
  reg  dirty0_13; // @[dcache.scala 50:21]
  reg  dirty0_14; // @[dcache.scala 50:21]
  reg  dirty0_15; // @[dcache.scala 50:21]
  reg  dirty0_16; // @[dcache.scala 50:21]
  reg  dirty0_17; // @[dcache.scala 50:21]
  reg  dirty0_18; // @[dcache.scala 50:21]
  reg  dirty0_19; // @[dcache.scala 50:21]
  reg  dirty0_20; // @[dcache.scala 50:21]
  reg  dirty0_21; // @[dcache.scala 50:21]
  reg  dirty0_22; // @[dcache.scala 50:21]
  reg  dirty0_23; // @[dcache.scala 50:21]
  reg  dirty0_24; // @[dcache.scala 50:21]
  reg  dirty0_25; // @[dcache.scala 50:21]
  reg  dirty0_26; // @[dcache.scala 50:21]
  reg  dirty0_27; // @[dcache.scala 50:21]
  reg  dirty0_28; // @[dcache.scala 50:21]
  reg  dirty0_29; // @[dcache.scala 50:21]
  reg  dirty0_30; // @[dcache.scala 50:21]
  reg  dirty0_31; // @[dcache.scala 50:21]
  reg  dirty0_32; // @[dcache.scala 50:21]
  reg  dirty0_33; // @[dcache.scala 50:21]
  reg  dirty0_34; // @[dcache.scala 50:21]
  reg  dirty0_35; // @[dcache.scala 50:21]
  reg  dirty0_36; // @[dcache.scala 50:21]
  reg  dirty0_37; // @[dcache.scala 50:21]
  reg  dirty0_38; // @[dcache.scala 50:21]
  reg  dirty0_39; // @[dcache.scala 50:21]
  reg  dirty0_40; // @[dcache.scala 50:21]
  reg  dirty0_41; // @[dcache.scala 50:21]
  reg  dirty0_42; // @[dcache.scala 50:21]
  reg  dirty0_43; // @[dcache.scala 50:21]
  reg  dirty0_44; // @[dcache.scala 50:21]
  reg  dirty0_45; // @[dcache.scala 50:21]
  reg  dirty0_46; // @[dcache.scala 50:21]
  reg  dirty0_47; // @[dcache.scala 50:21]
  reg  dirty0_48; // @[dcache.scala 50:21]
  reg  dirty0_49; // @[dcache.scala 50:21]
  reg  dirty0_50; // @[dcache.scala 50:21]
  reg  dirty0_51; // @[dcache.scala 50:21]
  reg  dirty0_52; // @[dcache.scala 50:21]
  reg  dirty0_53; // @[dcache.scala 50:21]
  reg  dirty0_54; // @[dcache.scala 50:21]
  reg  dirty0_55; // @[dcache.scala 50:21]
  reg  dirty0_56; // @[dcache.scala 50:21]
  reg  dirty0_57; // @[dcache.scala 50:21]
  reg  dirty0_58; // @[dcache.scala 50:21]
  reg  dirty0_59; // @[dcache.scala 50:21]
  reg  dirty0_60; // @[dcache.scala 50:21]
  reg  dirty0_61; // @[dcache.scala 50:21]
  reg  dirty0_62; // @[dcache.scala 50:21]
  reg  dirty0_63; // @[dcache.scala 50:21]
  reg  dirty0_64; // @[dcache.scala 50:21]
  reg  dirty0_65; // @[dcache.scala 50:21]
  reg  dirty0_66; // @[dcache.scala 50:21]
  reg  dirty0_67; // @[dcache.scala 50:21]
  reg  dirty0_68; // @[dcache.scala 50:21]
  reg  dirty0_69; // @[dcache.scala 50:21]
  reg  dirty0_70; // @[dcache.scala 50:21]
  reg  dirty0_71; // @[dcache.scala 50:21]
  reg  dirty0_72; // @[dcache.scala 50:21]
  reg  dirty0_73; // @[dcache.scala 50:21]
  reg  dirty0_74; // @[dcache.scala 50:21]
  reg  dirty0_75; // @[dcache.scala 50:21]
  reg  dirty0_76; // @[dcache.scala 50:21]
  reg  dirty0_77; // @[dcache.scala 50:21]
  reg  dirty0_78; // @[dcache.scala 50:21]
  reg  dirty0_79; // @[dcache.scala 50:21]
  reg  dirty0_80; // @[dcache.scala 50:21]
  reg  dirty0_81; // @[dcache.scala 50:21]
  reg  dirty0_82; // @[dcache.scala 50:21]
  reg  dirty0_83; // @[dcache.scala 50:21]
  reg  dirty0_84; // @[dcache.scala 50:21]
  reg  dirty0_85; // @[dcache.scala 50:21]
  reg  dirty0_86; // @[dcache.scala 50:21]
  reg  dirty0_87; // @[dcache.scala 50:21]
  reg  dirty0_88; // @[dcache.scala 50:21]
  reg  dirty0_89; // @[dcache.scala 50:21]
  reg  dirty0_90; // @[dcache.scala 50:21]
  reg  dirty0_91; // @[dcache.scala 50:21]
  reg  dirty0_92; // @[dcache.scala 50:21]
  reg  dirty0_93; // @[dcache.scala 50:21]
  reg  dirty0_94; // @[dcache.scala 50:21]
  reg  dirty0_95; // @[dcache.scala 50:21]
  reg  dirty0_96; // @[dcache.scala 50:21]
  reg  dirty0_97; // @[dcache.scala 50:21]
  reg  dirty0_98; // @[dcache.scala 50:21]
  reg  dirty0_99; // @[dcache.scala 50:21]
  reg  dirty0_100; // @[dcache.scala 50:21]
  reg  dirty0_101; // @[dcache.scala 50:21]
  reg  dirty0_102; // @[dcache.scala 50:21]
  reg  dirty0_103; // @[dcache.scala 50:21]
  reg  dirty0_104; // @[dcache.scala 50:21]
  reg  dirty0_105; // @[dcache.scala 50:21]
  reg  dirty0_106; // @[dcache.scala 50:21]
  reg  dirty0_107; // @[dcache.scala 50:21]
  reg  dirty0_108; // @[dcache.scala 50:21]
  reg  dirty0_109; // @[dcache.scala 50:21]
  reg  dirty0_110; // @[dcache.scala 50:21]
  reg  dirty0_111; // @[dcache.scala 50:21]
  reg  dirty0_112; // @[dcache.scala 50:21]
  reg  dirty0_113; // @[dcache.scala 50:21]
  reg  dirty0_114; // @[dcache.scala 50:21]
  reg  dirty0_115; // @[dcache.scala 50:21]
  reg  dirty0_116; // @[dcache.scala 50:21]
  reg  dirty0_117; // @[dcache.scala 50:21]
  reg  dirty0_118; // @[dcache.scala 50:21]
  reg  dirty0_119; // @[dcache.scala 50:21]
  reg  dirty0_120; // @[dcache.scala 50:21]
  reg  dirty0_121; // @[dcache.scala 50:21]
  reg  dirty0_122; // @[dcache.scala 50:21]
  reg  dirty0_123; // @[dcache.scala 50:21]
  reg  dirty0_124; // @[dcache.scala 50:21]
  reg  dirty0_125; // @[dcache.scala 50:21]
  reg  dirty0_126; // @[dcache.scala 50:21]
  reg  dirty0_127; // @[dcache.scala 50:21]
  reg  dirty1_0; // @[dcache.scala 51:21]
  reg  dirty1_1; // @[dcache.scala 51:21]
  reg  dirty1_2; // @[dcache.scala 51:21]
  reg  dirty1_3; // @[dcache.scala 51:21]
  reg  dirty1_4; // @[dcache.scala 51:21]
  reg  dirty1_5; // @[dcache.scala 51:21]
  reg  dirty1_6; // @[dcache.scala 51:21]
  reg  dirty1_7; // @[dcache.scala 51:21]
  reg  dirty1_8; // @[dcache.scala 51:21]
  reg  dirty1_9; // @[dcache.scala 51:21]
  reg  dirty1_10; // @[dcache.scala 51:21]
  reg  dirty1_11; // @[dcache.scala 51:21]
  reg  dirty1_12; // @[dcache.scala 51:21]
  reg  dirty1_13; // @[dcache.scala 51:21]
  reg  dirty1_14; // @[dcache.scala 51:21]
  reg  dirty1_15; // @[dcache.scala 51:21]
  reg  dirty1_16; // @[dcache.scala 51:21]
  reg  dirty1_17; // @[dcache.scala 51:21]
  reg  dirty1_18; // @[dcache.scala 51:21]
  reg  dirty1_19; // @[dcache.scala 51:21]
  reg  dirty1_20; // @[dcache.scala 51:21]
  reg  dirty1_21; // @[dcache.scala 51:21]
  reg  dirty1_22; // @[dcache.scala 51:21]
  reg  dirty1_23; // @[dcache.scala 51:21]
  reg  dirty1_24; // @[dcache.scala 51:21]
  reg  dirty1_25; // @[dcache.scala 51:21]
  reg  dirty1_26; // @[dcache.scala 51:21]
  reg  dirty1_27; // @[dcache.scala 51:21]
  reg  dirty1_28; // @[dcache.scala 51:21]
  reg  dirty1_29; // @[dcache.scala 51:21]
  reg  dirty1_30; // @[dcache.scala 51:21]
  reg  dirty1_31; // @[dcache.scala 51:21]
  reg  dirty1_32; // @[dcache.scala 51:21]
  reg  dirty1_33; // @[dcache.scala 51:21]
  reg  dirty1_34; // @[dcache.scala 51:21]
  reg  dirty1_35; // @[dcache.scala 51:21]
  reg  dirty1_36; // @[dcache.scala 51:21]
  reg  dirty1_37; // @[dcache.scala 51:21]
  reg  dirty1_38; // @[dcache.scala 51:21]
  reg  dirty1_39; // @[dcache.scala 51:21]
  reg  dirty1_40; // @[dcache.scala 51:21]
  reg  dirty1_41; // @[dcache.scala 51:21]
  reg  dirty1_42; // @[dcache.scala 51:21]
  reg  dirty1_43; // @[dcache.scala 51:21]
  reg  dirty1_44; // @[dcache.scala 51:21]
  reg  dirty1_45; // @[dcache.scala 51:21]
  reg  dirty1_46; // @[dcache.scala 51:21]
  reg  dirty1_47; // @[dcache.scala 51:21]
  reg  dirty1_48; // @[dcache.scala 51:21]
  reg  dirty1_49; // @[dcache.scala 51:21]
  reg  dirty1_50; // @[dcache.scala 51:21]
  reg  dirty1_51; // @[dcache.scala 51:21]
  reg  dirty1_52; // @[dcache.scala 51:21]
  reg  dirty1_53; // @[dcache.scala 51:21]
  reg  dirty1_54; // @[dcache.scala 51:21]
  reg  dirty1_55; // @[dcache.scala 51:21]
  reg  dirty1_56; // @[dcache.scala 51:21]
  reg  dirty1_57; // @[dcache.scala 51:21]
  reg  dirty1_58; // @[dcache.scala 51:21]
  reg  dirty1_59; // @[dcache.scala 51:21]
  reg  dirty1_60; // @[dcache.scala 51:21]
  reg  dirty1_61; // @[dcache.scala 51:21]
  reg  dirty1_62; // @[dcache.scala 51:21]
  reg  dirty1_63; // @[dcache.scala 51:21]
  reg  dirty1_64; // @[dcache.scala 51:21]
  reg  dirty1_65; // @[dcache.scala 51:21]
  reg  dirty1_66; // @[dcache.scala 51:21]
  reg  dirty1_67; // @[dcache.scala 51:21]
  reg  dirty1_68; // @[dcache.scala 51:21]
  reg  dirty1_69; // @[dcache.scala 51:21]
  reg  dirty1_70; // @[dcache.scala 51:21]
  reg  dirty1_71; // @[dcache.scala 51:21]
  reg  dirty1_72; // @[dcache.scala 51:21]
  reg  dirty1_73; // @[dcache.scala 51:21]
  reg  dirty1_74; // @[dcache.scala 51:21]
  reg  dirty1_75; // @[dcache.scala 51:21]
  reg  dirty1_76; // @[dcache.scala 51:21]
  reg  dirty1_77; // @[dcache.scala 51:21]
  reg  dirty1_78; // @[dcache.scala 51:21]
  reg  dirty1_79; // @[dcache.scala 51:21]
  reg  dirty1_80; // @[dcache.scala 51:21]
  reg  dirty1_81; // @[dcache.scala 51:21]
  reg  dirty1_82; // @[dcache.scala 51:21]
  reg  dirty1_83; // @[dcache.scala 51:21]
  reg  dirty1_84; // @[dcache.scala 51:21]
  reg  dirty1_85; // @[dcache.scala 51:21]
  reg  dirty1_86; // @[dcache.scala 51:21]
  reg  dirty1_87; // @[dcache.scala 51:21]
  reg  dirty1_88; // @[dcache.scala 51:21]
  reg  dirty1_89; // @[dcache.scala 51:21]
  reg  dirty1_90; // @[dcache.scala 51:21]
  reg  dirty1_91; // @[dcache.scala 51:21]
  reg  dirty1_92; // @[dcache.scala 51:21]
  reg  dirty1_93; // @[dcache.scala 51:21]
  reg  dirty1_94; // @[dcache.scala 51:21]
  reg  dirty1_95; // @[dcache.scala 51:21]
  reg  dirty1_96; // @[dcache.scala 51:21]
  reg  dirty1_97; // @[dcache.scala 51:21]
  reg  dirty1_98; // @[dcache.scala 51:21]
  reg  dirty1_99; // @[dcache.scala 51:21]
  reg  dirty1_100; // @[dcache.scala 51:21]
  reg  dirty1_101; // @[dcache.scala 51:21]
  reg  dirty1_102; // @[dcache.scala 51:21]
  reg  dirty1_103; // @[dcache.scala 51:21]
  reg  dirty1_104; // @[dcache.scala 51:21]
  reg  dirty1_105; // @[dcache.scala 51:21]
  reg  dirty1_106; // @[dcache.scala 51:21]
  reg  dirty1_107; // @[dcache.scala 51:21]
  reg  dirty1_108; // @[dcache.scala 51:21]
  reg  dirty1_109; // @[dcache.scala 51:21]
  reg  dirty1_110; // @[dcache.scala 51:21]
  reg  dirty1_111; // @[dcache.scala 51:21]
  reg  dirty1_112; // @[dcache.scala 51:21]
  reg  dirty1_113; // @[dcache.scala 51:21]
  reg  dirty1_114; // @[dcache.scala 51:21]
  reg  dirty1_115; // @[dcache.scala 51:21]
  reg  dirty1_116; // @[dcache.scala 51:21]
  reg  dirty1_117; // @[dcache.scala 51:21]
  reg  dirty1_118; // @[dcache.scala 51:21]
  reg  dirty1_119; // @[dcache.scala 51:21]
  reg  dirty1_120; // @[dcache.scala 51:21]
  reg  dirty1_121; // @[dcache.scala 51:21]
  reg  dirty1_122; // @[dcache.scala 51:21]
  reg  dirty1_123; // @[dcache.scala 51:21]
  reg  dirty1_124; // @[dcache.scala 51:21]
  reg  dirty1_125; // @[dcache.scala 51:21]
  reg  dirty1_126; // @[dcache.scala 51:21]
  reg  dirty1_127; // @[dcache.scala 51:21]
  reg  victim; // @[dcache.scala 59:17]
  reg [127:0] read_from_mem_buf; // @[dcache.scala 61:32]
  reg [2:0] write_state; // @[dcache.scala 68:26]
  reg [1:0] state; // @[dcache.scala 72:20]
  wire  write_done = io_mem_master_writeResp_valid & io_mem_master_writeResp_ready; // @[dcache.scala 75:49]
  wire  read_done = io_mem_master_readData_valid & io_mem_master_readData_ready; // @[dcache.scala 76:47]
  wire  _should_write_back_T = state == 2'h2; // @[dcache.scala 79:29]
  wire  _uncache_T_3 = cpu_mem_Maddr == 64'ha000004c; // @[dcache.scala 128:20]
  wire  _uncache_T_4 = cpu_mem_Maddr == 64'ha0000048 | _uncache_T_3; // @[dcache.scala 127:38]
  wire  _uncache_T_5 = cpu_mem_Maddr == 64'ha0000060; // @[dcache.scala 129:20]
  wire  _uncache_T_6 = _uncache_T_4 | _uncache_T_5; // @[dcache.scala 128:42]
  wire  _uncache_T_7 = cpu_mem_Maddr == 64'ha0000100; // @[dcache.scala 130:20]
  wire  _uncache_T_8 = _uncache_T_6 | _uncache_T_7; // @[dcache.scala 129:38]
  wire  _uncache_T_11 = cpu_mem_Maddr == 64'ha0000102; // @[dcache.scala 131:20]
  wire  _uncache_T_12 = _uncache_T_8 | _uncache_T_11; // @[dcache.scala 130:37]
  wire  _uncache_T_15 = cpu_mem_Maddr == 64'ha0000104; // @[dcache.scala 132:20]
  wire  _uncache_T_16 = _uncache_T_12 | _uncache_T_15; // @[dcache.scala 131:41]
  wire  _uncache_T_19 = cpu_mem_Maddr >= 64'ha1000000 & cpu_mem_Maddr < VGA_MEM_BLK_E; // @[dcache.scala 133:38]
  wire  uncache = _uncache_T_16 | _uncache_T_19; // @[dcache.scala 132:41]
  wire  _should_write_back_T_3 = ~uncache; // @[dcache.scala 79:106]
  wire [6:0] index = cpu_mem_Maddr[10:4]; // @[dcache.scala 115:23]
  wire  _GEN_1 = 7'h1 == index ? valid1_1 : valid1_0; // @[dcache.scala 80:{46,46}]
  wire  _GEN_2 = 7'h2 == index ? valid1_2 : _GEN_1; // @[dcache.scala 80:{46,46}]
  wire  _GEN_3 = 7'h3 == index ? valid1_3 : _GEN_2; // @[dcache.scala 80:{46,46}]
  wire  _GEN_4 = 7'h4 == index ? valid1_4 : _GEN_3; // @[dcache.scala 80:{46,46}]
  wire  _GEN_5 = 7'h5 == index ? valid1_5 : _GEN_4; // @[dcache.scala 80:{46,46}]
  wire  _GEN_6 = 7'h6 == index ? valid1_6 : _GEN_5; // @[dcache.scala 80:{46,46}]
  wire  _GEN_7 = 7'h7 == index ? valid1_7 : _GEN_6; // @[dcache.scala 80:{46,46}]
  wire  _GEN_8 = 7'h8 == index ? valid1_8 : _GEN_7; // @[dcache.scala 80:{46,46}]
  wire  _GEN_9 = 7'h9 == index ? valid1_9 : _GEN_8; // @[dcache.scala 80:{46,46}]
  wire  _GEN_10 = 7'ha == index ? valid1_10 : _GEN_9; // @[dcache.scala 80:{46,46}]
  wire  _GEN_11 = 7'hb == index ? valid1_11 : _GEN_10; // @[dcache.scala 80:{46,46}]
  wire  _GEN_12 = 7'hc == index ? valid1_12 : _GEN_11; // @[dcache.scala 80:{46,46}]
  wire  _GEN_13 = 7'hd == index ? valid1_13 : _GEN_12; // @[dcache.scala 80:{46,46}]
  wire  _GEN_14 = 7'he == index ? valid1_14 : _GEN_13; // @[dcache.scala 80:{46,46}]
  wire  _GEN_15 = 7'hf == index ? valid1_15 : _GEN_14; // @[dcache.scala 80:{46,46}]
  wire  _GEN_16 = 7'h10 == index ? valid1_16 : _GEN_15; // @[dcache.scala 80:{46,46}]
  wire  _GEN_17 = 7'h11 == index ? valid1_17 : _GEN_16; // @[dcache.scala 80:{46,46}]
  wire  _GEN_18 = 7'h12 == index ? valid1_18 : _GEN_17; // @[dcache.scala 80:{46,46}]
  wire  _GEN_19 = 7'h13 == index ? valid1_19 : _GEN_18; // @[dcache.scala 80:{46,46}]
  wire  _GEN_20 = 7'h14 == index ? valid1_20 : _GEN_19; // @[dcache.scala 80:{46,46}]
  wire  _GEN_21 = 7'h15 == index ? valid1_21 : _GEN_20; // @[dcache.scala 80:{46,46}]
  wire  _GEN_22 = 7'h16 == index ? valid1_22 : _GEN_21; // @[dcache.scala 80:{46,46}]
  wire  _GEN_23 = 7'h17 == index ? valid1_23 : _GEN_22; // @[dcache.scala 80:{46,46}]
  wire  _GEN_24 = 7'h18 == index ? valid1_24 : _GEN_23; // @[dcache.scala 80:{46,46}]
  wire  _GEN_25 = 7'h19 == index ? valid1_25 : _GEN_24; // @[dcache.scala 80:{46,46}]
  wire  _GEN_26 = 7'h1a == index ? valid1_26 : _GEN_25; // @[dcache.scala 80:{46,46}]
  wire  _GEN_27 = 7'h1b == index ? valid1_27 : _GEN_26; // @[dcache.scala 80:{46,46}]
  wire  _GEN_28 = 7'h1c == index ? valid1_28 : _GEN_27; // @[dcache.scala 80:{46,46}]
  wire  _GEN_29 = 7'h1d == index ? valid1_29 : _GEN_28; // @[dcache.scala 80:{46,46}]
  wire  _GEN_30 = 7'h1e == index ? valid1_30 : _GEN_29; // @[dcache.scala 80:{46,46}]
  wire  _GEN_31 = 7'h1f == index ? valid1_31 : _GEN_30; // @[dcache.scala 80:{46,46}]
  wire  _GEN_32 = 7'h20 == index ? valid1_32 : _GEN_31; // @[dcache.scala 80:{46,46}]
  wire  _GEN_33 = 7'h21 == index ? valid1_33 : _GEN_32; // @[dcache.scala 80:{46,46}]
  wire  _GEN_34 = 7'h22 == index ? valid1_34 : _GEN_33; // @[dcache.scala 80:{46,46}]
  wire  _GEN_35 = 7'h23 == index ? valid1_35 : _GEN_34; // @[dcache.scala 80:{46,46}]
  wire  _GEN_36 = 7'h24 == index ? valid1_36 : _GEN_35; // @[dcache.scala 80:{46,46}]
  wire  _GEN_37 = 7'h25 == index ? valid1_37 : _GEN_36; // @[dcache.scala 80:{46,46}]
  wire  _GEN_38 = 7'h26 == index ? valid1_38 : _GEN_37; // @[dcache.scala 80:{46,46}]
  wire  _GEN_39 = 7'h27 == index ? valid1_39 : _GEN_38; // @[dcache.scala 80:{46,46}]
  wire  _GEN_40 = 7'h28 == index ? valid1_40 : _GEN_39; // @[dcache.scala 80:{46,46}]
  wire  _GEN_41 = 7'h29 == index ? valid1_41 : _GEN_40; // @[dcache.scala 80:{46,46}]
  wire  _GEN_42 = 7'h2a == index ? valid1_42 : _GEN_41; // @[dcache.scala 80:{46,46}]
  wire  _GEN_43 = 7'h2b == index ? valid1_43 : _GEN_42; // @[dcache.scala 80:{46,46}]
  wire  _GEN_44 = 7'h2c == index ? valid1_44 : _GEN_43; // @[dcache.scala 80:{46,46}]
  wire  _GEN_45 = 7'h2d == index ? valid1_45 : _GEN_44; // @[dcache.scala 80:{46,46}]
  wire  _GEN_46 = 7'h2e == index ? valid1_46 : _GEN_45; // @[dcache.scala 80:{46,46}]
  wire  _GEN_47 = 7'h2f == index ? valid1_47 : _GEN_46; // @[dcache.scala 80:{46,46}]
  wire  _GEN_48 = 7'h30 == index ? valid1_48 : _GEN_47; // @[dcache.scala 80:{46,46}]
  wire  _GEN_49 = 7'h31 == index ? valid1_49 : _GEN_48; // @[dcache.scala 80:{46,46}]
  wire  _GEN_50 = 7'h32 == index ? valid1_50 : _GEN_49; // @[dcache.scala 80:{46,46}]
  wire  _GEN_51 = 7'h33 == index ? valid1_51 : _GEN_50; // @[dcache.scala 80:{46,46}]
  wire  _GEN_52 = 7'h34 == index ? valid1_52 : _GEN_51; // @[dcache.scala 80:{46,46}]
  wire  _GEN_53 = 7'h35 == index ? valid1_53 : _GEN_52; // @[dcache.scala 80:{46,46}]
  wire  _GEN_54 = 7'h36 == index ? valid1_54 : _GEN_53; // @[dcache.scala 80:{46,46}]
  wire  _GEN_55 = 7'h37 == index ? valid1_55 : _GEN_54; // @[dcache.scala 80:{46,46}]
  wire  _GEN_56 = 7'h38 == index ? valid1_56 : _GEN_55; // @[dcache.scala 80:{46,46}]
  wire  _GEN_57 = 7'h39 == index ? valid1_57 : _GEN_56; // @[dcache.scala 80:{46,46}]
  wire  _GEN_58 = 7'h3a == index ? valid1_58 : _GEN_57; // @[dcache.scala 80:{46,46}]
  wire  _GEN_59 = 7'h3b == index ? valid1_59 : _GEN_58; // @[dcache.scala 80:{46,46}]
  wire  _GEN_60 = 7'h3c == index ? valid1_60 : _GEN_59; // @[dcache.scala 80:{46,46}]
  wire  _GEN_61 = 7'h3d == index ? valid1_61 : _GEN_60; // @[dcache.scala 80:{46,46}]
  wire  _GEN_62 = 7'h3e == index ? valid1_62 : _GEN_61; // @[dcache.scala 80:{46,46}]
  wire  _GEN_63 = 7'h3f == index ? valid1_63 : _GEN_62; // @[dcache.scala 80:{46,46}]
  wire  _GEN_64 = 7'h40 == index ? valid1_64 : _GEN_63; // @[dcache.scala 80:{46,46}]
  wire  _GEN_65 = 7'h41 == index ? valid1_65 : _GEN_64; // @[dcache.scala 80:{46,46}]
  wire  _GEN_66 = 7'h42 == index ? valid1_66 : _GEN_65; // @[dcache.scala 80:{46,46}]
  wire  _GEN_67 = 7'h43 == index ? valid1_67 : _GEN_66; // @[dcache.scala 80:{46,46}]
  wire  _GEN_68 = 7'h44 == index ? valid1_68 : _GEN_67; // @[dcache.scala 80:{46,46}]
  wire  _GEN_69 = 7'h45 == index ? valid1_69 : _GEN_68; // @[dcache.scala 80:{46,46}]
  wire  _GEN_70 = 7'h46 == index ? valid1_70 : _GEN_69; // @[dcache.scala 80:{46,46}]
  wire  _GEN_71 = 7'h47 == index ? valid1_71 : _GEN_70; // @[dcache.scala 80:{46,46}]
  wire  _GEN_72 = 7'h48 == index ? valid1_72 : _GEN_71; // @[dcache.scala 80:{46,46}]
  wire  _GEN_73 = 7'h49 == index ? valid1_73 : _GEN_72; // @[dcache.scala 80:{46,46}]
  wire  _GEN_74 = 7'h4a == index ? valid1_74 : _GEN_73; // @[dcache.scala 80:{46,46}]
  wire  _GEN_75 = 7'h4b == index ? valid1_75 : _GEN_74; // @[dcache.scala 80:{46,46}]
  wire  _GEN_76 = 7'h4c == index ? valid1_76 : _GEN_75; // @[dcache.scala 80:{46,46}]
  wire  _GEN_77 = 7'h4d == index ? valid1_77 : _GEN_76; // @[dcache.scala 80:{46,46}]
  wire  _GEN_78 = 7'h4e == index ? valid1_78 : _GEN_77; // @[dcache.scala 80:{46,46}]
  wire  _GEN_79 = 7'h4f == index ? valid1_79 : _GEN_78; // @[dcache.scala 80:{46,46}]
  wire  _GEN_80 = 7'h50 == index ? valid1_80 : _GEN_79; // @[dcache.scala 80:{46,46}]
  wire  _GEN_81 = 7'h51 == index ? valid1_81 : _GEN_80; // @[dcache.scala 80:{46,46}]
  wire  _GEN_82 = 7'h52 == index ? valid1_82 : _GEN_81; // @[dcache.scala 80:{46,46}]
  wire  _GEN_83 = 7'h53 == index ? valid1_83 : _GEN_82; // @[dcache.scala 80:{46,46}]
  wire  _GEN_84 = 7'h54 == index ? valid1_84 : _GEN_83; // @[dcache.scala 80:{46,46}]
  wire  _GEN_85 = 7'h55 == index ? valid1_85 : _GEN_84; // @[dcache.scala 80:{46,46}]
  wire  _GEN_86 = 7'h56 == index ? valid1_86 : _GEN_85; // @[dcache.scala 80:{46,46}]
  wire  _GEN_87 = 7'h57 == index ? valid1_87 : _GEN_86; // @[dcache.scala 80:{46,46}]
  wire  _GEN_88 = 7'h58 == index ? valid1_88 : _GEN_87; // @[dcache.scala 80:{46,46}]
  wire  _GEN_89 = 7'h59 == index ? valid1_89 : _GEN_88; // @[dcache.scala 80:{46,46}]
  wire  _GEN_90 = 7'h5a == index ? valid1_90 : _GEN_89; // @[dcache.scala 80:{46,46}]
  wire  _GEN_91 = 7'h5b == index ? valid1_91 : _GEN_90; // @[dcache.scala 80:{46,46}]
  wire  _GEN_92 = 7'h5c == index ? valid1_92 : _GEN_91; // @[dcache.scala 80:{46,46}]
  wire  _GEN_93 = 7'h5d == index ? valid1_93 : _GEN_92; // @[dcache.scala 80:{46,46}]
  wire  _GEN_94 = 7'h5e == index ? valid1_94 : _GEN_93; // @[dcache.scala 80:{46,46}]
  wire  _GEN_95 = 7'h5f == index ? valid1_95 : _GEN_94; // @[dcache.scala 80:{46,46}]
  wire  _GEN_96 = 7'h60 == index ? valid1_96 : _GEN_95; // @[dcache.scala 80:{46,46}]
  wire  _GEN_97 = 7'h61 == index ? valid1_97 : _GEN_96; // @[dcache.scala 80:{46,46}]
  wire  _GEN_98 = 7'h62 == index ? valid1_98 : _GEN_97; // @[dcache.scala 80:{46,46}]
  wire  _GEN_99 = 7'h63 == index ? valid1_99 : _GEN_98; // @[dcache.scala 80:{46,46}]
  wire  _GEN_100 = 7'h64 == index ? valid1_100 : _GEN_99; // @[dcache.scala 80:{46,46}]
  wire  _GEN_101 = 7'h65 == index ? valid1_101 : _GEN_100; // @[dcache.scala 80:{46,46}]
  wire  _GEN_102 = 7'h66 == index ? valid1_102 : _GEN_101; // @[dcache.scala 80:{46,46}]
  wire  _GEN_103 = 7'h67 == index ? valid1_103 : _GEN_102; // @[dcache.scala 80:{46,46}]
  wire  _GEN_104 = 7'h68 == index ? valid1_104 : _GEN_103; // @[dcache.scala 80:{46,46}]
  wire  _GEN_105 = 7'h69 == index ? valid1_105 : _GEN_104; // @[dcache.scala 80:{46,46}]
  wire  _GEN_106 = 7'h6a == index ? valid1_106 : _GEN_105; // @[dcache.scala 80:{46,46}]
  wire  _GEN_107 = 7'h6b == index ? valid1_107 : _GEN_106; // @[dcache.scala 80:{46,46}]
  wire  _GEN_108 = 7'h6c == index ? valid1_108 : _GEN_107; // @[dcache.scala 80:{46,46}]
  wire  _GEN_109 = 7'h6d == index ? valid1_109 : _GEN_108; // @[dcache.scala 80:{46,46}]
  wire  _GEN_110 = 7'h6e == index ? valid1_110 : _GEN_109; // @[dcache.scala 80:{46,46}]
  wire  _GEN_111 = 7'h6f == index ? valid1_111 : _GEN_110; // @[dcache.scala 80:{46,46}]
  wire  _GEN_112 = 7'h70 == index ? valid1_112 : _GEN_111; // @[dcache.scala 80:{46,46}]
  wire  _GEN_113 = 7'h71 == index ? valid1_113 : _GEN_112; // @[dcache.scala 80:{46,46}]
  wire  _GEN_114 = 7'h72 == index ? valid1_114 : _GEN_113; // @[dcache.scala 80:{46,46}]
  wire  _GEN_115 = 7'h73 == index ? valid1_115 : _GEN_114; // @[dcache.scala 80:{46,46}]
  wire  _GEN_116 = 7'h74 == index ? valid1_116 : _GEN_115; // @[dcache.scala 80:{46,46}]
  wire  _GEN_117 = 7'h75 == index ? valid1_117 : _GEN_116; // @[dcache.scala 80:{46,46}]
  wire  _GEN_118 = 7'h76 == index ? valid1_118 : _GEN_117; // @[dcache.scala 80:{46,46}]
  wire  _GEN_119 = 7'h77 == index ? valid1_119 : _GEN_118; // @[dcache.scala 80:{46,46}]
  wire  _GEN_120 = 7'h78 == index ? valid1_120 : _GEN_119; // @[dcache.scala 80:{46,46}]
  wire  _GEN_121 = 7'h79 == index ? valid1_121 : _GEN_120; // @[dcache.scala 80:{46,46}]
  wire  _GEN_122 = 7'h7a == index ? valid1_122 : _GEN_121; // @[dcache.scala 80:{46,46}]
  wire  _GEN_123 = 7'h7b == index ? valid1_123 : _GEN_122; // @[dcache.scala 80:{46,46}]
  wire  _GEN_124 = 7'h7c == index ? valid1_124 : _GEN_123; // @[dcache.scala 80:{46,46}]
  wire  _GEN_125 = 7'h7d == index ? valid1_125 : _GEN_124; // @[dcache.scala 80:{46,46}]
  wire  _GEN_126 = 7'h7e == index ? valid1_126 : _GEN_125; // @[dcache.scala 80:{46,46}]
  wire  _GEN_127 = 7'h7f == index ? valid1_127 : _GEN_126; // @[dcache.scala 80:{46,46}]
  wire  _GEN_129 = 7'h1 == index ? valid0_1 : valid0_0; // @[dcache.scala 80:{70,70}]
  wire  _GEN_130 = 7'h2 == index ? valid0_2 : _GEN_129; // @[dcache.scala 80:{70,70}]
  wire  _GEN_131 = 7'h3 == index ? valid0_3 : _GEN_130; // @[dcache.scala 80:{70,70}]
  wire  _GEN_132 = 7'h4 == index ? valid0_4 : _GEN_131; // @[dcache.scala 80:{70,70}]
  wire  _GEN_133 = 7'h5 == index ? valid0_5 : _GEN_132; // @[dcache.scala 80:{70,70}]
  wire  _GEN_134 = 7'h6 == index ? valid0_6 : _GEN_133; // @[dcache.scala 80:{70,70}]
  wire  _GEN_135 = 7'h7 == index ? valid0_7 : _GEN_134; // @[dcache.scala 80:{70,70}]
  wire  _GEN_136 = 7'h8 == index ? valid0_8 : _GEN_135; // @[dcache.scala 80:{70,70}]
  wire  _GEN_137 = 7'h9 == index ? valid0_9 : _GEN_136; // @[dcache.scala 80:{70,70}]
  wire  _GEN_138 = 7'ha == index ? valid0_10 : _GEN_137; // @[dcache.scala 80:{70,70}]
  wire  _GEN_139 = 7'hb == index ? valid0_11 : _GEN_138; // @[dcache.scala 80:{70,70}]
  wire  _GEN_140 = 7'hc == index ? valid0_12 : _GEN_139; // @[dcache.scala 80:{70,70}]
  wire  _GEN_141 = 7'hd == index ? valid0_13 : _GEN_140; // @[dcache.scala 80:{70,70}]
  wire  _GEN_142 = 7'he == index ? valid0_14 : _GEN_141; // @[dcache.scala 80:{70,70}]
  wire  _GEN_143 = 7'hf == index ? valid0_15 : _GEN_142; // @[dcache.scala 80:{70,70}]
  wire  _GEN_144 = 7'h10 == index ? valid0_16 : _GEN_143; // @[dcache.scala 80:{70,70}]
  wire  _GEN_145 = 7'h11 == index ? valid0_17 : _GEN_144; // @[dcache.scala 80:{70,70}]
  wire  _GEN_146 = 7'h12 == index ? valid0_18 : _GEN_145; // @[dcache.scala 80:{70,70}]
  wire  _GEN_147 = 7'h13 == index ? valid0_19 : _GEN_146; // @[dcache.scala 80:{70,70}]
  wire  _GEN_148 = 7'h14 == index ? valid0_20 : _GEN_147; // @[dcache.scala 80:{70,70}]
  wire  _GEN_149 = 7'h15 == index ? valid0_21 : _GEN_148; // @[dcache.scala 80:{70,70}]
  wire  _GEN_150 = 7'h16 == index ? valid0_22 : _GEN_149; // @[dcache.scala 80:{70,70}]
  wire  _GEN_151 = 7'h17 == index ? valid0_23 : _GEN_150; // @[dcache.scala 80:{70,70}]
  wire  _GEN_152 = 7'h18 == index ? valid0_24 : _GEN_151; // @[dcache.scala 80:{70,70}]
  wire  _GEN_153 = 7'h19 == index ? valid0_25 : _GEN_152; // @[dcache.scala 80:{70,70}]
  wire  _GEN_154 = 7'h1a == index ? valid0_26 : _GEN_153; // @[dcache.scala 80:{70,70}]
  wire  _GEN_155 = 7'h1b == index ? valid0_27 : _GEN_154; // @[dcache.scala 80:{70,70}]
  wire  _GEN_156 = 7'h1c == index ? valid0_28 : _GEN_155; // @[dcache.scala 80:{70,70}]
  wire  _GEN_157 = 7'h1d == index ? valid0_29 : _GEN_156; // @[dcache.scala 80:{70,70}]
  wire  _GEN_158 = 7'h1e == index ? valid0_30 : _GEN_157; // @[dcache.scala 80:{70,70}]
  wire  _GEN_159 = 7'h1f == index ? valid0_31 : _GEN_158; // @[dcache.scala 80:{70,70}]
  wire  _GEN_160 = 7'h20 == index ? valid0_32 : _GEN_159; // @[dcache.scala 80:{70,70}]
  wire  _GEN_161 = 7'h21 == index ? valid0_33 : _GEN_160; // @[dcache.scala 80:{70,70}]
  wire  _GEN_162 = 7'h22 == index ? valid0_34 : _GEN_161; // @[dcache.scala 80:{70,70}]
  wire  _GEN_163 = 7'h23 == index ? valid0_35 : _GEN_162; // @[dcache.scala 80:{70,70}]
  wire  _GEN_164 = 7'h24 == index ? valid0_36 : _GEN_163; // @[dcache.scala 80:{70,70}]
  wire  _GEN_165 = 7'h25 == index ? valid0_37 : _GEN_164; // @[dcache.scala 80:{70,70}]
  wire  _GEN_166 = 7'h26 == index ? valid0_38 : _GEN_165; // @[dcache.scala 80:{70,70}]
  wire  _GEN_167 = 7'h27 == index ? valid0_39 : _GEN_166; // @[dcache.scala 80:{70,70}]
  wire  _GEN_168 = 7'h28 == index ? valid0_40 : _GEN_167; // @[dcache.scala 80:{70,70}]
  wire  _GEN_169 = 7'h29 == index ? valid0_41 : _GEN_168; // @[dcache.scala 80:{70,70}]
  wire  _GEN_170 = 7'h2a == index ? valid0_42 : _GEN_169; // @[dcache.scala 80:{70,70}]
  wire  _GEN_171 = 7'h2b == index ? valid0_43 : _GEN_170; // @[dcache.scala 80:{70,70}]
  wire  _GEN_172 = 7'h2c == index ? valid0_44 : _GEN_171; // @[dcache.scala 80:{70,70}]
  wire  _GEN_173 = 7'h2d == index ? valid0_45 : _GEN_172; // @[dcache.scala 80:{70,70}]
  wire  _GEN_174 = 7'h2e == index ? valid0_46 : _GEN_173; // @[dcache.scala 80:{70,70}]
  wire  _GEN_175 = 7'h2f == index ? valid0_47 : _GEN_174; // @[dcache.scala 80:{70,70}]
  wire  _GEN_176 = 7'h30 == index ? valid0_48 : _GEN_175; // @[dcache.scala 80:{70,70}]
  wire  _GEN_177 = 7'h31 == index ? valid0_49 : _GEN_176; // @[dcache.scala 80:{70,70}]
  wire  _GEN_178 = 7'h32 == index ? valid0_50 : _GEN_177; // @[dcache.scala 80:{70,70}]
  wire  _GEN_179 = 7'h33 == index ? valid0_51 : _GEN_178; // @[dcache.scala 80:{70,70}]
  wire  _GEN_180 = 7'h34 == index ? valid0_52 : _GEN_179; // @[dcache.scala 80:{70,70}]
  wire  _GEN_181 = 7'h35 == index ? valid0_53 : _GEN_180; // @[dcache.scala 80:{70,70}]
  wire  _GEN_182 = 7'h36 == index ? valid0_54 : _GEN_181; // @[dcache.scala 80:{70,70}]
  wire  _GEN_183 = 7'h37 == index ? valid0_55 : _GEN_182; // @[dcache.scala 80:{70,70}]
  wire  _GEN_184 = 7'h38 == index ? valid0_56 : _GEN_183; // @[dcache.scala 80:{70,70}]
  wire  _GEN_185 = 7'h39 == index ? valid0_57 : _GEN_184; // @[dcache.scala 80:{70,70}]
  wire  _GEN_186 = 7'h3a == index ? valid0_58 : _GEN_185; // @[dcache.scala 80:{70,70}]
  wire  _GEN_187 = 7'h3b == index ? valid0_59 : _GEN_186; // @[dcache.scala 80:{70,70}]
  wire  _GEN_188 = 7'h3c == index ? valid0_60 : _GEN_187; // @[dcache.scala 80:{70,70}]
  wire  _GEN_189 = 7'h3d == index ? valid0_61 : _GEN_188; // @[dcache.scala 80:{70,70}]
  wire  _GEN_190 = 7'h3e == index ? valid0_62 : _GEN_189; // @[dcache.scala 80:{70,70}]
  wire  _GEN_191 = 7'h3f == index ? valid0_63 : _GEN_190; // @[dcache.scala 80:{70,70}]
  wire  _GEN_192 = 7'h40 == index ? valid0_64 : _GEN_191; // @[dcache.scala 80:{70,70}]
  wire  _GEN_193 = 7'h41 == index ? valid0_65 : _GEN_192; // @[dcache.scala 80:{70,70}]
  wire  _GEN_194 = 7'h42 == index ? valid0_66 : _GEN_193; // @[dcache.scala 80:{70,70}]
  wire  _GEN_195 = 7'h43 == index ? valid0_67 : _GEN_194; // @[dcache.scala 80:{70,70}]
  wire  _GEN_196 = 7'h44 == index ? valid0_68 : _GEN_195; // @[dcache.scala 80:{70,70}]
  wire  _GEN_197 = 7'h45 == index ? valid0_69 : _GEN_196; // @[dcache.scala 80:{70,70}]
  wire  _GEN_198 = 7'h46 == index ? valid0_70 : _GEN_197; // @[dcache.scala 80:{70,70}]
  wire  _GEN_199 = 7'h47 == index ? valid0_71 : _GEN_198; // @[dcache.scala 80:{70,70}]
  wire  _GEN_200 = 7'h48 == index ? valid0_72 : _GEN_199; // @[dcache.scala 80:{70,70}]
  wire  _GEN_201 = 7'h49 == index ? valid0_73 : _GEN_200; // @[dcache.scala 80:{70,70}]
  wire  _GEN_202 = 7'h4a == index ? valid0_74 : _GEN_201; // @[dcache.scala 80:{70,70}]
  wire  _GEN_203 = 7'h4b == index ? valid0_75 : _GEN_202; // @[dcache.scala 80:{70,70}]
  wire  _GEN_204 = 7'h4c == index ? valid0_76 : _GEN_203; // @[dcache.scala 80:{70,70}]
  wire  _GEN_205 = 7'h4d == index ? valid0_77 : _GEN_204; // @[dcache.scala 80:{70,70}]
  wire  _GEN_206 = 7'h4e == index ? valid0_78 : _GEN_205; // @[dcache.scala 80:{70,70}]
  wire  _GEN_207 = 7'h4f == index ? valid0_79 : _GEN_206; // @[dcache.scala 80:{70,70}]
  wire  _GEN_208 = 7'h50 == index ? valid0_80 : _GEN_207; // @[dcache.scala 80:{70,70}]
  wire  _GEN_209 = 7'h51 == index ? valid0_81 : _GEN_208; // @[dcache.scala 80:{70,70}]
  wire  _GEN_210 = 7'h52 == index ? valid0_82 : _GEN_209; // @[dcache.scala 80:{70,70}]
  wire  _GEN_211 = 7'h53 == index ? valid0_83 : _GEN_210; // @[dcache.scala 80:{70,70}]
  wire  _GEN_212 = 7'h54 == index ? valid0_84 : _GEN_211; // @[dcache.scala 80:{70,70}]
  wire  _GEN_213 = 7'h55 == index ? valid0_85 : _GEN_212; // @[dcache.scala 80:{70,70}]
  wire  _GEN_214 = 7'h56 == index ? valid0_86 : _GEN_213; // @[dcache.scala 80:{70,70}]
  wire  _GEN_215 = 7'h57 == index ? valid0_87 : _GEN_214; // @[dcache.scala 80:{70,70}]
  wire  _GEN_216 = 7'h58 == index ? valid0_88 : _GEN_215; // @[dcache.scala 80:{70,70}]
  wire  _GEN_217 = 7'h59 == index ? valid0_89 : _GEN_216; // @[dcache.scala 80:{70,70}]
  wire  _GEN_218 = 7'h5a == index ? valid0_90 : _GEN_217; // @[dcache.scala 80:{70,70}]
  wire  _GEN_219 = 7'h5b == index ? valid0_91 : _GEN_218; // @[dcache.scala 80:{70,70}]
  wire  _GEN_220 = 7'h5c == index ? valid0_92 : _GEN_219; // @[dcache.scala 80:{70,70}]
  wire  _GEN_221 = 7'h5d == index ? valid0_93 : _GEN_220; // @[dcache.scala 80:{70,70}]
  wire  _GEN_222 = 7'h5e == index ? valid0_94 : _GEN_221; // @[dcache.scala 80:{70,70}]
  wire  _GEN_223 = 7'h5f == index ? valid0_95 : _GEN_222; // @[dcache.scala 80:{70,70}]
  wire  _GEN_224 = 7'h60 == index ? valid0_96 : _GEN_223; // @[dcache.scala 80:{70,70}]
  wire  _GEN_225 = 7'h61 == index ? valid0_97 : _GEN_224; // @[dcache.scala 80:{70,70}]
  wire  _GEN_226 = 7'h62 == index ? valid0_98 : _GEN_225; // @[dcache.scala 80:{70,70}]
  wire  _GEN_227 = 7'h63 == index ? valid0_99 : _GEN_226; // @[dcache.scala 80:{70,70}]
  wire  _GEN_228 = 7'h64 == index ? valid0_100 : _GEN_227; // @[dcache.scala 80:{70,70}]
  wire  _GEN_229 = 7'h65 == index ? valid0_101 : _GEN_228; // @[dcache.scala 80:{70,70}]
  wire  _GEN_230 = 7'h66 == index ? valid0_102 : _GEN_229; // @[dcache.scala 80:{70,70}]
  wire  _GEN_231 = 7'h67 == index ? valid0_103 : _GEN_230; // @[dcache.scala 80:{70,70}]
  wire  _GEN_232 = 7'h68 == index ? valid0_104 : _GEN_231; // @[dcache.scala 80:{70,70}]
  wire  _GEN_233 = 7'h69 == index ? valid0_105 : _GEN_232; // @[dcache.scala 80:{70,70}]
  wire  _GEN_234 = 7'h6a == index ? valid0_106 : _GEN_233; // @[dcache.scala 80:{70,70}]
  wire  _GEN_235 = 7'h6b == index ? valid0_107 : _GEN_234; // @[dcache.scala 80:{70,70}]
  wire  _GEN_236 = 7'h6c == index ? valid0_108 : _GEN_235; // @[dcache.scala 80:{70,70}]
  wire  _GEN_237 = 7'h6d == index ? valid0_109 : _GEN_236; // @[dcache.scala 80:{70,70}]
  wire  _GEN_238 = 7'h6e == index ? valid0_110 : _GEN_237; // @[dcache.scala 80:{70,70}]
  wire  _GEN_239 = 7'h6f == index ? valid0_111 : _GEN_238; // @[dcache.scala 80:{70,70}]
  wire  _GEN_240 = 7'h70 == index ? valid0_112 : _GEN_239; // @[dcache.scala 80:{70,70}]
  wire  _GEN_241 = 7'h71 == index ? valid0_113 : _GEN_240; // @[dcache.scala 80:{70,70}]
  wire  _GEN_242 = 7'h72 == index ? valid0_114 : _GEN_241; // @[dcache.scala 80:{70,70}]
  wire  _GEN_243 = 7'h73 == index ? valid0_115 : _GEN_242; // @[dcache.scala 80:{70,70}]
  wire  _GEN_244 = 7'h74 == index ? valid0_116 : _GEN_243; // @[dcache.scala 80:{70,70}]
  wire  _GEN_245 = 7'h75 == index ? valid0_117 : _GEN_244; // @[dcache.scala 80:{70,70}]
  wire  _GEN_246 = 7'h76 == index ? valid0_118 : _GEN_245; // @[dcache.scala 80:{70,70}]
  wire  _GEN_247 = 7'h77 == index ? valid0_119 : _GEN_246; // @[dcache.scala 80:{70,70}]
  wire  _GEN_248 = 7'h78 == index ? valid0_120 : _GEN_247; // @[dcache.scala 80:{70,70}]
  wire  _GEN_249 = 7'h79 == index ? valid0_121 : _GEN_248; // @[dcache.scala 80:{70,70}]
  wire  _GEN_250 = 7'h7a == index ? valid0_122 : _GEN_249; // @[dcache.scala 80:{70,70}]
  wire  _GEN_251 = 7'h7b == index ? valid0_123 : _GEN_250; // @[dcache.scala 80:{70,70}]
  wire  _GEN_252 = 7'h7c == index ? valid0_124 : _GEN_251; // @[dcache.scala 80:{70,70}]
  wire  _GEN_253 = 7'h7d == index ? valid0_125 : _GEN_252; // @[dcache.scala 80:{70,70}]
  wire  _GEN_254 = 7'h7e == index ? valid0_126 : _GEN_253; // @[dcache.scala 80:{70,70}]
  wire  _GEN_255 = 7'h7f == index ? valid0_127 : _GEN_254; // @[dcache.scala 80:{70,70}]
  wire  _should_write_back_T_8 = victim ? _GEN_127 : _GEN_255; // @[dcache.scala 80:8]
  wire  _should_write_back_T_9 = state == 2'h2 & io_mem_master_readData_valid & io_mem_master_readData_ready & ~uncache
     & _should_write_back_T_8; // @[dcache.scala 79:115]
  wire  _GEN_257 = 7'h1 == index ? dirty1_1 : dirty1_0; // @[dcache.scala 80:{80,80}]
  wire  _GEN_258 = 7'h2 == index ? dirty1_2 : _GEN_257; // @[dcache.scala 80:{80,80}]
  wire  _GEN_259 = 7'h3 == index ? dirty1_3 : _GEN_258; // @[dcache.scala 80:{80,80}]
  wire  _GEN_260 = 7'h4 == index ? dirty1_4 : _GEN_259; // @[dcache.scala 80:{80,80}]
  wire  _GEN_261 = 7'h5 == index ? dirty1_5 : _GEN_260; // @[dcache.scala 80:{80,80}]
  wire  _GEN_262 = 7'h6 == index ? dirty1_6 : _GEN_261; // @[dcache.scala 80:{80,80}]
  wire  _GEN_263 = 7'h7 == index ? dirty1_7 : _GEN_262; // @[dcache.scala 80:{80,80}]
  wire  _GEN_264 = 7'h8 == index ? dirty1_8 : _GEN_263; // @[dcache.scala 80:{80,80}]
  wire  _GEN_265 = 7'h9 == index ? dirty1_9 : _GEN_264; // @[dcache.scala 80:{80,80}]
  wire  _GEN_266 = 7'ha == index ? dirty1_10 : _GEN_265; // @[dcache.scala 80:{80,80}]
  wire  _GEN_267 = 7'hb == index ? dirty1_11 : _GEN_266; // @[dcache.scala 80:{80,80}]
  wire  _GEN_268 = 7'hc == index ? dirty1_12 : _GEN_267; // @[dcache.scala 80:{80,80}]
  wire  _GEN_269 = 7'hd == index ? dirty1_13 : _GEN_268; // @[dcache.scala 80:{80,80}]
  wire  _GEN_270 = 7'he == index ? dirty1_14 : _GEN_269; // @[dcache.scala 80:{80,80}]
  wire  _GEN_271 = 7'hf == index ? dirty1_15 : _GEN_270; // @[dcache.scala 80:{80,80}]
  wire  _GEN_272 = 7'h10 == index ? dirty1_16 : _GEN_271; // @[dcache.scala 80:{80,80}]
  wire  _GEN_273 = 7'h11 == index ? dirty1_17 : _GEN_272; // @[dcache.scala 80:{80,80}]
  wire  _GEN_274 = 7'h12 == index ? dirty1_18 : _GEN_273; // @[dcache.scala 80:{80,80}]
  wire  _GEN_275 = 7'h13 == index ? dirty1_19 : _GEN_274; // @[dcache.scala 80:{80,80}]
  wire  _GEN_276 = 7'h14 == index ? dirty1_20 : _GEN_275; // @[dcache.scala 80:{80,80}]
  wire  _GEN_277 = 7'h15 == index ? dirty1_21 : _GEN_276; // @[dcache.scala 80:{80,80}]
  wire  _GEN_278 = 7'h16 == index ? dirty1_22 : _GEN_277; // @[dcache.scala 80:{80,80}]
  wire  _GEN_279 = 7'h17 == index ? dirty1_23 : _GEN_278; // @[dcache.scala 80:{80,80}]
  wire  _GEN_280 = 7'h18 == index ? dirty1_24 : _GEN_279; // @[dcache.scala 80:{80,80}]
  wire  _GEN_281 = 7'h19 == index ? dirty1_25 : _GEN_280; // @[dcache.scala 80:{80,80}]
  wire  _GEN_282 = 7'h1a == index ? dirty1_26 : _GEN_281; // @[dcache.scala 80:{80,80}]
  wire  _GEN_283 = 7'h1b == index ? dirty1_27 : _GEN_282; // @[dcache.scala 80:{80,80}]
  wire  _GEN_284 = 7'h1c == index ? dirty1_28 : _GEN_283; // @[dcache.scala 80:{80,80}]
  wire  _GEN_285 = 7'h1d == index ? dirty1_29 : _GEN_284; // @[dcache.scala 80:{80,80}]
  wire  _GEN_286 = 7'h1e == index ? dirty1_30 : _GEN_285; // @[dcache.scala 80:{80,80}]
  wire  _GEN_287 = 7'h1f == index ? dirty1_31 : _GEN_286; // @[dcache.scala 80:{80,80}]
  wire  _GEN_288 = 7'h20 == index ? dirty1_32 : _GEN_287; // @[dcache.scala 80:{80,80}]
  wire  _GEN_289 = 7'h21 == index ? dirty1_33 : _GEN_288; // @[dcache.scala 80:{80,80}]
  wire  _GEN_290 = 7'h22 == index ? dirty1_34 : _GEN_289; // @[dcache.scala 80:{80,80}]
  wire  _GEN_291 = 7'h23 == index ? dirty1_35 : _GEN_290; // @[dcache.scala 80:{80,80}]
  wire  _GEN_292 = 7'h24 == index ? dirty1_36 : _GEN_291; // @[dcache.scala 80:{80,80}]
  wire  _GEN_293 = 7'h25 == index ? dirty1_37 : _GEN_292; // @[dcache.scala 80:{80,80}]
  wire  _GEN_294 = 7'h26 == index ? dirty1_38 : _GEN_293; // @[dcache.scala 80:{80,80}]
  wire  _GEN_295 = 7'h27 == index ? dirty1_39 : _GEN_294; // @[dcache.scala 80:{80,80}]
  wire  _GEN_296 = 7'h28 == index ? dirty1_40 : _GEN_295; // @[dcache.scala 80:{80,80}]
  wire  _GEN_297 = 7'h29 == index ? dirty1_41 : _GEN_296; // @[dcache.scala 80:{80,80}]
  wire  _GEN_298 = 7'h2a == index ? dirty1_42 : _GEN_297; // @[dcache.scala 80:{80,80}]
  wire  _GEN_299 = 7'h2b == index ? dirty1_43 : _GEN_298; // @[dcache.scala 80:{80,80}]
  wire  _GEN_300 = 7'h2c == index ? dirty1_44 : _GEN_299; // @[dcache.scala 80:{80,80}]
  wire  _GEN_301 = 7'h2d == index ? dirty1_45 : _GEN_300; // @[dcache.scala 80:{80,80}]
  wire  _GEN_302 = 7'h2e == index ? dirty1_46 : _GEN_301; // @[dcache.scala 80:{80,80}]
  wire  _GEN_303 = 7'h2f == index ? dirty1_47 : _GEN_302; // @[dcache.scala 80:{80,80}]
  wire  _GEN_304 = 7'h30 == index ? dirty1_48 : _GEN_303; // @[dcache.scala 80:{80,80}]
  wire  _GEN_305 = 7'h31 == index ? dirty1_49 : _GEN_304; // @[dcache.scala 80:{80,80}]
  wire  _GEN_306 = 7'h32 == index ? dirty1_50 : _GEN_305; // @[dcache.scala 80:{80,80}]
  wire  _GEN_307 = 7'h33 == index ? dirty1_51 : _GEN_306; // @[dcache.scala 80:{80,80}]
  wire  _GEN_308 = 7'h34 == index ? dirty1_52 : _GEN_307; // @[dcache.scala 80:{80,80}]
  wire  _GEN_309 = 7'h35 == index ? dirty1_53 : _GEN_308; // @[dcache.scala 80:{80,80}]
  wire  _GEN_310 = 7'h36 == index ? dirty1_54 : _GEN_309; // @[dcache.scala 80:{80,80}]
  wire  _GEN_311 = 7'h37 == index ? dirty1_55 : _GEN_310; // @[dcache.scala 80:{80,80}]
  wire  _GEN_312 = 7'h38 == index ? dirty1_56 : _GEN_311; // @[dcache.scala 80:{80,80}]
  wire  _GEN_313 = 7'h39 == index ? dirty1_57 : _GEN_312; // @[dcache.scala 80:{80,80}]
  wire  _GEN_314 = 7'h3a == index ? dirty1_58 : _GEN_313; // @[dcache.scala 80:{80,80}]
  wire  _GEN_315 = 7'h3b == index ? dirty1_59 : _GEN_314; // @[dcache.scala 80:{80,80}]
  wire  _GEN_316 = 7'h3c == index ? dirty1_60 : _GEN_315; // @[dcache.scala 80:{80,80}]
  wire  _GEN_317 = 7'h3d == index ? dirty1_61 : _GEN_316; // @[dcache.scala 80:{80,80}]
  wire  _GEN_318 = 7'h3e == index ? dirty1_62 : _GEN_317; // @[dcache.scala 80:{80,80}]
  wire  _GEN_319 = 7'h3f == index ? dirty1_63 : _GEN_318; // @[dcache.scala 80:{80,80}]
  wire  _GEN_320 = 7'h40 == index ? dirty1_64 : _GEN_319; // @[dcache.scala 80:{80,80}]
  wire  _GEN_321 = 7'h41 == index ? dirty1_65 : _GEN_320; // @[dcache.scala 80:{80,80}]
  wire  _GEN_322 = 7'h42 == index ? dirty1_66 : _GEN_321; // @[dcache.scala 80:{80,80}]
  wire  _GEN_323 = 7'h43 == index ? dirty1_67 : _GEN_322; // @[dcache.scala 80:{80,80}]
  wire  _GEN_324 = 7'h44 == index ? dirty1_68 : _GEN_323; // @[dcache.scala 80:{80,80}]
  wire  _GEN_325 = 7'h45 == index ? dirty1_69 : _GEN_324; // @[dcache.scala 80:{80,80}]
  wire  _GEN_326 = 7'h46 == index ? dirty1_70 : _GEN_325; // @[dcache.scala 80:{80,80}]
  wire  _GEN_327 = 7'h47 == index ? dirty1_71 : _GEN_326; // @[dcache.scala 80:{80,80}]
  wire  _GEN_328 = 7'h48 == index ? dirty1_72 : _GEN_327; // @[dcache.scala 80:{80,80}]
  wire  _GEN_329 = 7'h49 == index ? dirty1_73 : _GEN_328; // @[dcache.scala 80:{80,80}]
  wire  _GEN_330 = 7'h4a == index ? dirty1_74 : _GEN_329; // @[dcache.scala 80:{80,80}]
  wire  _GEN_331 = 7'h4b == index ? dirty1_75 : _GEN_330; // @[dcache.scala 80:{80,80}]
  wire  _GEN_332 = 7'h4c == index ? dirty1_76 : _GEN_331; // @[dcache.scala 80:{80,80}]
  wire  _GEN_333 = 7'h4d == index ? dirty1_77 : _GEN_332; // @[dcache.scala 80:{80,80}]
  wire  _GEN_334 = 7'h4e == index ? dirty1_78 : _GEN_333; // @[dcache.scala 80:{80,80}]
  wire  _GEN_335 = 7'h4f == index ? dirty1_79 : _GEN_334; // @[dcache.scala 80:{80,80}]
  wire  _GEN_336 = 7'h50 == index ? dirty1_80 : _GEN_335; // @[dcache.scala 80:{80,80}]
  wire  _GEN_337 = 7'h51 == index ? dirty1_81 : _GEN_336; // @[dcache.scala 80:{80,80}]
  wire  _GEN_338 = 7'h52 == index ? dirty1_82 : _GEN_337; // @[dcache.scala 80:{80,80}]
  wire  _GEN_339 = 7'h53 == index ? dirty1_83 : _GEN_338; // @[dcache.scala 80:{80,80}]
  wire  _GEN_340 = 7'h54 == index ? dirty1_84 : _GEN_339; // @[dcache.scala 80:{80,80}]
  wire  _GEN_341 = 7'h55 == index ? dirty1_85 : _GEN_340; // @[dcache.scala 80:{80,80}]
  wire  _GEN_342 = 7'h56 == index ? dirty1_86 : _GEN_341; // @[dcache.scala 80:{80,80}]
  wire  _GEN_343 = 7'h57 == index ? dirty1_87 : _GEN_342; // @[dcache.scala 80:{80,80}]
  wire  _GEN_344 = 7'h58 == index ? dirty1_88 : _GEN_343; // @[dcache.scala 80:{80,80}]
  wire  _GEN_345 = 7'h59 == index ? dirty1_89 : _GEN_344; // @[dcache.scala 80:{80,80}]
  wire  _GEN_346 = 7'h5a == index ? dirty1_90 : _GEN_345; // @[dcache.scala 80:{80,80}]
  wire  _GEN_347 = 7'h5b == index ? dirty1_91 : _GEN_346; // @[dcache.scala 80:{80,80}]
  wire  _GEN_348 = 7'h5c == index ? dirty1_92 : _GEN_347; // @[dcache.scala 80:{80,80}]
  wire  _GEN_349 = 7'h5d == index ? dirty1_93 : _GEN_348; // @[dcache.scala 80:{80,80}]
  wire  _GEN_350 = 7'h5e == index ? dirty1_94 : _GEN_349; // @[dcache.scala 80:{80,80}]
  wire  _GEN_351 = 7'h5f == index ? dirty1_95 : _GEN_350; // @[dcache.scala 80:{80,80}]
  wire  _GEN_352 = 7'h60 == index ? dirty1_96 : _GEN_351; // @[dcache.scala 80:{80,80}]
  wire  _GEN_353 = 7'h61 == index ? dirty1_97 : _GEN_352; // @[dcache.scala 80:{80,80}]
  wire  _GEN_354 = 7'h62 == index ? dirty1_98 : _GEN_353; // @[dcache.scala 80:{80,80}]
  wire  _GEN_355 = 7'h63 == index ? dirty1_99 : _GEN_354; // @[dcache.scala 80:{80,80}]
  wire  _GEN_356 = 7'h64 == index ? dirty1_100 : _GEN_355; // @[dcache.scala 80:{80,80}]
  wire  _GEN_357 = 7'h65 == index ? dirty1_101 : _GEN_356; // @[dcache.scala 80:{80,80}]
  wire  _GEN_358 = 7'h66 == index ? dirty1_102 : _GEN_357; // @[dcache.scala 80:{80,80}]
  wire  _GEN_359 = 7'h67 == index ? dirty1_103 : _GEN_358; // @[dcache.scala 80:{80,80}]
  wire  _GEN_360 = 7'h68 == index ? dirty1_104 : _GEN_359; // @[dcache.scala 80:{80,80}]
  wire  _GEN_361 = 7'h69 == index ? dirty1_105 : _GEN_360; // @[dcache.scala 80:{80,80}]
  wire  _GEN_362 = 7'h6a == index ? dirty1_106 : _GEN_361; // @[dcache.scala 80:{80,80}]
  wire  _GEN_363 = 7'h6b == index ? dirty1_107 : _GEN_362; // @[dcache.scala 80:{80,80}]
  wire  _GEN_364 = 7'h6c == index ? dirty1_108 : _GEN_363; // @[dcache.scala 80:{80,80}]
  wire  _GEN_365 = 7'h6d == index ? dirty1_109 : _GEN_364; // @[dcache.scala 80:{80,80}]
  wire  _GEN_366 = 7'h6e == index ? dirty1_110 : _GEN_365; // @[dcache.scala 80:{80,80}]
  wire  _GEN_367 = 7'h6f == index ? dirty1_111 : _GEN_366; // @[dcache.scala 80:{80,80}]
  wire  _GEN_368 = 7'h70 == index ? dirty1_112 : _GEN_367; // @[dcache.scala 80:{80,80}]
  wire  _GEN_369 = 7'h71 == index ? dirty1_113 : _GEN_368; // @[dcache.scala 80:{80,80}]
  wire  _GEN_370 = 7'h72 == index ? dirty1_114 : _GEN_369; // @[dcache.scala 80:{80,80}]
  wire  _GEN_371 = 7'h73 == index ? dirty1_115 : _GEN_370; // @[dcache.scala 80:{80,80}]
  wire  _GEN_372 = 7'h74 == index ? dirty1_116 : _GEN_371; // @[dcache.scala 80:{80,80}]
  wire  _GEN_373 = 7'h75 == index ? dirty1_117 : _GEN_372; // @[dcache.scala 80:{80,80}]
  wire  _GEN_374 = 7'h76 == index ? dirty1_118 : _GEN_373; // @[dcache.scala 80:{80,80}]
  wire  _GEN_375 = 7'h77 == index ? dirty1_119 : _GEN_374; // @[dcache.scala 80:{80,80}]
  wire  _GEN_376 = 7'h78 == index ? dirty1_120 : _GEN_375; // @[dcache.scala 80:{80,80}]
  wire  _GEN_377 = 7'h79 == index ? dirty1_121 : _GEN_376; // @[dcache.scala 80:{80,80}]
  wire  _GEN_378 = 7'h7a == index ? dirty1_122 : _GEN_377; // @[dcache.scala 80:{80,80}]
  wire  _GEN_379 = 7'h7b == index ? dirty1_123 : _GEN_378; // @[dcache.scala 80:{80,80}]
  wire  _GEN_380 = 7'h7c == index ? dirty1_124 : _GEN_379; // @[dcache.scala 80:{80,80}]
  wire  _GEN_381 = 7'h7d == index ? dirty1_125 : _GEN_380; // @[dcache.scala 80:{80,80}]
  wire  _GEN_382 = 7'h7e == index ? dirty1_126 : _GEN_381; // @[dcache.scala 80:{80,80}]
  wire  _GEN_383 = 7'h7f == index ? dirty1_127 : _GEN_382; // @[dcache.scala 80:{80,80}]
  wire  _GEN_385 = 7'h1 == index ? dirty0_1 : dirty0_0; // @[dcache.scala 80:{80,80}]
  wire  _GEN_386 = 7'h2 == index ? dirty0_2 : _GEN_385; // @[dcache.scala 80:{80,80}]
  wire  _GEN_387 = 7'h3 == index ? dirty0_3 : _GEN_386; // @[dcache.scala 80:{80,80}]
  wire  _GEN_388 = 7'h4 == index ? dirty0_4 : _GEN_387; // @[dcache.scala 80:{80,80}]
  wire  _GEN_389 = 7'h5 == index ? dirty0_5 : _GEN_388; // @[dcache.scala 80:{80,80}]
  wire  _GEN_390 = 7'h6 == index ? dirty0_6 : _GEN_389; // @[dcache.scala 80:{80,80}]
  wire  _GEN_391 = 7'h7 == index ? dirty0_7 : _GEN_390; // @[dcache.scala 80:{80,80}]
  wire  _GEN_392 = 7'h8 == index ? dirty0_8 : _GEN_391; // @[dcache.scala 80:{80,80}]
  wire  _GEN_393 = 7'h9 == index ? dirty0_9 : _GEN_392; // @[dcache.scala 80:{80,80}]
  wire  _GEN_394 = 7'ha == index ? dirty0_10 : _GEN_393; // @[dcache.scala 80:{80,80}]
  wire  _GEN_395 = 7'hb == index ? dirty0_11 : _GEN_394; // @[dcache.scala 80:{80,80}]
  wire  _GEN_396 = 7'hc == index ? dirty0_12 : _GEN_395; // @[dcache.scala 80:{80,80}]
  wire  _GEN_397 = 7'hd == index ? dirty0_13 : _GEN_396; // @[dcache.scala 80:{80,80}]
  wire  _GEN_398 = 7'he == index ? dirty0_14 : _GEN_397; // @[dcache.scala 80:{80,80}]
  wire  _GEN_399 = 7'hf == index ? dirty0_15 : _GEN_398; // @[dcache.scala 80:{80,80}]
  wire  _GEN_400 = 7'h10 == index ? dirty0_16 : _GEN_399; // @[dcache.scala 80:{80,80}]
  wire  _GEN_401 = 7'h11 == index ? dirty0_17 : _GEN_400; // @[dcache.scala 80:{80,80}]
  wire  _GEN_402 = 7'h12 == index ? dirty0_18 : _GEN_401; // @[dcache.scala 80:{80,80}]
  wire  _GEN_403 = 7'h13 == index ? dirty0_19 : _GEN_402; // @[dcache.scala 80:{80,80}]
  wire  _GEN_404 = 7'h14 == index ? dirty0_20 : _GEN_403; // @[dcache.scala 80:{80,80}]
  wire  _GEN_405 = 7'h15 == index ? dirty0_21 : _GEN_404; // @[dcache.scala 80:{80,80}]
  wire  _GEN_406 = 7'h16 == index ? dirty0_22 : _GEN_405; // @[dcache.scala 80:{80,80}]
  wire  _GEN_407 = 7'h17 == index ? dirty0_23 : _GEN_406; // @[dcache.scala 80:{80,80}]
  wire  _GEN_408 = 7'h18 == index ? dirty0_24 : _GEN_407; // @[dcache.scala 80:{80,80}]
  wire  _GEN_409 = 7'h19 == index ? dirty0_25 : _GEN_408; // @[dcache.scala 80:{80,80}]
  wire  _GEN_410 = 7'h1a == index ? dirty0_26 : _GEN_409; // @[dcache.scala 80:{80,80}]
  wire  _GEN_411 = 7'h1b == index ? dirty0_27 : _GEN_410; // @[dcache.scala 80:{80,80}]
  wire  _GEN_412 = 7'h1c == index ? dirty0_28 : _GEN_411; // @[dcache.scala 80:{80,80}]
  wire  _GEN_413 = 7'h1d == index ? dirty0_29 : _GEN_412; // @[dcache.scala 80:{80,80}]
  wire  _GEN_414 = 7'h1e == index ? dirty0_30 : _GEN_413; // @[dcache.scala 80:{80,80}]
  wire  _GEN_415 = 7'h1f == index ? dirty0_31 : _GEN_414; // @[dcache.scala 80:{80,80}]
  wire  _GEN_416 = 7'h20 == index ? dirty0_32 : _GEN_415; // @[dcache.scala 80:{80,80}]
  wire  _GEN_417 = 7'h21 == index ? dirty0_33 : _GEN_416; // @[dcache.scala 80:{80,80}]
  wire  _GEN_418 = 7'h22 == index ? dirty0_34 : _GEN_417; // @[dcache.scala 80:{80,80}]
  wire  _GEN_419 = 7'h23 == index ? dirty0_35 : _GEN_418; // @[dcache.scala 80:{80,80}]
  wire  _GEN_420 = 7'h24 == index ? dirty0_36 : _GEN_419; // @[dcache.scala 80:{80,80}]
  wire  _GEN_421 = 7'h25 == index ? dirty0_37 : _GEN_420; // @[dcache.scala 80:{80,80}]
  wire  _GEN_422 = 7'h26 == index ? dirty0_38 : _GEN_421; // @[dcache.scala 80:{80,80}]
  wire  _GEN_423 = 7'h27 == index ? dirty0_39 : _GEN_422; // @[dcache.scala 80:{80,80}]
  wire  _GEN_424 = 7'h28 == index ? dirty0_40 : _GEN_423; // @[dcache.scala 80:{80,80}]
  wire  _GEN_425 = 7'h29 == index ? dirty0_41 : _GEN_424; // @[dcache.scala 80:{80,80}]
  wire  _GEN_426 = 7'h2a == index ? dirty0_42 : _GEN_425; // @[dcache.scala 80:{80,80}]
  wire  _GEN_427 = 7'h2b == index ? dirty0_43 : _GEN_426; // @[dcache.scala 80:{80,80}]
  wire  _GEN_428 = 7'h2c == index ? dirty0_44 : _GEN_427; // @[dcache.scala 80:{80,80}]
  wire  _GEN_429 = 7'h2d == index ? dirty0_45 : _GEN_428; // @[dcache.scala 80:{80,80}]
  wire  _GEN_430 = 7'h2e == index ? dirty0_46 : _GEN_429; // @[dcache.scala 80:{80,80}]
  wire  _GEN_431 = 7'h2f == index ? dirty0_47 : _GEN_430; // @[dcache.scala 80:{80,80}]
  wire  _GEN_432 = 7'h30 == index ? dirty0_48 : _GEN_431; // @[dcache.scala 80:{80,80}]
  wire  _GEN_433 = 7'h31 == index ? dirty0_49 : _GEN_432; // @[dcache.scala 80:{80,80}]
  wire  _GEN_434 = 7'h32 == index ? dirty0_50 : _GEN_433; // @[dcache.scala 80:{80,80}]
  wire  _GEN_435 = 7'h33 == index ? dirty0_51 : _GEN_434; // @[dcache.scala 80:{80,80}]
  wire  _GEN_436 = 7'h34 == index ? dirty0_52 : _GEN_435; // @[dcache.scala 80:{80,80}]
  wire  _GEN_437 = 7'h35 == index ? dirty0_53 : _GEN_436; // @[dcache.scala 80:{80,80}]
  wire  _GEN_438 = 7'h36 == index ? dirty0_54 : _GEN_437; // @[dcache.scala 80:{80,80}]
  wire  _GEN_439 = 7'h37 == index ? dirty0_55 : _GEN_438; // @[dcache.scala 80:{80,80}]
  wire  _GEN_440 = 7'h38 == index ? dirty0_56 : _GEN_439; // @[dcache.scala 80:{80,80}]
  wire  _GEN_441 = 7'h39 == index ? dirty0_57 : _GEN_440; // @[dcache.scala 80:{80,80}]
  wire  _GEN_442 = 7'h3a == index ? dirty0_58 : _GEN_441; // @[dcache.scala 80:{80,80}]
  wire  _GEN_443 = 7'h3b == index ? dirty0_59 : _GEN_442; // @[dcache.scala 80:{80,80}]
  wire  _GEN_444 = 7'h3c == index ? dirty0_60 : _GEN_443; // @[dcache.scala 80:{80,80}]
  wire  _GEN_445 = 7'h3d == index ? dirty0_61 : _GEN_444; // @[dcache.scala 80:{80,80}]
  wire  _GEN_446 = 7'h3e == index ? dirty0_62 : _GEN_445; // @[dcache.scala 80:{80,80}]
  wire  _GEN_447 = 7'h3f == index ? dirty0_63 : _GEN_446; // @[dcache.scala 80:{80,80}]
  wire  _GEN_448 = 7'h40 == index ? dirty0_64 : _GEN_447; // @[dcache.scala 80:{80,80}]
  wire  _GEN_449 = 7'h41 == index ? dirty0_65 : _GEN_448; // @[dcache.scala 80:{80,80}]
  wire  _GEN_450 = 7'h42 == index ? dirty0_66 : _GEN_449; // @[dcache.scala 80:{80,80}]
  wire  _GEN_451 = 7'h43 == index ? dirty0_67 : _GEN_450; // @[dcache.scala 80:{80,80}]
  wire  _GEN_452 = 7'h44 == index ? dirty0_68 : _GEN_451; // @[dcache.scala 80:{80,80}]
  wire  _GEN_453 = 7'h45 == index ? dirty0_69 : _GEN_452; // @[dcache.scala 80:{80,80}]
  wire  _GEN_454 = 7'h46 == index ? dirty0_70 : _GEN_453; // @[dcache.scala 80:{80,80}]
  wire  _GEN_455 = 7'h47 == index ? dirty0_71 : _GEN_454; // @[dcache.scala 80:{80,80}]
  wire  _GEN_456 = 7'h48 == index ? dirty0_72 : _GEN_455; // @[dcache.scala 80:{80,80}]
  wire  _GEN_457 = 7'h49 == index ? dirty0_73 : _GEN_456; // @[dcache.scala 80:{80,80}]
  wire  _GEN_458 = 7'h4a == index ? dirty0_74 : _GEN_457; // @[dcache.scala 80:{80,80}]
  wire  _GEN_459 = 7'h4b == index ? dirty0_75 : _GEN_458; // @[dcache.scala 80:{80,80}]
  wire  _GEN_460 = 7'h4c == index ? dirty0_76 : _GEN_459; // @[dcache.scala 80:{80,80}]
  wire  _GEN_461 = 7'h4d == index ? dirty0_77 : _GEN_460; // @[dcache.scala 80:{80,80}]
  wire  _GEN_462 = 7'h4e == index ? dirty0_78 : _GEN_461; // @[dcache.scala 80:{80,80}]
  wire  _GEN_463 = 7'h4f == index ? dirty0_79 : _GEN_462; // @[dcache.scala 80:{80,80}]
  wire  _GEN_464 = 7'h50 == index ? dirty0_80 : _GEN_463; // @[dcache.scala 80:{80,80}]
  wire  _GEN_465 = 7'h51 == index ? dirty0_81 : _GEN_464; // @[dcache.scala 80:{80,80}]
  wire  _GEN_466 = 7'h52 == index ? dirty0_82 : _GEN_465; // @[dcache.scala 80:{80,80}]
  wire  _GEN_467 = 7'h53 == index ? dirty0_83 : _GEN_466; // @[dcache.scala 80:{80,80}]
  wire  _GEN_468 = 7'h54 == index ? dirty0_84 : _GEN_467; // @[dcache.scala 80:{80,80}]
  wire  _GEN_469 = 7'h55 == index ? dirty0_85 : _GEN_468; // @[dcache.scala 80:{80,80}]
  wire  _GEN_470 = 7'h56 == index ? dirty0_86 : _GEN_469; // @[dcache.scala 80:{80,80}]
  wire  _GEN_471 = 7'h57 == index ? dirty0_87 : _GEN_470; // @[dcache.scala 80:{80,80}]
  wire  _GEN_472 = 7'h58 == index ? dirty0_88 : _GEN_471; // @[dcache.scala 80:{80,80}]
  wire  _GEN_473 = 7'h59 == index ? dirty0_89 : _GEN_472; // @[dcache.scala 80:{80,80}]
  wire  _GEN_474 = 7'h5a == index ? dirty0_90 : _GEN_473; // @[dcache.scala 80:{80,80}]
  wire  _GEN_475 = 7'h5b == index ? dirty0_91 : _GEN_474; // @[dcache.scala 80:{80,80}]
  wire  _GEN_476 = 7'h5c == index ? dirty0_92 : _GEN_475; // @[dcache.scala 80:{80,80}]
  wire  _GEN_477 = 7'h5d == index ? dirty0_93 : _GEN_476; // @[dcache.scala 80:{80,80}]
  wire  _GEN_478 = 7'h5e == index ? dirty0_94 : _GEN_477; // @[dcache.scala 80:{80,80}]
  wire  _GEN_479 = 7'h5f == index ? dirty0_95 : _GEN_478; // @[dcache.scala 80:{80,80}]
  wire  _GEN_480 = 7'h60 == index ? dirty0_96 : _GEN_479; // @[dcache.scala 80:{80,80}]
  wire  _GEN_481 = 7'h61 == index ? dirty0_97 : _GEN_480; // @[dcache.scala 80:{80,80}]
  wire  _GEN_482 = 7'h62 == index ? dirty0_98 : _GEN_481; // @[dcache.scala 80:{80,80}]
  wire  _GEN_483 = 7'h63 == index ? dirty0_99 : _GEN_482; // @[dcache.scala 80:{80,80}]
  wire  _GEN_484 = 7'h64 == index ? dirty0_100 : _GEN_483; // @[dcache.scala 80:{80,80}]
  wire  _GEN_485 = 7'h65 == index ? dirty0_101 : _GEN_484; // @[dcache.scala 80:{80,80}]
  wire  _GEN_486 = 7'h66 == index ? dirty0_102 : _GEN_485; // @[dcache.scala 80:{80,80}]
  wire  _GEN_487 = 7'h67 == index ? dirty0_103 : _GEN_486; // @[dcache.scala 80:{80,80}]
  wire  _GEN_488 = 7'h68 == index ? dirty0_104 : _GEN_487; // @[dcache.scala 80:{80,80}]
  wire  _GEN_489 = 7'h69 == index ? dirty0_105 : _GEN_488; // @[dcache.scala 80:{80,80}]
  wire  _GEN_490 = 7'h6a == index ? dirty0_106 : _GEN_489; // @[dcache.scala 80:{80,80}]
  wire  _GEN_491 = 7'h6b == index ? dirty0_107 : _GEN_490; // @[dcache.scala 80:{80,80}]
  wire  _GEN_492 = 7'h6c == index ? dirty0_108 : _GEN_491; // @[dcache.scala 80:{80,80}]
  wire  _GEN_493 = 7'h6d == index ? dirty0_109 : _GEN_492; // @[dcache.scala 80:{80,80}]
  wire  _GEN_494 = 7'h6e == index ? dirty0_110 : _GEN_493; // @[dcache.scala 80:{80,80}]
  wire  _GEN_495 = 7'h6f == index ? dirty0_111 : _GEN_494; // @[dcache.scala 80:{80,80}]
  wire  _GEN_496 = 7'h70 == index ? dirty0_112 : _GEN_495; // @[dcache.scala 80:{80,80}]
  wire  _GEN_497 = 7'h71 == index ? dirty0_113 : _GEN_496; // @[dcache.scala 80:{80,80}]
  wire  _GEN_498 = 7'h72 == index ? dirty0_114 : _GEN_497; // @[dcache.scala 80:{80,80}]
  wire  _GEN_499 = 7'h73 == index ? dirty0_115 : _GEN_498; // @[dcache.scala 80:{80,80}]
  wire  _GEN_500 = 7'h74 == index ? dirty0_116 : _GEN_499; // @[dcache.scala 80:{80,80}]
  wire  _GEN_501 = 7'h75 == index ? dirty0_117 : _GEN_500; // @[dcache.scala 80:{80,80}]
  wire  _GEN_502 = 7'h76 == index ? dirty0_118 : _GEN_501; // @[dcache.scala 80:{80,80}]
  wire  _GEN_503 = 7'h77 == index ? dirty0_119 : _GEN_502; // @[dcache.scala 80:{80,80}]
  wire  _GEN_504 = 7'h78 == index ? dirty0_120 : _GEN_503; // @[dcache.scala 80:{80,80}]
  wire  _GEN_505 = 7'h79 == index ? dirty0_121 : _GEN_504; // @[dcache.scala 80:{80,80}]
  wire  _GEN_506 = 7'h7a == index ? dirty0_122 : _GEN_505; // @[dcache.scala 80:{80,80}]
  wire  _GEN_507 = 7'h7b == index ? dirty0_123 : _GEN_506; // @[dcache.scala 80:{80,80}]
  wire  _GEN_508 = 7'h7c == index ? dirty0_124 : _GEN_507; // @[dcache.scala 80:{80,80}]
  wire  _GEN_509 = 7'h7d == index ? dirty0_125 : _GEN_508; // @[dcache.scala 80:{80,80}]
  wire  _GEN_510 = 7'h7e == index ? dirty0_126 : _GEN_509; // @[dcache.scala 80:{80,80}]
  wire  _GEN_511 = 7'h7f == index ? dirty0_127 : _GEN_510; // @[dcache.scala 80:{80,80}]
  wire  _should_write_back_T_11 = victim ? _GEN_383 : _GEN_511; // @[dcache.scala 80:80]
  wire  should_write_back = _should_write_back_T_9 & _should_write_back_T_11; // @[dcache.scala 80:74]
  wire  _write_back_is_finishing_T = ~cpu_mem_Mwout; // @[dcache.scala 86:42]
  wire  write_back_is_finishing = write_done & ~cpu_mem_Mwout & cpu_mem_Men; // @[dcache.scala 86:57]
  wire  _next_state_T = state == 2'h0; // @[dcache.scala 186:12]
  wire  _next_state_T_1 = state == 2'h1; // @[dcache.scala 188:12]
  wire [52:0] _GEN_520 = 7'h1 == index ? tags0_1 : tags0_0; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_521 = 7'h2 == index ? tags0_2 : _GEN_520; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_522 = 7'h3 == index ? tags0_3 : _GEN_521; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_523 = 7'h4 == index ? tags0_4 : _GEN_522; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_524 = 7'h5 == index ? tags0_5 : _GEN_523; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_525 = 7'h6 == index ? tags0_6 : _GEN_524; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_526 = 7'h7 == index ? tags0_7 : _GEN_525; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_527 = 7'h8 == index ? tags0_8 : _GEN_526; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_528 = 7'h9 == index ? tags0_9 : _GEN_527; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_529 = 7'ha == index ? tags0_10 : _GEN_528; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_530 = 7'hb == index ? tags0_11 : _GEN_529; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_531 = 7'hc == index ? tags0_12 : _GEN_530; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_532 = 7'hd == index ? tags0_13 : _GEN_531; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_533 = 7'he == index ? tags0_14 : _GEN_532; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_534 = 7'hf == index ? tags0_15 : _GEN_533; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_535 = 7'h10 == index ? tags0_16 : _GEN_534; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_536 = 7'h11 == index ? tags0_17 : _GEN_535; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_537 = 7'h12 == index ? tags0_18 : _GEN_536; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_538 = 7'h13 == index ? tags0_19 : _GEN_537; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_539 = 7'h14 == index ? tags0_20 : _GEN_538; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_540 = 7'h15 == index ? tags0_21 : _GEN_539; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_541 = 7'h16 == index ? tags0_22 : _GEN_540; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_542 = 7'h17 == index ? tags0_23 : _GEN_541; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_543 = 7'h18 == index ? tags0_24 : _GEN_542; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_544 = 7'h19 == index ? tags0_25 : _GEN_543; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_545 = 7'h1a == index ? tags0_26 : _GEN_544; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_546 = 7'h1b == index ? tags0_27 : _GEN_545; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_547 = 7'h1c == index ? tags0_28 : _GEN_546; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_548 = 7'h1d == index ? tags0_29 : _GEN_547; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_549 = 7'h1e == index ? tags0_30 : _GEN_548; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_550 = 7'h1f == index ? tags0_31 : _GEN_549; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_551 = 7'h20 == index ? tags0_32 : _GEN_550; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_552 = 7'h21 == index ? tags0_33 : _GEN_551; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_553 = 7'h22 == index ? tags0_34 : _GEN_552; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_554 = 7'h23 == index ? tags0_35 : _GEN_553; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_555 = 7'h24 == index ? tags0_36 : _GEN_554; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_556 = 7'h25 == index ? tags0_37 : _GEN_555; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_557 = 7'h26 == index ? tags0_38 : _GEN_556; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_558 = 7'h27 == index ? tags0_39 : _GEN_557; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_559 = 7'h28 == index ? tags0_40 : _GEN_558; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_560 = 7'h29 == index ? tags0_41 : _GEN_559; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_561 = 7'h2a == index ? tags0_42 : _GEN_560; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_562 = 7'h2b == index ? tags0_43 : _GEN_561; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_563 = 7'h2c == index ? tags0_44 : _GEN_562; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_564 = 7'h2d == index ? tags0_45 : _GEN_563; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_565 = 7'h2e == index ? tags0_46 : _GEN_564; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_566 = 7'h2f == index ? tags0_47 : _GEN_565; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_567 = 7'h30 == index ? tags0_48 : _GEN_566; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_568 = 7'h31 == index ? tags0_49 : _GEN_567; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_569 = 7'h32 == index ? tags0_50 : _GEN_568; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_570 = 7'h33 == index ? tags0_51 : _GEN_569; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_571 = 7'h34 == index ? tags0_52 : _GEN_570; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_572 = 7'h35 == index ? tags0_53 : _GEN_571; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_573 = 7'h36 == index ? tags0_54 : _GEN_572; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_574 = 7'h37 == index ? tags0_55 : _GEN_573; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_575 = 7'h38 == index ? tags0_56 : _GEN_574; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_576 = 7'h39 == index ? tags0_57 : _GEN_575; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_577 = 7'h3a == index ? tags0_58 : _GEN_576; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_578 = 7'h3b == index ? tags0_59 : _GEN_577; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_579 = 7'h3c == index ? tags0_60 : _GEN_578; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_580 = 7'h3d == index ? tags0_61 : _GEN_579; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_581 = 7'h3e == index ? tags0_62 : _GEN_580; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_582 = 7'h3f == index ? tags0_63 : _GEN_581; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_583 = 7'h40 == index ? tags0_64 : _GEN_582; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_584 = 7'h41 == index ? tags0_65 : _GEN_583; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_585 = 7'h42 == index ? tags0_66 : _GEN_584; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_586 = 7'h43 == index ? tags0_67 : _GEN_585; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_587 = 7'h44 == index ? tags0_68 : _GEN_586; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_588 = 7'h45 == index ? tags0_69 : _GEN_587; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_589 = 7'h46 == index ? tags0_70 : _GEN_588; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_590 = 7'h47 == index ? tags0_71 : _GEN_589; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_591 = 7'h48 == index ? tags0_72 : _GEN_590; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_592 = 7'h49 == index ? tags0_73 : _GEN_591; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_593 = 7'h4a == index ? tags0_74 : _GEN_592; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_594 = 7'h4b == index ? tags0_75 : _GEN_593; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_595 = 7'h4c == index ? tags0_76 : _GEN_594; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_596 = 7'h4d == index ? tags0_77 : _GEN_595; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_597 = 7'h4e == index ? tags0_78 : _GEN_596; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_598 = 7'h4f == index ? tags0_79 : _GEN_597; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_599 = 7'h50 == index ? tags0_80 : _GEN_598; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_600 = 7'h51 == index ? tags0_81 : _GEN_599; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_601 = 7'h52 == index ? tags0_82 : _GEN_600; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_602 = 7'h53 == index ? tags0_83 : _GEN_601; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_603 = 7'h54 == index ? tags0_84 : _GEN_602; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_604 = 7'h55 == index ? tags0_85 : _GEN_603; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_605 = 7'h56 == index ? tags0_86 : _GEN_604; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_606 = 7'h57 == index ? tags0_87 : _GEN_605; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_607 = 7'h58 == index ? tags0_88 : _GEN_606; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_608 = 7'h59 == index ? tags0_89 : _GEN_607; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_609 = 7'h5a == index ? tags0_90 : _GEN_608; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_610 = 7'h5b == index ? tags0_91 : _GEN_609; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_611 = 7'h5c == index ? tags0_92 : _GEN_610; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_612 = 7'h5d == index ? tags0_93 : _GEN_611; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_613 = 7'h5e == index ? tags0_94 : _GEN_612; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_614 = 7'h5f == index ? tags0_95 : _GEN_613; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_615 = 7'h60 == index ? tags0_96 : _GEN_614; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_616 = 7'h61 == index ? tags0_97 : _GEN_615; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_617 = 7'h62 == index ? tags0_98 : _GEN_616; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_618 = 7'h63 == index ? tags0_99 : _GEN_617; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_619 = 7'h64 == index ? tags0_100 : _GEN_618; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_620 = 7'h65 == index ? tags0_101 : _GEN_619; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_621 = 7'h66 == index ? tags0_102 : _GEN_620; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_622 = 7'h67 == index ? tags0_103 : _GEN_621; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_623 = 7'h68 == index ? tags0_104 : _GEN_622; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_624 = 7'h69 == index ? tags0_105 : _GEN_623; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_625 = 7'h6a == index ? tags0_106 : _GEN_624; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_626 = 7'h6b == index ? tags0_107 : _GEN_625; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_627 = 7'h6c == index ? tags0_108 : _GEN_626; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_628 = 7'h6d == index ? tags0_109 : _GEN_627; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_629 = 7'h6e == index ? tags0_110 : _GEN_628; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_630 = 7'h6f == index ? tags0_111 : _GEN_629; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_631 = 7'h70 == index ? tags0_112 : _GEN_630; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_632 = 7'h71 == index ? tags0_113 : _GEN_631; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_633 = 7'h72 == index ? tags0_114 : _GEN_632; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_634 = 7'h73 == index ? tags0_115 : _GEN_633; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_635 = 7'h74 == index ? tags0_116 : _GEN_634; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_636 = 7'h75 == index ? tags0_117 : _GEN_635; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_637 = 7'h76 == index ? tags0_118 : _GEN_636; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_638 = 7'h77 == index ? tags0_119 : _GEN_637; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_639 = 7'h78 == index ? tags0_120 : _GEN_638; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_640 = 7'h79 == index ? tags0_121 : _GEN_639; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_641 = 7'h7a == index ? tags0_122 : _GEN_640; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_642 = 7'h7b == index ? tags0_123 : _GEN_641; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_643 = 7'h7c == index ? tags0_124 : _GEN_642; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_644 = 7'h7d == index ? tags0_125 : _GEN_643; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_645 = 7'h7e == index ? tags0_126 : _GEN_644; // @[dcache.scala 117:{48,48}]
  wire [52:0] _GEN_646 = 7'h7f == index ? tags0_127 : _GEN_645; // @[dcache.scala 117:{48,48}]
  wire [52:0] tag = cpu_mem_Maddr[63:11]; // @[dcache.scala 114:21]
  wire  hit_bank_0 = _GEN_255 & _GEN_646 == tag & _should_write_back_T_3; // @[dcache.scala 117:67]
  wire [52:0] _GEN_648 = 7'h1 == index ? tags1_1 : tags1_0; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_649 = 7'h2 == index ? tags1_2 : _GEN_648; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_650 = 7'h3 == index ? tags1_3 : _GEN_649; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_651 = 7'h4 == index ? tags1_4 : _GEN_650; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_652 = 7'h5 == index ? tags1_5 : _GEN_651; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_653 = 7'h6 == index ? tags1_6 : _GEN_652; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_654 = 7'h7 == index ? tags1_7 : _GEN_653; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_655 = 7'h8 == index ? tags1_8 : _GEN_654; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_656 = 7'h9 == index ? tags1_9 : _GEN_655; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_657 = 7'ha == index ? tags1_10 : _GEN_656; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_658 = 7'hb == index ? tags1_11 : _GEN_657; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_659 = 7'hc == index ? tags1_12 : _GEN_658; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_660 = 7'hd == index ? tags1_13 : _GEN_659; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_661 = 7'he == index ? tags1_14 : _GEN_660; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_662 = 7'hf == index ? tags1_15 : _GEN_661; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_663 = 7'h10 == index ? tags1_16 : _GEN_662; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_664 = 7'h11 == index ? tags1_17 : _GEN_663; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_665 = 7'h12 == index ? tags1_18 : _GEN_664; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_666 = 7'h13 == index ? tags1_19 : _GEN_665; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_667 = 7'h14 == index ? tags1_20 : _GEN_666; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_668 = 7'h15 == index ? tags1_21 : _GEN_667; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_669 = 7'h16 == index ? tags1_22 : _GEN_668; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_670 = 7'h17 == index ? tags1_23 : _GEN_669; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_671 = 7'h18 == index ? tags1_24 : _GEN_670; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_672 = 7'h19 == index ? tags1_25 : _GEN_671; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_673 = 7'h1a == index ? tags1_26 : _GEN_672; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_674 = 7'h1b == index ? tags1_27 : _GEN_673; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_675 = 7'h1c == index ? tags1_28 : _GEN_674; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_676 = 7'h1d == index ? tags1_29 : _GEN_675; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_677 = 7'h1e == index ? tags1_30 : _GEN_676; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_678 = 7'h1f == index ? tags1_31 : _GEN_677; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_679 = 7'h20 == index ? tags1_32 : _GEN_678; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_680 = 7'h21 == index ? tags1_33 : _GEN_679; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_681 = 7'h22 == index ? tags1_34 : _GEN_680; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_682 = 7'h23 == index ? tags1_35 : _GEN_681; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_683 = 7'h24 == index ? tags1_36 : _GEN_682; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_684 = 7'h25 == index ? tags1_37 : _GEN_683; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_685 = 7'h26 == index ? tags1_38 : _GEN_684; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_686 = 7'h27 == index ? tags1_39 : _GEN_685; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_687 = 7'h28 == index ? tags1_40 : _GEN_686; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_688 = 7'h29 == index ? tags1_41 : _GEN_687; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_689 = 7'h2a == index ? tags1_42 : _GEN_688; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_690 = 7'h2b == index ? tags1_43 : _GEN_689; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_691 = 7'h2c == index ? tags1_44 : _GEN_690; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_692 = 7'h2d == index ? tags1_45 : _GEN_691; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_693 = 7'h2e == index ? tags1_46 : _GEN_692; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_694 = 7'h2f == index ? tags1_47 : _GEN_693; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_695 = 7'h30 == index ? tags1_48 : _GEN_694; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_696 = 7'h31 == index ? tags1_49 : _GEN_695; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_697 = 7'h32 == index ? tags1_50 : _GEN_696; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_698 = 7'h33 == index ? tags1_51 : _GEN_697; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_699 = 7'h34 == index ? tags1_52 : _GEN_698; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_700 = 7'h35 == index ? tags1_53 : _GEN_699; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_701 = 7'h36 == index ? tags1_54 : _GEN_700; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_702 = 7'h37 == index ? tags1_55 : _GEN_701; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_703 = 7'h38 == index ? tags1_56 : _GEN_702; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_704 = 7'h39 == index ? tags1_57 : _GEN_703; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_705 = 7'h3a == index ? tags1_58 : _GEN_704; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_706 = 7'h3b == index ? tags1_59 : _GEN_705; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_707 = 7'h3c == index ? tags1_60 : _GEN_706; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_708 = 7'h3d == index ? tags1_61 : _GEN_707; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_709 = 7'h3e == index ? tags1_62 : _GEN_708; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_710 = 7'h3f == index ? tags1_63 : _GEN_709; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_711 = 7'h40 == index ? tags1_64 : _GEN_710; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_712 = 7'h41 == index ? tags1_65 : _GEN_711; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_713 = 7'h42 == index ? tags1_66 : _GEN_712; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_714 = 7'h43 == index ? tags1_67 : _GEN_713; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_715 = 7'h44 == index ? tags1_68 : _GEN_714; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_716 = 7'h45 == index ? tags1_69 : _GEN_715; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_717 = 7'h46 == index ? tags1_70 : _GEN_716; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_718 = 7'h47 == index ? tags1_71 : _GEN_717; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_719 = 7'h48 == index ? tags1_72 : _GEN_718; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_720 = 7'h49 == index ? tags1_73 : _GEN_719; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_721 = 7'h4a == index ? tags1_74 : _GEN_720; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_722 = 7'h4b == index ? tags1_75 : _GEN_721; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_723 = 7'h4c == index ? tags1_76 : _GEN_722; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_724 = 7'h4d == index ? tags1_77 : _GEN_723; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_725 = 7'h4e == index ? tags1_78 : _GEN_724; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_726 = 7'h4f == index ? tags1_79 : _GEN_725; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_727 = 7'h50 == index ? tags1_80 : _GEN_726; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_728 = 7'h51 == index ? tags1_81 : _GEN_727; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_729 = 7'h52 == index ? tags1_82 : _GEN_728; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_730 = 7'h53 == index ? tags1_83 : _GEN_729; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_731 = 7'h54 == index ? tags1_84 : _GEN_730; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_732 = 7'h55 == index ? tags1_85 : _GEN_731; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_733 = 7'h56 == index ? tags1_86 : _GEN_732; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_734 = 7'h57 == index ? tags1_87 : _GEN_733; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_735 = 7'h58 == index ? tags1_88 : _GEN_734; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_736 = 7'h59 == index ? tags1_89 : _GEN_735; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_737 = 7'h5a == index ? tags1_90 : _GEN_736; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_738 = 7'h5b == index ? tags1_91 : _GEN_737; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_739 = 7'h5c == index ? tags1_92 : _GEN_738; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_740 = 7'h5d == index ? tags1_93 : _GEN_739; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_741 = 7'h5e == index ? tags1_94 : _GEN_740; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_742 = 7'h5f == index ? tags1_95 : _GEN_741; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_743 = 7'h60 == index ? tags1_96 : _GEN_742; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_744 = 7'h61 == index ? tags1_97 : _GEN_743; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_745 = 7'h62 == index ? tags1_98 : _GEN_744; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_746 = 7'h63 == index ? tags1_99 : _GEN_745; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_747 = 7'h64 == index ? tags1_100 : _GEN_746; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_748 = 7'h65 == index ? tags1_101 : _GEN_747; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_749 = 7'h66 == index ? tags1_102 : _GEN_748; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_750 = 7'h67 == index ? tags1_103 : _GEN_749; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_751 = 7'h68 == index ? tags1_104 : _GEN_750; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_752 = 7'h69 == index ? tags1_105 : _GEN_751; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_753 = 7'h6a == index ? tags1_106 : _GEN_752; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_754 = 7'h6b == index ? tags1_107 : _GEN_753; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_755 = 7'h6c == index ? tags1_108 : _GEN_754; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_756 = 7'h6d == index ? tags1_109 : _GEN_755; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_757 = 7'h6e == index ? tags1_110 : _GEN_756; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_758 = 7'h6f == index ? tags1_111 : _GEN_757; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_759 = 7'h70 == index ? tags1_112 : _GEN_758; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_760 = 7'h71 == index ? tags1_113 : _GEN_759; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_761 = 7'h72 == index ? tags1_114 : _GEN_760; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_762 = 7'h73 == index ? tags1_115 : _GEN_761; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_763 = 7'h74 == index ? tags1_116 : _GEN_762; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_764 = 7'h75 == index ? tags1_117 : _GEN_763; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_765 = 7'h76 == index ? tags1_118 : _GEN_764; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_766 = 7'h77 == index ? tags1_119 : _GEN_765; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_767 = 7'h78 == index ? tags1_120 : _GEN_766; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_768 = 7'h79 == index ? tags1_121 : _GEN_767; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_769 = 7'h7a == index ? tags1_122 : _GEN_768; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_770 = 7'h7b == index ? tags1_123 : _GEN_769; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_771 = 7'h7c == index ? tags1_124 : _GEN_770; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_772 = 7'h7d == index ? tags1_125 : _GEN_771; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_773 = 7'h7e == index ? tags1_126 : _GEN_772; // @[dcache.scala 118:{48,48}]
  wire [52:0] _GEN_774 = 7'h7f == index ? tags1_127 : _GEN_773; // @[dcache.scala 118:{48,48}]
  wire  hit_bank_1 = _GEN_127 & _GEN_774 == tag & _should_write_back_T_3; // @[dcache.scala 118:67]
  wire  hit = (hit_bank_0 | hit_bank_1) & _should_write_back_T_3; // @[dcache.scala 119:37]
  wire  _next_state_T_2 = ~hit; // @[dcache.scala 188:27]
  wire  _next_state_T_5 = state == 2'h1 & ~hit & cpu_mem_Men & new_req; // @[dcache.scala 188:48]
  wire  _next_state_T_7 = _should_write_back_T & write_done; // @[dcache.scala 189:22]
  wire  _next_state_T_9 = _should_write_back_T & read_done; // @[dcache.scala 190:22]
  wire  _next_state_T_11 = _should_write_back_T & read_done & ~should_write_back; // @[dcache.scala 190:35]
  wire  _next_state_T_14 = _next_state_T_9 & should_write_back; // @[dcache.scala 191:35]
  wire [1:0] _next_state_T_15 = _next_state_T_14 ? 2'h2 : state; // @[Mux.scala 101:16]
  wire [1:0] _next_state_T_16 = _next_state_T_11 ? 2'h1 : _next_state_T_15; // @[Mux.scala 101:16]
  wire [1:0] _next_state_T_17 = _next_state_T_7 ? 2'h1 : _next_state_T_16; // @[Mux.scala 101:16]
  wire [1:0] _next_state_T_18 = _next_state_T_5 ? 2'h2 : _next_state_T_17; // @[Mux.scala 101:16]
  wire [1:0] next_state = _next_state_T ? 2'h1 : _next_state_T_18; // @[Mux.scala 101:16]
  wire  _T = next_state == 2'h1; // @[dcache.scala 88:16]
  wire [127:0] _read_data_T_1 = hit_bank_1 ? data_array_1_io_o_rdata : 128'h0; // @[Mux.scala 101:16]
  wire [127:0] _read_data_T_2 = hit_bank_0 ? data_array_0_io_o_rdata : _read_data_T_1; // @[Mux.scala 101:16]
  wire [127:0] _read_data_T_4 = _should_write_back_T ? io_mem_master_readData_bits_data : 128'h0; // @[Mux.scala 101:16]
  wire [127:0] read_data = _next_state_T_1 ? _read_data_T_2 : _read_data_T_4; // @[Mux.scala 101:16]
  wire [6:0] _io_cpu_mem_MdataIn_T_1 = {cpu_mem_Maddr[3:0], 3'h0}; // @[dcache.scala 100:53]
  wire [127:0] _io_cpu_mem_MdataIn_T_2 = read_data >> _io_cpu_mem_MdataIn_T_1; // @[dcache.scala 100:32]
  wire  _io_cpu_mem_data_valid_T = next_state != 2'h2; // @[dcache.scala 111:38]
  wire  _io_cpu_mem_data_valid_T_6 = write_state == 3'h1; // @[dcache.scala 111:109]
  wire  _victim_T_1 = ~_GEN_255; // @[dcache.scala 121:6]
  wire  _victim_T_5 = _GEN_255 & ~_GEN_127; // @[dcache.scala 122:27]
  wire  _strb_T = cpu_mem_Mlen == 32'h1; // @[dcache.scala 139:19]
  wire  _strb_T_1 = cpu_mem_Mlen == 32'h2; // @[dcache.scala 140:19]
  wire  _strb_T_2 = cpu_mem_Mlen == 32'h3; // @[dcache.scala 141:19]
  wire  _strb_T_3 = cpu_mem_Mlen == 32'h4; // @[dcache.scala 142:19]
  wire  _strb_T_4 = cpu_mem_Mlen == 32'h8; // @[dcache.scala 143:19]
  wire  _strb_T_5 = cpu_mem_Mlen == 32'h10; // @[dcache.scala 144:19]
  wire [15:0] _strb_T_6 = _strb_T_5 ? 16'hffff : 16'h0; // @[Mux.scala 101:16]
  wire [15:0] _strb_T_7 = _strb_T_4 ? 16'hff : _strb_T_6; // @[Mux.scala 101:16]
  wire [15:0] _strb_T_8 = _strb_T_3 ? 16'hf : _strb_T_7; // @[Mux.scala 101:16]
  wire [15:0] _strb_T_9 = _strb_T_2 ? 16'h7 : _strb_T_8; // @[Mux.scala 101:16]
  wire [15:0] _strb_T_10 = _strb_T_1 ? 16'h3 : _strb_T_9; // @[Mux.scala 101:16]
  wire [15:0] strb = _strb_T ? 16'h1 : _strb_T_10; // @[Mux.scala 101:16]
  wire [30:0] _GEN_0 = {{15'd0}, strb}; // @[dcache.scala 149:27]
  wire [30:0] _strb_aligned_T = _GEN_0 << cpu_mem_Maddr[3:0]; // @[dcache.scala 149:27]
  wire  _data_array_0_io_i_wen_T_9 = ~victim; // @[dcache.scala 152:157]
  wire [15:0] strb_aligned = _strb_aligned_T[15:0]; // @[dcache.scala 146:24 149:18]
  wire [190:0] _GEN_128 = {{127'd0}, cpu_mem_MdataOut}; // @[dcache.scala 155:104]
  wire [190:0] _data_array_0_io_i_wdata_T_2 = _GEN_128 << _io_cpu_mem_MdataIn_T_1; // @[dcache.scala 155:104]
  wire [190:0] _data_array_0_io_i_wdata_T_3 = hit ? _data_array_0_io_i_wdata_T_2 : {{63'd0},
    io_mem_master_readData_bits_data}; // @[dcache.scala 155:82]
  wire [190:0] _data_array_0_io_i_wdata_T_4 = write_back_is_finishing ? {{63'd0}, read_from_mem_buf} :
    _data_array_0_io_i_wdata_T_3; // @[dcache.scala 155:36]
  wire  _T_3 = _T & _should_write_back_T; // @[dcache.scala 158:30]
  wire  _GEN_3336 = 7'h0 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_775 = 7'h0 == index | valid0_0; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3337 = 7'h1 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_776 = 7'h1 == index | valid0_1; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3338 = 7'h2 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_777 = 7'h2 == index | valid0_2; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3339 = 7'h3 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_778 = 7'h3 == index | valid0_3; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3340 = 7'h4 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_779 = 7'h4 == index | valid0_4; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3341 = 7'h5 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_780 = 7'h5 == index | valid0_5; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3342 = 7'h6 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_781 = 7'h6 == index | valid0_6; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3343 = 7'h7 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_782 = 7'h7 == index | valid0_7; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3344 = 7'h8 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_783 = 7'h8 == index | valid0_8; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3345 = 7'h9 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_784 = 7'h9 == index | valid0_9; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3346 = 7'ha == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_785 = 7'ha == index | valid0_10; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3347 = 7'hb == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_786 = 7'hb == index | valid0_11; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3348 = 7'hc == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_787 = 7'hc == index | valid0_12; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3349 = 7'hd == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_788 = 7'hd == index | valid0_13; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3350 = 7'he == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_789 = 7'he == index | valid0_14; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3351 = 7'hf == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_790 = 7'hf == index | valid0_15; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3352 = 7'h10 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_791 = 7'h10 == index | valid0_16; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3353 = 7'h11 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_792 = 7'h11 == index | valid0_17; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3354 = 7'h12 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_793 = 7'h12 == index | valid0_18; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3355 = 7'h13 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_794 = 7'h13 == index | valid0_19; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3356 = 7'h14 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_795 = 7'h14 == index | valid0_20; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3357 = 7'h15 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_796 = 7'h15 == index | valid0_21; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3358 = 7'h16 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_797 = 7'h16 == index | valid0_22; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3359 = 7'h17 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_798 = 7'h17 == index | valid0_23; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3360 = 7'h18 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_799 = 7'h18 == index | valid0_24; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3361 = 7'h19 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_800 = 7'h19 == index | valid0_25; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3362 = 7'h1a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_801 = 7'h1a == index | valid0_26; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3363 = 7'h1b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_802 = 7'h1b == index | valid0_27; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3364 = 7'h1c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_803 = 7'h1c == index | valid0_28; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3365 = 7'h1d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_804 = 7'h1d == index | valid0_29; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3366 = 7'h1e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_805 = 7'h1e == index | valid0_30; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3367 = 7'h1f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_806 = 7'h1f == index | valid0_31; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3368 = 7'h20 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_807 = 7'h20 == index | valid0_32; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3369 = 7'h21 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_808 = 7'h21 == index | valid0_33; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3370 = 7'h22 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_809 = 7'h22 == index | valid0_34; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3371 = 7'h23 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_810 = 7'h23 == index | valid0_35; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3372 = 7'h24 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_811 = 7'h24 == index | valid0_36; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3373 = 7'h25 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_812 = 7'h25 == index | valid0_37; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3374 = 7'h26 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_813 = 7'h26 == index | valid0_38; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3375 = 7'h27 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_814 = 7'h27 == index | valid0_39; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3376 = 7'h28 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_815 = 7'h28 == index | valid0_40; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3377 = 7'h29 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_816 = 7'h29 == index | valid0_41; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3378 = 7'h2a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_817 = 7'h2a == index | valid0_42; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3379 = 7'h2b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_818 = 7'h2b == index | valid0_43; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3380 = 7'h2c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_819 = 7'h2c == index | valid0_44; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3381 = 7'h2d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_820 = 7'h2d == index | valid0_45; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3382 = 7'h2e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_821 = 7'h2e == index | valid0_46; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3383 = 7'h2f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_822 = 7'h2f == index | valid0_47; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3384 = 7'h30 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_823 = 7'h30 == index | valid0_48; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3385 = 7'h31 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_824 = 7'h31 == index | valid0_49; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3386 = 7'h32 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_825 = 7'h32 == index | valid0_50; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3387 = 7'h33 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_826 = 7'h33 == index | valid0_51; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3388 = 7'h34 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_827 = 7'h34 == index | valid0_52; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3389 = 7'h35 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_828 = 7'h35 == index | valid0_53; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3390 = 7'h36 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_829 = 7'h36 == index | valid0_54; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3391 = 7'h37 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_830 = 7'h37 == index | valid0_55; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3392 = 7'h38 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_831 = 7'h38 == index | valid0_56; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3393 = 7'h39 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_832 = 7'h39 == index | valid0_57; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3394 = 7'h3a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_833 = 7'h3a == index | valid0_58; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3395 = 7'h3b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_834 = 7'h3b == index | valid0_59; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3396 = 7'h3c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_835 = 7'h3c == index | valid0_60; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3397 = 7'h3d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_836 = 7'h3d == index | valid0_61; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3398 = 7'h3e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_837 = 7'h3e == index | valid0_62; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3399 = 7'h3f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_838 = 7'h3f == index | valid0_63; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3400 = 7'h40 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_839 = 7'h40 == index | valid0_64; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3401 = 7'h41 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_840 = 7'h41 == index | valid0_65; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3402 = 7'h42 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_841 = 7'h42 == index | valid0_66; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3403 = 7'h43 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_842 = 7'h43 == index | valid0_67; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3404 = 7'h44 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_843 = 7'h44 == index | valid0_68; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3405 = 7'h45 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_844 = 7'h45 == index | valid0_69; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3406 = 7'h46 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_845 = 7'h46 == index | valid0_70; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3407 = 7'h47 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_846 = 7'h47 == index | valid0_71; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3408 = 7'h48 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_847 = 7'h48 == index | valid0_72; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3409 = 7'h49 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_848 = 7'h49 == index | valid0_73; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3410 = 7'h4a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_849 = 7'h4a == index | valid0_74; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3411 = 7'h4b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_850 = 7'h4b == index | valid0_75; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3412 = 7'h4c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_851 = 7'h4c == index | valid0_76; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3413 = 7'h4d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_852 = 7'h4d == index | valid0_77; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3414 = 7'h4e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_853 = 7'h4e == index | valid0_78; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3415 = 7'h4f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_854 = 7'h4f == index | valid0_79; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3416 = 7'h50 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_855 = 7'h50 == index | valid0_80; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3417 = 7'h51 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_856 = 7'h51 == index | valid0_81; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3418 = 7'h52 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_857 = 7'h52 == index | valid0_82; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3419 = 7'h53 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_858 = 7'h53 == index | valid0_83; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3420 = 7'h54 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_859 = 7'h54 == index | valid0_84; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3421 = 7'h55 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_860 = 7'h55 == index | valid0_85; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3422 = 7'h56 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_861 = 7'h56 == index | valid0_86; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3423 = 7'h57 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_862 = 7'h57 == index | valid0_87; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3424 = 7'h58 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_863 = 7'h58 == index | valid0_88; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3425 = 7'h59 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_864 = 7'h59 == index | valid0_89; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3426 = 7'h5a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_865 = 7'h5a == index | valid0_90; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3427 = 7'h5b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_866 = 7'h5b == index | valid0_91; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3428 = 7'h5c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_867 = 7'h5c == index | valid0_92; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3429 = 7'h5d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_868 = 7'h5d == index | valid0_93; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3430 = 7'h5e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_869 = 7'h5e == index | valid0_94; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3431 = 7'h5f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_870 = 7'h5f == index | valid0_95; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3432 = 7'h60 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_871 = 7'h60 == index | valid0_96; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3433 = 7'h61 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_872 = 7'h61 == index | valid0_97; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3434 = 7'h62 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_873 = 7'h62 == index | valid0_98; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3435 = 7'h63 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_874 = 7'h63 == index | valid0_99; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3436 = 7'h64 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_875 = 7'h64 == index | valid0_100; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3437 = 7'h65 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_876 = 7'h65 == index | valid0_101; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3438 = 7'h66 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_877 = 7'h66 == index | valid0_102; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3439 = 7'h67 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_878 = 7'h67 == index | valid0_103; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3440 = 7'h68 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_879 = 7'h68 == index | valid0_104; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3441 = 7'h69 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_880 = 7'h69 == index | valid0_105; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3442 = 7'h6a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_881 = 7'h6a == index | valid0_106; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3443 = 7'h6b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_882 = 7'h6b == index | valid0_107; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3444 = 7'h6c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_883 = 7'h6c == index | valid0_108; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3445 = 7'h6d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_884 = 7'h6d == index | valid0_109; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3446 = 7'h6e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_885 = 7'h6e == index | valid0_110; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3447 = 7'h6f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_886 = 7'h6f == index | valid0_111; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3448 = 7'h70 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_887 = 7'h70 == index | valid0_112; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3449 = 7'h71 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_888 = 7'h71 == index | valid0_113; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3450 = 7'h72 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_889 = 7'h72 == index | valid0_114; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3451 = 7'h73 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_890 = 7'h73 == index | valid0_115; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3452 = 7'h74 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_891 = 7'h74 == index | valid0_116; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3453 = 7'h75 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_892 = 7'h75 == index | valid0_117; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3454 = 7'h76 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_893 = 7'h76 == index | valid0_118; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3455 = 7'h77 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_894 = 7'h77 == index | valid0_119; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3456 = 7'h78 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_895 = 7'h78 == index | valid0_120; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3457 = 7'h79 == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_896 = 7'h79 == index | valid0_121; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3458 = 7'h7a == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_897 = 7'h7a == index | valid0_122; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3459 = 7'h7b == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_898 = 7'h7b == index | valid0_123; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3460 = 7'h7c == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_899 = 7'h7c == index | valid0_124; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3461 = 7'h7d == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_900 = 7'h7d == index | valid0_125; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3462 = 7'h7e == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_901 = 7'h7e == index | valid0_126; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_3463 = 7'h7f == index; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_902 = 7'h7f == index | valid0_127; // @[dcache.scala 159:{19,19} 48:21]
  wire  _GEN_903 = 7'h0 == index ? 1'h0 : dirty0_0; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_904 = 7'h1 == index ? 1'h0 : dirty0_1; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_905 = 7'h2 == index ? 1'h0 : dirty0_2; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_906 = 7'h3 == index ? 1'h0 : dirty0_3; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_907 = 7'h4 == index ? 1'h0 : dirty0_4; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_908 = 7'h5 == index ? 1'h0 : dirty0_5; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_909 = 7'h6 == index ? 1'h0 : dirty0_6; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_910 = 7'h7 == index ? 1'h0 : dirty0_7; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_911 = 7'h8 == index ? 1'h0 : dirty0_8; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_912 = 7'h9 == index ? 1'h0 : dirty0_9; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_913 = 7'ha == index ? 1'h0 : dirty0_10; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_914 = 7'hb == index ? 1'h0 : dirty0_11; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_915 = 7'hc == index ? 1'h0 : dirty0_12; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_916 = 7'hd == index ? 1'h0 : dirty0_13; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_917 = 7'he == index ? 1'h0 : dirty0_14; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_918 = 7'hf == index ? 1'h0 : dirty0_15; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_919 = 7'h10 == index ? 1'h0 : dirty0_16; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_920 = 7'h11 == index ? 1'h0 : dirty0_17; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_921 = 7'h12 == index ? 1'h0 : dirty0_18; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_922 = 7'h13 == index ? 1'h0 : dirty0_19; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_923 = 7'h14 == index ? 1'h0 : dirty0_20; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_924 = 7'h15 == index ? 1'h0 : dirty0_21; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_925 = 7'h16 == index ? 1'h0 : dirty0_22; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_926 = 7'h17 == index ? 1'h0 : dirty0_23; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_927 = 7'h18 == index ? 1'h0 : dirty0_24; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_928 = 7'h19 == index ? 1'h0 : dirty0_25; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_929 = 7'h1a == index ? 1'h0 : dirty0_26; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_930 = 7'h1b == index ? 1'h0 : dirty0_27; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_931 = 7'h1c == index ? 1'h0 : dirty0_28; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_932 = 7'h1d == index ? 1'h0 : dirty0_29; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_933 = 7'h1e == index ? 1'h0 : dirty0_30; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_934 = 7'h1f == index ? 1'h0 : dirty0_31; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_935 = 7'h20 == index ? 1'h0 : dirty0_32; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_936 = 7'h21 == index ? 1'h0 : dirty0_33; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_937 = 7'h22 == index ? 1'h0 : dirty0_34; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_938 = 7'h23 == index ? 1'h0 : dirty0_35; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_939 = 7'h24 == index ? 1'h0 : dirty0_36; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_940 = 7'h25 == index ? 1'h0 : dirty0_37; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_941 = 7'h26 == index ? 1'h0 : dirty0_38; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_942 = 7'h27 == index ? 1'h0 : dirty0_39; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_943 = 7'h28 == index ? 1'h0 : dirty0_40; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_944 = 7'h29 == index ? 1'h0 : dirty0_41; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_945 = 7'h2a == index ? 1'h0 : dirty0_42; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_946 = 7'h2b == index ? 1'h0 : dirty0_43; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_947 = 7'h2c == index ? 1'h0 : dirty0_44; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_948 = 7'h2d == index ? 1'h0 : dirty0_45; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_949 = 7'h2e == index ? 1'h0 : dirty0_46; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_950 = 7'h2f == index ? 1'h0 : dirty0_47; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_951 = 7'h30 == index ? 1'h0 : dirty0_48; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_952 = 7'h31 == index ? 1'h0 : dirty0_49; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_953 = 7'h32 == index ? 1'h0 : dirty0_50; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_954 = 7'h33 == index ? 1'h0 : dirty0_51; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_955 = 7'h34 == index ? 1'h0 : dirty0_52; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_956 = 7'h35 == index ? 1'h0 : dirty0_53; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_957 = 7'h36 == index ? 1'h0 : dirty0_54; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_958 = 7'h37 == index ? 1'h0 : dirty0_55; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_959 = 7'h38 == index ? 1'h0 : dirty0_56; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_960 = 7'h39 == index ? 1'h0 : dirty0_57; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_961 = 7'h3a == index ? 1'h0 : dirty0_58; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_962 = 7'h3b == index ? 1'h0 : dirty0_59; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_963 = 7'h3c == index ? 1'h0 : dirty0_60; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_964 = 7'h3d == index ? 1'h0 : dirty0_61; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_965 = 7'h3e == index ? 1'h0 : dirty0_62; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_966 = 7'h3f == index ? 1'h0 : dirty0_63; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_967 = 7'h40 == index ? 1'h0 : dirty0_64; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_968 = 7'h41 == index ? 1'h0 : dirty0_65; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_969 = 7'h42 == index ? 1'h0 : dirty0_66; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_970 = 7'h43 == index ? 1'h0 : dirty0_67; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_971 = 7'h44 == index ? 1'h0 : dirty0_68; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_972 = 7'h45 == index ? 1'h0 : dirty0_69; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_973 = 7'h46 == index ? 1'h0 : dirty0_70; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_974 = 7'h47 == index ? 1'h0 : dirty0_71; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_975 = 7'h48 == index ? 1'h0 : dirty0_72; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_976 = 7'h49 == index ? 1'h0 : dirty0_73; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_977 = 7'h4a == index ? 1'h0 : dirty0_74; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_978 = 7'h4b == index ? 1'h0 : dirty0_75; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_979 = 7'h4c == index ? 1'h0 : dirty0_76; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_980 = 7'h4d == index ? 1'h0 : dirty0_77; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_981 = 7'h4e == index ? 1'h0 : dirty0_78; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_982 = 7'h4f == index ? 1'h0 : dirty0_79; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_983 = 7'h50 == index ? 1'h0 : dirty0_80; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_984 = 7'h51 == index ? 1'h0 : dirty0_81; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_985 = 7'h52 == index ? 1'h0 : dirty0_82; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_986 = 7'h53 == index ? 1'h0 : dirty0_83; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_987 = 7'h54 == index ? 1'h0 : dirty0_84; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_988 = 7'h55 == index ? 1'h0 : dirty0_85; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_989 = 7'h56 == index ? 1'h0 : dirty0_86; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_990 = 7'h57 == index ? 1'h0 : dirty0_87; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_991 = 7'h58 == index ? 1'h0 : dirty0_88; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_992 = 7'h59 == index ? 1'h0 : dirty0_89; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_993 = 7'h5a == index ? 1'h0 : dirty0_90; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_994 = 7'h5b == index ? 1'h0 : dirty0_91; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_995 = 7'h5c == index ? 1'h0 : dirty0_92; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_996 = 7'h5d == index ? 1'h0 : dirty0_93; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_997 = 7'h5e == index ? 1'h0 : dirty0_94; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_998 = 7'h5f == index ? 1'h0 : dirty0_95; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_999 = 7'h60 == index ? 1'h0 : dirty0_96; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1000 = 7'h61 == index ? 1'h0 : dirty0_97; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1001 = 7'h62 == index ? 1'h0 : dirty0_98; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1002 = 7'h63 == index ? 1'h0 : dirty0_99; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1003 = 7'h64 == index ? 1'h0 : dirty0_100; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1004 = 7'h65 == index ? 1'h0 : dirty0_101; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1005 = 7'h66 == index ? 1'h0 : dirty0_102; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1006 = 7'h67 == index ? 1'h0 : dirty0_103; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1007 = 7'h68 == index ? 1'h0 : dirty0_104; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1008 = 7'h69 == index ? 1'h0 : dirty0_105; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1009 = 7'h6a == index ? 1'h0 : dirty0_106; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1010 = 7'h6b == index ? 1'h0 : dirty0_107; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1011 = 7'h6c == index ? 1'h0 : dirty0_108; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1012 = 7'h6d == index ? 1'h0 : dirty0_109; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1013 = 7'h6e == index ? 1'h0 : dirty0_110; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1014 = 7'h6f == index ? 1'h0 : dirty0_111; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1015 = 7'h70 == index ? 1'h0 : dirty0_112; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1016 = 7'h71 == index ? 1'h0 : dirty0_113; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1017 = 7'h72 == index ? 1'h0 : dirty0_114; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1018 = 7'h73 == index ? 1'h0 : dirty0_115; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1019 = 7'h74 == index ? 1'h0 : dirty0_116; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1020 = 7'h75 == index ? 1'h0 : dirty0_117; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1021 = 7'h76 == index ? 1'h0 : dirty0_118; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1022 = 7'h77 == index ? 1'h0 : dirty0_119; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1023 = 7'h78 == index ? 1'h0 : dirty0_120; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1024 = 7'h79 == index ? 1'h0 : dirty0_121; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1025 = 7'h7a == index ? 1'h0 : dirty0_122; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1026 = 7'h7b == index ? 1'h0 : dirty0_123; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1027 = 7'h7c == index ? 1'h0 : dirty0_124; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1028 = 7'h7d == index ? 1'h0 : dirty0_125; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1029 = 7'h7e == index ? 1'h0 : dirty0_126; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1030 = 7'h7f == index ? 1'h0 : dirty0_127; // @[dcache.scala 160:{19,19} 50:21]
  wire  _GEN_1287 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_903 :
    dirty0_0; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1288 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_904 :
    dirty0_1; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1289 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_905 :
    dirty0_2; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1290 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_906 :
    dirty0_3; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1291 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_907 :
    dirty0_4; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1292 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_908 :
    dirty0_5; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1293 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_909 :
    dirty0_6; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1294 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_910 :
    dirty0_7; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1295 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_911 :
    dirty0_8; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1296 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_912 :
    dirty0_9; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1297 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_913 :
    dirty0_10; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1298 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_914 :
    dirty0_11; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1299 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_915 :
    dirty0_12; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1300 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_916 :
    dirty0_13; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1301 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_917 :
    dirty0_14; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1302 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_918 :
    dirty0_15; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1303 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_919 :
    dirty0_16; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1304 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_920 :
    dirty0_17; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1305 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_921 :
    dirty0_18; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1306 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_922 :
    dirty0_19; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1307 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_923 :
    dirty0_20; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1308 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_924 :
    dirty0_21; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1309 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_925 :
    dirty0_22; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1310 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_926 :
    dirty0_23; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1311 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_927 :
    dirty0_24; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1312 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_928 :
    dirty0_25; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1313 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_929 :
    dirty0_26; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1314 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_930 :
    dirty0_27; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1315 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_931 :
    dirty0_28; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1316 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_932 :
    dirty0_29; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1317 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_933 :
    dirty0_30; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1318 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_934 :
    dirty0_31; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1319 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_935 :
    dirty0_32; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1320 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_936 :
    dirty0_33; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1321 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_937 :
    dirty0_34; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1322 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_938 :
    dirty0_35; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1323 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_939 :
    dirty0_36; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1324 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_940 :
    dirty0_37; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1325 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_941 :
    dirty0_38; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1326 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_942 :
    dirty0_39; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1327 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_943 :
    dirty0_40; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1328 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_944 :
    dirty0_41; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1329 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_945 :
    dirty0_42; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1330 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_946 :
    dirty0_43; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1331 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_947 :
    dirty0_44; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1332 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_948 :
    dirty0_45; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1333 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_949 :
    dirty0_46; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1334 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_950 :
    dirty0_47; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1335 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_951 :
    dirty0_48; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1336 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_952 :
    dirty0_49; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1337 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_953 :
    dirty0_50; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1338 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_954 :
    dirty0_51; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1339 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_955 :
    dirty0_52; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1340 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_956 :
    dirty0_53; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1341 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_957 :
    dirty0_54; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1342 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_958 :
    dirty0_55; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1343 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_959 :
    dirty0_56; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1344 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_960 :
    dirty0_57; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1345 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_961 :
    dirty0_58; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1346 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_962 :
    dirty0_59; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1347 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_963 :
    dirty0_60; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1348 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_964 :
    dirty0_61; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1349 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_965 :
    dirty0_62; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1350 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_966 :
    dirty0_63; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1351 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_967 :
    dirty0_64; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1352 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_968 :
    dirty0_65; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1353 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_969 :
    dirty0_66; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1354 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_970 :
    dirty0_67; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1355 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_971 :
    dirty0_68; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1356 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_972 :
    dirty0_69; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1357 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_973 :
    dirty0_70; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1358 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_974 :
    dirty0_71; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1359 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_975 :
    dirty0_72; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1360 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_976 :
    dirty0_73; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1361 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_977 :
    dirty0_74; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1362 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_978 :
    dirty0_75; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1363 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_979 :
    dirty0_76; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1364 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_980 :
    dirty0_77; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1365 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_981 :
    dirty0_78; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1366 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_982 :
    dirty0_79; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1367 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_983 :
    dirty0_80; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1368 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_984 :
    dirty0_81; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1369 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_985 :
    dirty0_82; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1370 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_986 :
    dirty0_83; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1371 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_987 :
    dirty0_84; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1372 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_988 :
    dirty0_85; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1373 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_989 :
    dirty0_86; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1374 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_990 :
    dirty0_87; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1375 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_991 :
    dirty0_88; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1376 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_992 :
    dirty0_89; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1377 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_993 :
    dirty0_90; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1378 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_994 :
    dirty0_91; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1379 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_995 :
    dirty0_92; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1380 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_996 :
    dirty0_93; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1381 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_997 :
    dirty0_94; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1382 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_998 :
    dirty0_95; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1383 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_999 :
    dirty0_96; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1384 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1000 :
    dirty0_97; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1385 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1001 :
    dirty0_98; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1386 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1002 :
    dirty0_99; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1387 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1003 :
    dirty0_100; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1388 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1004 :
    dirty0_101; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1389 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1005 :
    dirty0_102; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1390 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1006 :
    dirty0_103; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1391 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1007 :
    dirty0_104; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1392 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1008 :
    dirty0_105; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1393 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1009 :
    dirty0_106; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1394 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1010 :
    dirty0_107; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1395 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1011 :
    dirty0_108; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1396 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1012 :
    dirty0_109; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1397 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1013 :
    dirty0_110; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1398 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1014 :
    dirty0_111; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1399 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1015 :
    dirty0_112; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1400 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1016 :
    dirty0_113; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1401 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1017 :
    dirty0_114; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1402 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1018 :
    dirty0_115; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1403 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1019 :
    dirty0_116; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1404 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1020 :
    dirty0_117; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1405 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1021 :
    dirty0_118; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1406 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1022 :
    dirty0_119; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1407 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1023 :
    dirty0_120; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1408 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1024 :
    dirty0_121; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1409 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1025 :
    dirty0_122; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1410 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1026 :
    dirty0_123; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1411 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1027 :
    dirty0_124; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1412 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1028 :
    dirty0_125; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1413 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1029 :
    dirty0_126; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1414 = _T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T ? _GEN_1030 :
    dirty0_127; // @[dcache.scala 158:91 50:21]
  wire  _GEN_1543 = _GEN_3336 | valid1_0; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1544 = _GEN_3337 | valid1_1; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1545 = _GEN_3338 | valid1_2; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1546 = _GEN_3339 | valid1_3; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1547 = _GEN_3340 | valid1_4; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1548 = _GEN_3341 | valid1_5; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1549 = _GEN_3342 | valid1_6; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1550 = _GEN_3343 | valid1_7; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1551 = _GEN_3344 | valid1_8; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1552 = _GEN_3345 | valid1_9; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1553 = _GEN_3346 | valid1_10; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1554 = _GEN_3347 | valid1_11; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1555 = _GEN_3348 | valid1_12; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1556 = _GEN_3349 | valid1_13; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1557 = _GEN_3350 | valid1_14; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1558 = _GEN_3351 | valid1_15; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1559 = _GEN_3352 | valid1_16; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1560 = _GEN_3353 | valid1_17; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1561 = _GEN_3354 | valid1_18; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1562 = _GEN_3355 | valid1_19; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1563 = _GEN_3356 | valid1_20; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1564 = _GEN_3357 | valid1_21; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1565 = _GEN_3358 | valid1_22; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1566 = _GEN_3359 | valid1_23; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1567 = _GEN_3360 | valid1_24; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1568 = _GEN_3361 | valid1_25; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1569 = _GEN_3362 | valid1_26; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1570 = _GEN_3363 | valid1_27; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1571 = _GEN_3364 | valid1_28; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1572 = _GEN_3365 | valid1_29; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1573 = _GEN_3366 | valid1_30; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1574 = _GEN_3367 | valid1_31; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1575 = _GEN_3368 | valid1_32; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1576 = _GEN_3369 | valid1_33; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1577 = _GEN_3370 | valid1_34; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1578 = _GEN_3371 | valid1_35; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1579 = _GEN_3372 | valid1_36; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1580 = _GEN_3373 | valid1_37; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1581 = _GEN_3374 | valid1_38; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1582 = _GEN_3375 | valid1_39; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1583 = _GEN_3376 | valid1_40; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1584 = _GEN_3377 | valid1_41; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1585 = _GEN_3378 | valid1_42; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1586 = _GEN_3379 | valid1_43; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1587 = _GEN_3380 | valid1_44; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1588 = _GEN_3381 | valid1_45; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1589 = _GEN_3382 | valid1_46; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1590 = _GEN_3383 | valid1_47; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1591 = _GEN_3384 | valid1_48; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1592 = _GEN_3385 | valid1_49; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1593 = _GEN_3386 | valid1_50; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1594 = _GEN_3387 | valid1_51; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1595 = _GEN_3388 | valid1_52; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1596 = _GEN_3389 | valid1_53; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1597 = _GEN_3390 | valid1_54; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1598 = _GEN_3391 | valid1_55; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1599 = _GEN_3392 | valid1_56; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1600 = _GEN_3393 | valid1_57; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1601 = _GEN_3394 | valid1_58; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1602 = _GEN_3395 | valid1_59; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1603 = _GEN_3396 | valid1_60; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1604 = _GEN_3397 | valid1_61; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1605 = _GEN_3398 | valid1_62; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1606 = _GEN_3399 | valid1_63; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1607 = _GEN_3400 | valid1_64; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1608 = _GEN_3401 | valid1_65; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1609 = _GEN_3402 | valid1_66; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1610 = _GEN_3403 | valid1_67; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1611 = _GEN_3404 | valid1_68; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1612 = _GEN_3405 | valid1_69; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1613 = _GEN_3406 | valid1_70; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1614 = _GEN_3407 | valid1_71; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1615 = _GEN_3408 | valid1_72; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1616 = _GEN_3409 | valid1_73; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1617 = _GEN_3410 | valid1_74; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1618 = _GEN_3411 | valid1_75; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1619 = _GEN_3412 | valid1_76; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1620 = _GEN_3413 | valid1_77; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1621 = _GEN_3414 | valid1_78; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1622 = _GEN_3415 | valid1_79; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1623 = _GEN_3416 | valid1_80; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1624 = _GEN_3417 | valid1_81; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1625 = _GEN_3418 | valid1_82; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1626 = _GEN_3419 | valid1_83; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1627 = _GEN_3420 | valid1_84; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1628 = _GEN_3421 | valid1_85; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1629 = _GEN_3422 | valid1_86; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1630 = _GEN_3423 | valid1_87; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1631 = _GEN_3424 | valid1_88; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1632 = _GEN_3425 | valid1_89; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1633 = _GEN_3426 | valid1_90; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1634 = _GEN_3427 | valid1_91; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1635 = _GEN_3428 | valid1_92; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1636 = _GEN_3429 | valid1_93; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1637 = _GEN_3430 | valid1_94; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1638 = _GEN_3431 | valid1_95; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1639 = _GEN_3432 | valid1_96; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1640 = _GEN_3433 | valid1_97; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1641 = _GEN_3434 | valid1_98; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1642 = _GEN_3435 | valid1_99; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1643 = _GEN_3436 | valid1_100; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1644 = _GEN_3437 | valid1_101; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1645 = _GEN_3438 | valid1_102; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1646 = _GEN_3439 | valid1_103; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1647 = _GEN_3440 | valid1_104; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1648 = _GEN_3441 | valid1_105; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1649 = _GEN_3442 | valid1_106; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1650 = _GEN_3443 | valid1_107; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1651 = _GEN_3444 | valid1_108; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1652 = _GEN_3445 | valid1_109; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1653 = _GEN_3446 | valid1_110; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1654 = _GEN_3447 | valid1_111; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1655 = _GEN_3448 | valid1_112; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1656 = _GEN_3449 | valid1_113; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1657 = _GEN_3450 | valid1_114; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1658 = _GEN_3451 | valid1_115; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1659 = _GEN_3452 | valid1_116; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1660 = _GEN_3453 | valid1_117; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1661 = _GEN_3454 | valid1_118; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1662 = _GEN_3455 | valid1_119; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1663 = _GEN_3456 | valid1_120; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1664 = _GEN_3457 | valid1_121; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1665 = _GEN_3458 | valid1_122; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1666 = _GEN_3459 | valid1_123; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1667 = _GEN_3460 | valid1_124; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1668 = _GEN_3461 | valid1_125; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1669 = _GEN_3462 | valid1_126; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1670 = _GEN_3463 | valid1_127; // @[dcache.scala 164:{19,19} 49:21]
  wire  _GEN_1671 = 7'h0 == index ? 1'h0 : dirty1_0; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1672 = 7'h1 == index ? 1'h0 : dirty1_1; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1673 = 7'h2 == index ? 1'h0 : dirty1_2; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1674 = 7'h3 == index ? 1'h0 : dirty1_3; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1675 = 7'h4 == index ? 1'h0 : dirty1_4; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1676 = 7'h5 == index ? 1'h0 : dirty1_5; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1677 = 7'h6 == index ? 1'h0 : dirty1_6; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1678 = 7'h7 == index ? 1'h0 : dirty1_7; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1679 = 7'h8 == index ? 1'h0 : dirty1_8; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1680 = 7'h9 == index ? 1'h0 : dirty1_9; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1681 = 7'ha == index ? 1'h0 : dirty1_10; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1682 = 7'hb == index ? 1'h0 : dirty1_11; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1683 = 7'hc == index ? 1'h0 : dirty1_12; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1684 = 7'hd == index ? 1'h0 : dirty1_13; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1685 = 7'he == index ? 1'h0 : dirty1_14; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1686 = 7'hf == index ? 1'h0 : dirty1_15; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1687 = 7'h10 == index ? 1'h0 : dirty1_16; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1688 = 7'h11 == index ? 1'h0 : dirty1_17; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1689 = 7'h12 == index ? 1'h0 : dirty1_18; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1690 = 7'h13 == index ? 1'h0 : dirty1_19; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1691 = 7'h14 == index ? 1'h0 : dirty1_20; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1692 = 7'h15 == index ? 1'h0 : dirty1_21; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1693 = 7'h16 == index ? 1'h0 : dirty1_22; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1694 = 7'h17 == index ? 1'h0 : dirty1_23; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1695 = 7'h18 == index ? 1'h0 : dirty1_24; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1696 = 7'h19 == index ? 1'h0 : dirty1_25; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1697 = 7'h1a == index ? 1'h0 : dirty1_26; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1698 = 7'h1b == index ? 1'h0 : dirty1_27; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1699 = 7'h1c == index ? 1'h0 : dirty1_28; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1700 = 7'h1d == index ? 1'h0 : dirty1_29; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1701 = 7'h1e == index ? 1'h0 : dirty1_30; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1702 = 7'h1f == index ? 1'h0 : dirty1_31; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1703 = 7'h20 == index ? 1'h0 : dirty1_32; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1704 = 7'h21 == index ? 1'h0 : dirty1_33; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1705 = 7'h22 == index ? 1'h0 : dirty1_34; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1706 = 7'h23 == index ? 1'h0 : dirty1_35; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1707 = 7'h24 == index ? 1'h0 : dirty1_36; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1708 = 7'h25 == index ? 1'h0 : dirty1_37; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1709 = 7'h26 == index ? 1'h0 : dirty1_38; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1710 = 7'h27 == index ? 1'h0 : dirty1_39; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1711 = 7'h28 == index ? 1'h0 : dirty1_40; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1712 = 7'h29 == index ? 1'h0 : dirty1_41; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1713 = 7'h2a == index ? 1'h0 : dirty1_42; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1714 = 7'h2b == index ? 1'h0 : dirty1_43; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1715 = 7'h2c == index ? 1'h0 : dirty1_44; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1716 = 7'h2d == index ? 1'h0 : dirty1_45; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1717 = 7'h2e == index ? 1'h0 : dirty1_46; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1718 = 7'h2f == index ? 1'h0 : dirty1_47; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1719 = 7'h30 == index ? 1'h0 : dirty1_48; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1720 = 7'h31 == index ? 1'h0 : dirty1_49; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1721 = 7'h32 == index ? 1'h0 : dirty1_50; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1722 = 7'h33 == index ? 1'h0 : dirty1_51; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1723 = 7'h34 == index ? 1'h0 : dirty1_52; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1724 = 7'h35 == index ? 1'h0 : dirty1_53; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1725 = 7'h36 == index ? 1'h0 : dirty1_54; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1726 = 7'h37 == index ? 1'h0 : dirty1_55; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1727 = 7'h38 == index ? 1'h0 : dirty1_56; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1728 = 7'h39 == index ? 1'h0 : dirty1_57; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1729 = 7'h3a == index ? 1'h0 : dirty1_58; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1730 = 7'h3b == index ? 1'h0 : dirty1_59; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1731 = 7'h3c == index ? 1'h0 : dirty1_60; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1732 = 7'h3d == index ? 1'h0 : dirty1_61; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1733 = 7'h3e == index ? 1'h0 : dirty1_62; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1734 = 7'h3f == index ? 1'h0 : dirty1_63; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1735 = 7'h40 == index ? 1'h0 : dirty1_64; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1736 = 7'h41 == index ? 1'h0 : dirty1_65; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1737 = 7'h42 == index ? 1'h0 : dirty1_66; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1738 = 7'h43 == index ? 1'h0 : dirty1_67; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1739 = 7'h44 == index ? 1'h0 : dirty1_68; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1740 = 7'h45 == index ? 1'h0 : dirty1_69; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1741 = 7'h46 == index ? 1'h0 : dirty1_70; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1742 = 7'h47 == index ? 1'h0 : dirty1_71; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1743 = 7'h48 == index ? 1'h0 : dirty1_72; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1744 = 7'h49 == index ? 1'h0 : dirty1_73; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1745 = 7'h4a == index ? 1'h0 : dirty1_74; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1746 = 7'h4b == index ? 1'h0 : dirty1_75; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1747 = 7'h4c == index ? 1'h0 : dirty1_76; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1748 = 7'h4d == index ? 1'h0 : dirty1_77; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1749 = 7'h4e == index ? 1'h0 : dirty1_78; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1750 = 7'h4f == index ? 1'h0 : dirty1_79; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1751 = 7'h50 == index ? 1'h0 : dirty1_80; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1752 = 7'h51 == index ? 1'h0 : dirty1_81; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1753 = 7'h52 == index ? 1'h0 : dirty1_82; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1754 = 7'h53 == index ? 1'h0 : dirty1_83; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1755 = 7'h54 == index ? 1'h0 : dirty1_84; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1756 = 7'h55 == index ? 1'h0 : dirty1_85; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1757 = 7'h56 == index ? 1'h0 : dirty1_86; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1758 = 7'h57 == index ? 1'h0 : dirty1_87; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1759 = 7'h58 == index ? 1'h0 : dirty1_88; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1760 = 7'h59 == index ? 1'h0 : dirty1_89; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1761 = 7'h5a == index ? 1'h0 : dirty1_90; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1762 = 7'h5b == index ? 1'h0 : dirty1_91; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1763 = 7'h5c == index ? 1'h0 : dirty1_92; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1764 = 7'h5d == index ? 1'h0 : dirty1_93; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1765 = 7'h5e == index ? 1'h0 : dirty1_94; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1766 = 7'h5f == index ? 1'h0 : dirty1_95; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1767 = 7'h60 == index ? 1'h0 : dirty1_96; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1768 = 7'h61 == index ? 1'h0 : dirty1_97; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1769 = 7'h62 == index ? 1'h0 : dirty1_98; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1770 = 7'h63 == index ? 1'h0 : dirty1_99; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1771 = 7'h64 == index ? 1'h0 : dirty1_100; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1772 = 7'h65 == index ? 1'h0 : dirty1_101; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1773 = 7'h66 == index ? 1'h0 : dirty1_102; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1774 = 7'h67 == index ? 1'h0 : dirty1_103; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1775 = 7'h68 == index ? 1'h0 : dirty1_104; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1776 = 7'h69 == index ? 1'h0 : dirty1_105; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1777 = 7'h6a == index ? 1'h0 : dirty1_106; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1778 = 7'h6b == index ? 1'h0 : dirty1_107; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1779 = 7'h6c == index ? 1'h0 : dirty1_108; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1780 = 7'h6d == index ? 1'h0 : dirty1_109; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1781 = 7'h6e == index ? 1'h0 : dirty1_110; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1782 = 7'h6f == index ? 1'h0 : dirty1_111; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1783 = 7'h70 == index ? 1'h0 : dirty1_112; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1784 = 7'h71 == index ? 1'h0 : dirty1_113; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1785 = 7'h72 == index ? 1'h0 : dirty1_114; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1786 = 7'h73 == index ? 1'h0 : dirty1_115; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1787 = 7'h74 == index ? 1'h0 : dirty1_116; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1788 = 7'h75 == index ? 1'h0 : dirty1_117; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1789 = 7'h76 == index ? 1'h0 : dirty1_118; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1790 = 7'h77 == index ? 1'h0 : dirty1_119; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1791 = 7'h78 == index ? 1'h0 : dirty1_120; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1792 = 7'h79 == index ? 1'h0 : dirty1_121; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1793 = 7'h7a == index ? 1'h0 : dirty1_122; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1794 = 7'h7b == index ? 1'h0 : dirty1_123; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1795 = 7'h7c == index ? 1'h0 : dirty1_124; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1796 = 7'h7d == index ? 1'h0 : dirty1_125; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1797 = 7'h7e == index ? 1'h0 : dirty1_126; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_1798 = 7'h7f == index ? 1'h0 : dirty1_127; // @[dcache.scala 165:{19,19} 51:21]
  wire  _GEN_2055 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1671 : dirty1_0; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2056 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1672 : dirty1_1; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2057 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1673 : dirty1_2; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2058 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1674 : dirty1_3; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2059 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1675 : dirty1_4; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2060 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1676 : dirty1_5; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2061 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1677 : dirty1_6; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2062 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1678 : dirty1_7; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2063 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1679 : dirty1_8; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2064 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1680 : dirty1_9; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2065 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1681 : dirty1_10; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2066 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1682 : dirty1_11; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2067 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1683 : dirty1_12; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2068 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1684 : dirty1_13; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2069 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1685 : dirty1_14; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2070 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1686 : dirty1_15; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2071 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1687 : dirty1_16; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2072 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1688 : dirty1_17; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2073 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1689 : dirty1_18; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2074 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1690 : dirty1_19; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2075 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1691 : dirty1_20; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2076 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1692 : dirty1_21; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2077 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1693 : dirty1_22; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2078 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1694 : dirty1_23; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2079 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1695 : dirty1_24; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2080 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1696 : dirty1_25; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2081 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1697 : dirty1_26; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2082 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1698 : dirty1_27; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2083 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1699 : dirty1_28; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2084 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1700 : dirty1_29; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2085 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1701 : dirty1_30; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2086 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1702 : dirty1_31; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2087 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1703 : dirty1_32; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2088 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1704 : dirty1_33; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2089 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1705 : dirty1_34; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2090 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1706 : dirty1_35; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2091 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1707 : dirty1_36; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2092 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1708 : dirty1_37; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2093 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1709 : dirty1_38; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2094 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1710 : dirty1_39; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2095 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1711 : dirty1_40; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2096 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1712 : dirty1_41; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2097 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1713 : dirty1_42; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2098 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1714 : dirty1_43; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2099 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1715 : dirty1_44; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2100 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1716 : dirty1_45; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2101 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1717 : dirty1_46; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2102 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1718 : dirty1_47; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2103 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1719 : dirty1_48; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2104 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1720 : dirty1_49; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2105 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1721 : dirty1_50; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2106 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1722 : dirty1_51; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2107 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1723 : dirty1_52; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2108 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1724 : dirty1_53; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2109 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1725 : dirty1_54; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2110 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1726 : dirty1_55; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2111 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1727 : dirty1_56; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2112 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1728 : dirty1_57; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2113 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1729 : dirty1_58; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2114 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1730 : dirty1_59; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2115 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1731 : dirty1_60; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2116 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1732 : dirty1_61; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2117 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1733 : dirty1_62; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2118 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1734 : dirty1_63; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2119 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1735 : dirty1_64; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2120 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1736 : dirty1_65; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2121 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1737 : dirty1_66; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2122 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1738 : dirty1_67; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2123 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1739 : dirty1_68; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2124 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1740 : dirty1_69; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2125 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1741 : dirty1_70; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2126 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1742 : dirty1_71; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2127 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1743 : dirty1_72; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2128 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1744 : dirty1_73; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2129 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1745 : dirty1_74; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2130 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1746 : dirty1_75; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2131 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1747 : dirty1_76; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2132 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1748 : dirty1_77; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2133 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1749 : dirty1_78; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2134 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1750 : dirty1_79; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2135 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1751 : dirty1_80; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2136 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1752 : dirty1_81; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2137 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1753 : dirty1_82; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2138 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1754 : dirty1_83; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2139 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1755 : dirty1_84; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2140 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1756 : dirty1_85; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2141 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1757 : dirty1_86; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2142 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1758 : dirty1_87; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2143 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1759 : dirty1_88; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2144 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1760 : dirty1_89; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2145 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1761 : dirty1_90; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2146 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1762 : dirty1_91; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2147 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1763 : dirty1_92; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2148 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1764 : dirty1_93; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2149 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1765 : dirty1_94; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2150 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1766 : dirty1_95; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2151 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1767 : dirty1_96; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2152 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1768 : dirty1_97; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2153 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1769 : dirty1_98; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2154 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1770 : dirty1_99; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2155 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1771 : dirty1_100; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2156 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1772 : dirty1_101; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2157 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1773 : dirty1_102; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2158 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1774 : dirty1_103; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2159 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1775 : dirty1_104; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2160 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1776 : dirty1_105; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2161 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1777 : dirty1_106; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2162 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1778 : dirty1_107; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2163 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1779 : dirty1_108; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2164 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1780 : dirty1_109; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2165 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1781 : dirty1_110; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2166 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1782 : dirty1_111; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2167 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1783 : dirty1_112; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2168 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1784 : dirty1_113; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2169 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1785 : dirty1_114; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2170 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1786 : dirty1_115; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2171 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1787 : dirty1_116; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2172 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1788 : dirty1_117; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2173 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1789 : dirty1_118; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2174 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1790 : dirty1_119; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2175 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1791 : dirty1_120; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2176 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1792 : dirty1_121; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2177 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1793 : dirty1_122; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2178 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1794 : dirty1_123; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2179 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1795 : dirty1_124; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2180 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1796 : dirty1_125; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2181 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1797 : dirty1_126; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2182 = _T_3 & victim & _write_back_is_finishing_T ? _GEN_1798 : dirty1_127; // @[dcache.scala 163:91 51:21]
  wire  _GEN_2311 = _GEN_3336 | _GEN_1287; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2312 = _GEN_3337 | _GEN_1288; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2313 = _GEN_3338 | _GEN_1289; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2314 = _GEN_3339 | _GEN_1290; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2315 = _GEN_3340 | _GEN_1291; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2316 = _GEN_3341 | _GEN_1292; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2317 = _GEN_3342 | _GEN_1293; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2318 = _GEN_3343 | _GEN_1294; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2319 = _GEN_3344 | _GEN_1295; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2320 = _GEN_3345 | _GEN_1296; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2321 = _GEN_3346 | _GEN_1297; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2322 = _GEN_3347 | _GEN_1298; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2323 = _GEN_3348 | _GEN_1299; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2324 = _GEN_3349 | _GEN_1300; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2325 = _GEN_3350 | _GEN_1301; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2326 = _GEN_3351 | _GEN_1302; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2327 = _GEN_3352 | _GEN_1303; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2328 = _GEN_3353 | _GEN_1304; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2329 = _GEN_3354 | _GEN_1305; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2330 = _GEN_3355 | _GEN_1306; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2331 = _GEN_3356 | _GEN_1307; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2332 = _GEN_3357 | _GEN_1308; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2333 = _GEN_3358 | _GEN_1309; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2334 = _GEN_3359 | _GEN_1310; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2335 = _GEN_3360 | _GEN_1311; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2336 = _GEN_3361 | _GEN_1312; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2337 = _GEN_3362 | _GEN_1313; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2338 = _GEN_3363 | _GEN_1314; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2339 = _GEN_3364 | _GEN_1315; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2340 = _GEN_3365 | _GEN_1316; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2341 = _GEN_3366 | _GEN_1317; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2342 = _GEN_3367 | _GEN_1318; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2343 = _GEN_3368 | _GEN_1319; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2344 = _GEN_3369 | _GEN_1320; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2345 = _GEN_3370 | _GEN_1321; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2346 = _GEN_3371 | _GEN_1322; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2347 = _GEN_3372 | _GEN_1323; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2348 = _GEN_3373 | _GEN_1324; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2349 = _GEN_3374 | _GEN_1325; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2350 = _GEN_3375 | _GEN_1326; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2351 = _GEN_3376 | _GEN_1327; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2352 = _GEN_3377 | _GEN_1328; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2353 = _GEN_3378 | _GEN_1329; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2354 = _GEN_3379 | _GEN_1330; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2355 = _GEN_3380 | _GEN_1331; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2356 = _GEN_3381 | _GEN_1332; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2357 = _GEN_3382 | _GEN_1333; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2358 = _GEN_3383 | _GEN_1334; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2359 = _GEN_3384 | _GEN_1335; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2360 = _GEN_3385 | _GEN_1336; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2361 = _GEN_3386 | _GEN_1337; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2362 = _GEN_3387 | _GEN_1338; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2363 = _GEN_3388 | _GEN_1339; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2364 = _GEN_3389 | _GEN_1340; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2365 = _GEN_3390 | _GEN_1341; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2366 = _GEN_3391 | _GEN_1342; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2367 = _GEN_3392 | _GEN_1343; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2368 = _GEN_3393 | _GEN_1344; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2369 = _GEN_3394 | _GEN_1345; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2370 = _GEN_3395 | _GEN_1346; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2371 = _GEN_3396 | _GEN_1347; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2372 = _GEN_3397 | _GEN_1348; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2373 = _GEN_3398 | _GEN_1349; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2374 = _GEN_3399 | _GEN_1350; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2375 = _GEN_3400 | _GEN_1351; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2376 = _GEN_3401 | _GEN_1352; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2377 = _GEN_3402 | _GEN_1353; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2378 = _GEN_3403 | _GEN_1354; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2379 = _GEN_3404 | _GEN_1355; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2380 = _GEN_3405 | _GEN_1356; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2381 = _GEN_3406 | _GEN_1357; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2382 = _GEN_3407 | _GEN_1358; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2383 = _GEN_3408 | _GEN_1359; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2384 = _GEN_3409 | _GEN_1360; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2385 = _GEN_3410 | _GEN_1361; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2386 = _GEN_3411 | _GEN_1362; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2387 = _GEN_3412 | _GEN_1363; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2388 = _GEN_3413 | _GEN_1364; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2389 = _GEN_3414 | _GEN_1365; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2390 = _GEN_3415 | _GEN_1366; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2391 = _GEN_3416 | _GEN_1367; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2392 = _GEN_3417 | _GEN_1368; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2393 = _GEN_3418 | _GEN_1369; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2394 = _GEN_3419 | _GEN_1370; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2395 = _GEN_3420 | _GEN_1371; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2396 = _GEN_3421 | _GEN_1372; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2397 = _GEN_3422 | _GEN_1373; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2398 = _GEN_3423 | _GEN_1374; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2399 = _GEN_3424 | _GEN_1375; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2400 = _GEN_3425 | _GEN_1376; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2401 = _GEN_3426 | _GEN_1377; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2402 = _GEN_3427 | _GEN_1378; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2403 = _GEN_3428 | _GEN_1379; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2404 = _GEN_3429 | _GEN_1380; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2405 = _GEN_3430 | _GEN_1381; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2406 = _GEN_3431 | _GEN_1382; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2407 = _GEN_3432 | _GEN_1383; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2408 = _GEN_3433 | _GEN_1384; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2409 = _GEN_3434 | _GEN_1385; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2410 = _GEN_3435 | _GEN_1386; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2411 = _GEN_3436 | _GEN_1387; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2412 = _GEN_3437 | _GEN_1388; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2413 = _GEN_3438 | _GEN_1389; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2414 = _GEN_3439 | _GEN_1390; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2415 = _GEN_3440 | _GEN_1391; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2416 = _GEN_3441 | _GEN_1392; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2417 = _GEN_3442 | _GEN_1393; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2418 = _GEN_3443 | _GEN_1394; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2419 = _GEN_3444 | _GEN_1395; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2420 = _GEN_3445 | _GEN_1396; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2421 = _GEN_3446 | _GEN_1397; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2422 = _GEN_3447 | _GEN_1398; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2423 = _GEN_3448 | _GEN_1399; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2424 = _GEN_3449 | _GEN_1400; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2425 = _GEN_3450 | _GEN_1401; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2426 = _GEN_3451 | _GEN_1402; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2427 = _GEN_3452 | _GEN_1403; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2428 = _GEN_3453 | _GEN_1404; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2429 = _GEN_3454 | _GEN_1405; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2430 = _GEN_3455 | _GEN_1406; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2431 = _GEN_3456 | _GEN_1407; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2432 = _GEN_3457 | _GEN_1408; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2433 = _GEN_3458 | _GEN_1409; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2434 = _GEN_3459 | _GEN_1410; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2435 = _GEN_3460 | _GEN_1411; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2436 = _GEN_3461 | _GEN_1412; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2437 = _GEN_3462 | _GEN_1413; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2438 = _GEN_3463 | _GEN_1414; // @[dcache.scala 169:{19,19}]
  wire  _GEN_2439 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2311 : _GEN_1287; // @[dcache.scala 168:42]
  wire  _GEN_2440 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2312 : _GEN_1288; // @[dcache.scala 168:42]
  wire  _GEN_2441 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2313 : _GEN_1289; // @[dcache.scala 168:42]
  wire  _GEN_2442 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2314 : _GEN_1290; // @[dcache.scala 168:42]
  wire  _GEN_2443 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2315 : _GEN_1291; // @[dcache.scala 168:42]
  wire  _GEN_2444 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2316 : _GEN_1292; // @[dcache.scala 168:42]
  wire  _GEN_2445 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2317 : _GEN_1293; // @[dcache.scala 168:42]
  wire  _GEN_2446 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2318 : _GEN_1294; // @[dcache.scala 168:42]
  wire  _GEN_2447 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2319 : _GEN_1295; // @[dcache.scala 168:42]
  wire  _GEN_2448 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2320 : _GEN_1296; // @[dcache.scala 168:42]
  wire  _GEN_2449 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2321 : _GEN_1297; // @[dcache.scala 168:42]
  wire  _GEN_2450 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2322 : _GEN_1298; // @[dcache.scala 168:42]
  wire  _GEN_2451 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2323 : _GEN_1299; // @[dcache.scala 168:42]
  wire  _GEN_2452 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2324 : _GEN_1300; // @[dcache.scala 168:42]
  wire  _GEN_2453 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2325 : _GEN_1301; // @[dcache.scala 168:42]
  wire  _GEN_2454 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2326 : _GEN_1302; // @[dcache.scala 168:42]
  wire  _GEN_2455 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2327 : _GEN_1303; // @[dcache.scala 168:42]
  wire  _GEN_2456 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2328 : _GEN_1304; // @[dcache.scala 168:42]
  wire  _GEN_2457 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2329 : _GEN_1305; // @[dcache.scala 168:42]
  wire  _GEN_2458 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2330 : _GEN_1306; // @[dcache.scala 168:42]
  wire  _GEN_2459 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2331 : _GEN_1307; // @[dcache.scala 168:42]
  wire  _GEN_2460 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2332 : _GEN_1308; // @[dcache.scala 168:42]
  wire  _GEN_2461 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2333 : _GEN_1309; // @[dcache.scala 168:42]
  wire  _GEN_2462 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2334 : _GEN_1310; // @[dcache.scala 168:42]
  wire  _GEN_2463 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2335 : _GEN_1311; // @[dcache.scala 168:42]
  wire  _GEN_2464 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2336 : _GEN_1312; // @[dcache.scala 168:42]
  wire  _GEN_2465 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2337 : _GEN_1313; // @[dcache.scala 168:42]
  wire  _GEN_2466 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2338 : _GEN_1314; // @[dcache.scala 168:42]
  wire  _GEN_2467 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2339 : _GEN_1315; // @[dcache.scala 168:42]
  wire  _GEN_2468 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2340 : _GEN_1316; // @[dcache.scala 168:42]
  wire  _GEN_2469 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2341 : _GEN_1317; // @[dcache.scala 168:42]
  wire  _GEN_2470 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2342 : _GEN_1318; // @[dcache.scala 168:42]
  wire  _GEN_2471 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2343 : _GEN_1319; // @[dcache.scala 168:42]
  wire  _GEN_2472 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2344 : _GEN_1320; // @[dcache.scala 168:42]
  wire  _GEN_2473 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2345 : _GEN_1321; // @[dcache.scala 168:42]
  wire  _GEN_2474 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2346 : _GEN_1322; // @[dcache.scala 168:42]
  wire  _GEN_2475 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2347 : _GEN_1323; // @[dcache.scala 168:42]
  wire  _GEN_2476 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2348 : _GEN_1324; // @[dcache.scala 168:42]
  wire  _GEN_2477 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2349 : _GEN_1325; // @[dcache.scala 168:42]
  wire  _GEN_2478 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2350 : _GEN_1326; // @[dcache.scala 168:42]
  wire  _GEN_2479 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2351 : _GEN_1327; // @[dcache.scala 168:42]
  wire  _GEN_2480 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2352 : _GEN_1328; // @[dcache.scala 168:42]
  wire  _GEN_2481 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2353 : _GEN_1329; // @[dcache.scala 168:42]
  wire  _GEN_2482 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2354 : _GEN_1330; // @[dcache.scala 168:42]
  wire  _GEN_2483 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2355 : _GEN_1331; // @[dcache.scala 168:42]
  wire  _GEN_2484 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2356 : _GEN_1332; // @[dcache.scala 168:42]
  wire  _GEN_2485 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2357 : _GEN_1333; // @[dcache.scala 168:42]
  wire  _GEN_2486 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2358 : _GEN_1334; // @[dcache.scala 168:42]
  wire  _GEN_2487 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2359 : _GEN_1335; // @[dcache.scala 168:42]
  wire  _GEN_2488 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2360 : _GEN_1336; // @[dcache.scala 168:42]
  wire  _GEN_2489 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2361 : _GEN_1337; // @[dcache.scala 168:42]
  wire  _GEN_2490 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2362 : _GEN_1338; // @[dcache.scala 168:42]
  wire  _GEN_2491 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2363 : _GEN_1339; // @[dcache.scala 168:42]
  wire  _GEN_2492 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2364 : _GEN_1340; // @[dcache.scala 168:42]
  wire  _GEN_2493 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2365 : _GEN_1341; // @[dcache.scala 168:42]
  wire  _GEN_2494 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2366 : _GEN_1342; // @[dcache.scala 168:42]
  wire  _GEN_2495 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2367 : _GEN_1343; // @[dcache.scala 168:42]
  wire  _GEN_2496 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2368 : _GEN_1344; // @[dcache.scala 168:42]
  wire  _GEN_2497 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2369 : _GEN_1345; // @[dcache.scala 168:42]
  wire  _GEN_2498 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2370 : _GEN_1346; // @[dcache.scala 168:42]
  wire  _GEN_2499 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2371 : _GEN_1347; // @[dcache.scala 168:42]
  wire  _GEN_2500 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2372 : _GEN_1348; // @[dcache.scala 168:42]
  wire  _GEN_2501 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2373 : _GEN_1349; // @[dcache.scala 168:42]
  wire  _GEN_2502 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2374 : _GEN_1350; // @[dcache.scala 168:42]
  wire  _GEN_2503 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2375 : _GEN_1351; // @[dcache.scala 168:42]
  wire  _GEN_2504 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2376 : _GEN_1352; // @[dcache.scala 168:42]
  wire  _GEN_2505 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2377 : _GEN_1353; // @[dcache.scala 168:42]
  wire  _GEN_2506 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2378 : _GEN_1354; // @[dcache.scala 168:42]
  wire  _GEN_2507 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2379 : _GEN_1355; // @[dcache.scala 168:42]
  wire  _GEN_2508 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2380 : _GEN_1356; // @[dcache.scala 168:42]
  wire  _GEN_2509 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2381 : _GEN_1357; // @[dcache.scala 168:42]
  wire  _GEN_2510 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2382 : _GEN_1358; // @[dcache.scala 168:42]
  wire  _GEN_2511 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2383 : _GEN_1359; // @[dcache.scala 168:42]
  wire  _GEN_2512 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2384 : _GEN_1360; // @[dcache.scala 168:42]
  wire  _GEN_2513 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2385 : _GEN_1361; // @[dcache.scala 168:42]
  wire  _GEN_2514 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2386 : _GEN_1362; // @[dcache.scala 168:42]
  wire  _GEN_2515 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2387 : _GEN_1363; // @[dcache.scala 168:42]
  wire  _GEN_2516 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2388 : _GEN_1364; // @[dcache.scala 168:42]
  wire  _GEN_2517 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2389 : _GEN_1365; // @[dcache.scala 168:42]
  wire  _GEN_2518 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2390 : _GEN_1366; // @[dcache.scala 168:42]
  wire  _GEN_2519 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2391 : _GEN_1367; // @[dcache.scala 168:42]
  wire  _GEN_2520 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2392 : _GEN_1368; // @[dcache.scala 168:42]
  wire  _GEN_2521 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2393 : _GEN_1369; // @[dcache.scala 168:42]
  wire  _GEN_2522 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2394 : _GEN_1370; // @[dcache.scala 168:42]
  wire  _GEN_2523 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2395 : _GEN_1371; // @[dcache.scala 168:42]
  wire  _GEN_2524 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2396 : _GEN_1372; // @[dcache.scala 168:42]
  wire  _GEN_2525 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2397 : _GEN_1373; // @[dcache.scala 168:42]
  wire  _GEN_2526 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2398 : _GEN_1374; // @[dcache.scala 168:42]
  wire  _GEN_2527 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2399 : _GEN_1375; // @[dcache.scala 168:42]
  wire  _GEN_2528 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2400 : _GEN_1376; // @[dcache.scala 168:42]
  wire  _GEN_2529 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2401 : _GEN_1377; // @[dcache.scala 168:42]
  wire  _GEN_2530 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2402 : _GEN_1378; // @[dcache.scala 168:42]
  wire  _GEN_2531 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2403 : _GEN_1379; // @[dcache.scala 168:42]
  wire  _GEN_2532 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2404 : _GEN_1380; // @[dcache.scala 168:42]
  wire  _GEN_2533 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2405 : _GEN_1381; // @[dcache.scala 168:42]
  wire  _GEN_2534 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2406 : _GEN_1382; // @[dcache.scala 168:42]
  wire  _GEN_2535 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2407 : _GEN_1383; // @[dcache.scala 168:42]
  wire  _GEN_2536 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2408 : _GEN_1384; // @[dcache.scala 168:42]
  wire  _GEN_2537 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2409 : _GEN_1385; // @[dcache.scala 168:42]
  wire  _GEN_2538 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2410 : _GEN_1386; // @[dcache.scala 168:42]
  wire  _GEN_2539 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2411 : _GEN_1387; // @[dcache.scala 168:42]
  wire  _GEN_2540 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2412 : _GEN_1388; // @[dcache.scala 168:42]
  wire  _GEN_2541 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2413 : _GEN_1389; // @[dcache.scala 168:42]
  wire  _GEN_2542 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2414 : _GEN_1390; // @[dcache.scala 168:42]
  wire  _GEN_2543 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2415 : _GEN_1391; // @[dcache.scala 168:42]
  wire  _GEN_2544 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2416 : _GEN_1392; // @[dcache.scala 168:42]
  wire  _GEN_2545 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2417 : _GEN_1393; // @[dcache.scala 168:42]
  wire  _GEN_2546 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2418 : _GEN_1394; // @[dcache.scala 168:42]
  wire  _GEN_2547 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2419 : _GEN_1395; // @[dcache.scala 168:42]
  wire  _GEN_2548 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2420 : _GEN_1396; // @[dcache.scala 168:42]
  wire  _GEN_2549 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2421 : _GEN_1397; // @[dcache.scala 168:42]
  wire  _GEN_2550 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2422 : _GEN_1398; // @[dcache.scala 168:42]
  wire  _GEN_2551 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2423 : _GEN_1399; // @[dcache.scala 168:42]
  wire  _GEN_2552 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2424 : _GEN_1400; // @[dcache.scala 168:42]
  wire  _GEN_2553 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2425 : _GEN_1401; // @[dcache.scala 168:42]
  wire  _GEN_2554 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2426 : _GEN_1402; // @[dcache.scala 168:42]
  wire  _GEN_2555 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2427 : _GEN_1403; // @[dcache.scala 168:42]
  wire  _GEN_2556 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2428 : _GEN_1404; // @[dcache.scala 168:42]
  wire  _GEN_2557 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2429 : _GEN_1405; // @[dcache.scala 168:42]
  wire  _GEN_2558 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2430 : _GEN_1406; // @[dcache.scala 168:42]
  wire  _GEN_2559 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2431 : _GEN_1407; // @[dcache.scala 168:42]
  wire  _GEN_2560 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2432 : _GEN_1408; // @[dcache.scala 168:42]
  wire  _GEN_2561 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2433 : _GEN_1409; // @[dcache.scala 168:42]
  wire  _GEN_2562 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2434 : _GEN_1410; // @[dcache.scala 168:42]
  wire  _GEN_2563 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2435 : _GEN_1411; // @[dcache.scala 168:42]
  wire  _GEN_2564 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2436 : _GEN_1412; // @[dcache.scala 168:42]
  wire  _GEN_2565 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2437 : _GEN_1413; // @[dcache.scala 168:42]
  wire  _GEN_2566 = cpu_mem_Mwout & hit_bank_0 ? _GEN_2438 : _GEN_1414; // @[dcache.scala 168:42]
  wire  _GEN_2567 = _GEN_3336 | _GEN_2055; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2568 = _GEN_3337 | _GEN_2056; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2569 = _GEN_3338 | _GEN_2057; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2570 = _GEN_3339 | _GEN_2058; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2571 = _GEN_3340 | _GEN_2059; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2572 = _GEN_3341 | _GEN_2060; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2573 = _GEN_3342 | _GEN_2061; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2574 = _GEN_3343 | _GEN_2062; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2575 = _GEN_3344 | _GEN_2063; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2576 = _GEN_3345 | _GEN_2064; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2577 = _GEN_3346 | _GEN_2065; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2578 = _GEN_3347 | _GEN_2066; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2579 = _GEN_3348 | _GEN_2067; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2580 = _GEN_3349 | _GEN_2068; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2581 = _GEN_3350 | _GEN_2069; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2582 = _GEN_3351 | _GEN_2070; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2583 = _GEN_3352 | _GEN_2071; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2584 = _GEN_3353 | _GEN_2072; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2585 = _GEN_3354 | _GEN_2073; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2586 = _GEN_3355 | _GEN_2074; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2587 = _GEN_3356 | _GEN_2075; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2588 = _GEN_3357 | _GEN_2076; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2589 = _GEN_3358 | _GEN_2077; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2590 = _GEN_3359 | _GEN_2078; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2591 = _GEN_3360 | _GEN_2079; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2592 = _GEN_3361 | _GEN_2080; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2593 = _GEN_3362 | _GEN_2081; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2594 = _GEN_3363 | _GEN_2082; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2595 = _GEN_3364 | _GEN_2083; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2596 = _GEN_3365 | _GEN_2084; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2597 = _GEN_3366 | _GEN_2085; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2598 = _GEN_3367 | _GEN_2086; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2599 = _GEN_3368 | _GEN_2087; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2600 = _GEN_3369 | _GEN_2088; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2601 = _GEN_3370 | _GEN_2089; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2602 = _GEN_3371 | _GEN_2090; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2603 = _GEN_3372 | _GEN_2091; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2604 = _GEN_3373 | _GEN_2092; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2605 = _GEN_3374 | _GEN_2093; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2606 = _GEN_3375 | _GEN_2094; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2607 = _GEN_3376 | _GEN_2095; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2608 = _GEN_3377 | _GEN_2096; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2609 = _GEN_3378 | _GEN_2097; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2610 = _GEN_3379 | _GEN_2098; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2611 = _GEN_3380 | _GEN_2099; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2612 = _GEN_3381 | _GEN_2100; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2613 = _GEN_3382 | _GEN_2101; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2614 = _GEN_3383 | _GEN_2102; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2615 = _GEN_3384 | _GEN_2103; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2616 = _GEN_3385 | _GEN_2104; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2617 = _GEN_3386 | _GEN_2105; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2618 = _GEN_3387 | _GEN_2106; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2619 = _GEN_3388 | _GEN_2107; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2620 = _GEN_3389 | _GEN_2108; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2621 = _GEN_3390 | _GEN_2109; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2622 = _GEN_3391 | _GEN_2110; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2623 = _GEN_3392 | _GEN_2111; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2624 = _GEN_3393 | _GEN_2112; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2625 = _GEN_3394 | _GEN_2113; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2626 = _GEN_3395 | _GEN_2114; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2627 = _GEN_3396 | _GEN_2115; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2628 = _GEN_3397 | _GEN_2116; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2629 = _GEN_3398 | _GEN_2117; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2630 = _GEN_3399 | _GEN_2118; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2631 = _GEN_3400 | _GEN_2119; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2632 = _GEN_3401 | _GEN_2120; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2633 = _GEN_3402 | _GEN_2121; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2634 = _GEN_3403 | _GEN_2122; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2635 = _GEN_3404 | _GEN_2123; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2636 = _GEN_3405 | _GEN_2124; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2637 = _GEN_3406 | _GEN_2125; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2638 = _GEN_3407 | _GEN_2126; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2639 = _GEN_3408 | _GEN_2127; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2640 = _GEN_3409 | _GEN_2128; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2641 = _GEN_3410 | _GEN_2129; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2642 = _GEN_3411 | _GEN_2130; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2643 = _GEN_3412 | _GEN_2131; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2644 = _GEN_3413 | _GEN_2132; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2645 = _GEN_3414 | _GEN_2133; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2646 = _GEN_3415 | _GEN_2134; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2647 = _GEN_3416 | _GEN_2135; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2648 = _GEN_3417 | _GEN_2136; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2649 = _GEN_3418 | _GEN_2137; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2650 = _GEN_3419 | _GEN_2138; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2651 = _GEN_3420 | _GEN_2139; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2652 = _GEN_3421 | _GEN_2140; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2653 = _GEN_3422 | _GEN_2141; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2654 = _GEN_3423 | _GEN_2142; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2655 = _GEN_3424 | _GEN_2143; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2656 = _GEN_3425 | _GEN_2144; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2657 = _GEN_3426 | _GEN_2145; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2658 = _GEN_3427 | _GEN_2146; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2659 = _GEN_3428 | _GEN_2147; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2660 = _GEN_3429 | _GEN_2148; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2661 = _GEN_3430 | _GEN_2149; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2662 = _GEN_3431 | _GEN_2150; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2663 = _GEN_3432 | _GEN_2151; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2664 = _GEN_3433 | _GEN_2152; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2665 = _GEN_3434 | _GEN_2153; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2666 = _GEN_3435 | _GEN_2154; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2667 = _GEN_3436 | _GEN_2155; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2668 = _GEN_3437 | _GEN_2156; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2669 = _GEN_3438 | _GEN_2157; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2670 = _GEN_3439 | _GEN_2158; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2671 = _GEN_3440 | _GEN_2159; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2672 = _GEN_3441 | _GEN_2160; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2673 = _GEN_3442 | _GEN_2161; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2674 = _GEN_3443 | _GEN_2162; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2675 = _GEN_3444 | _GEN_2163; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2676 = _GEN_3445 | _GEN_2164; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2677 = _GEN_3446 | _GEN_2165; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2678 = _GEN_3447 | _GEN_2166; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2679 = _GEN_3448 | _GEN_2167; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2680 = _GEN_3449 | _GEN_2168; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2681 = _GEN_3450 | _GEN_2169; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2682 = _GEN_3451 | _GEN_2170; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2683 = _GEN_3452 | _GEN_2171; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2684 = _GEN_3453 | _GEN_2172; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2685 = _GEN_3454 | _GEN_2173; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2686 = _GEN_3455 | _GEN_2174; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2687 = _GEN_3456 | _GEN_2175; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2688 = _GEN_3457 | _GEN_2176; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2689 = _GEN_3458 | _GEN_2177; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2690 = _GEN_3459 | _GEN_2178; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2691 = _GEN_3460 | _GEN_2179; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2692 = _GEN_3461 | _GEN_2180; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2693 = _GEN_3462 | _GEN_2181; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2694 = _GEN_3463 | _GEN_2182; // @[dcache.scala 172:{19,19}]
  wire  _GEN_2695 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2567 : _GEN_2055; // @[dcache.scala 171:42]
  wire  _GEN_2696 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2568 : _GEN_2056; // @[dcache.scala 171:42]
  wire  _GEN_2697 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2569 : _GEN_2057; // @[dcache.scala 171:42]
  wire  _GEN_2698 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2570 : _GEN_2058; // @[dcache.scala 171:42]
  wire  _GEN_2699 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2571 : _GEN_2059; // @[dcache.scala 171:42]
  wire  _GEN_2700 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2572 : _GEN_2060; // @[dcache.scala 171:42]
  wire  _GEN_2701 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2573 : _GEN_2061; // @[dcache.scala 171:42]
  wire  _GEN_2702 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2574 : _GEN_2062; // @[dcache.scala 171:42]
  wire  _GEN_2703 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2575 : _GEN_2063; // @[dcache.scala 171:42]
  wire  _GEN_2704 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2576 : _GEN_2064; // @[dcache.scala 171:42]
  wire  _GEN_2705 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2577 : _GEN_2065; // @[dcache.scala 171:42]
  wire  _GEN_2706 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2578 : _GEN_2066; // @[dcache.scala 171:42]
  wire  _GEN_2707 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2579 : _GEN_2067; // @[dcache.scala 171:42]
  wire  _GEN_2708 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2580 : _GEN_2068; // @[dcache.scala 171:42]
  wire  _GEN_2709 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2581 : _GEN_2069; // @[dcache.scala 171:42]
  wire  _GEN_2710 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2582 : _GEN_2070; // @[dcache.scala 171:42]
  wire  _GEN_2711 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2583 : _GEN_2071; // @[dcache.scala 171:42]
  wire  _GEN_2712 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2584 : _GEN_2072; // @[dcache.scala 171:42]
  wire  _GEN_2713 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2585 : _GEN_2073; // @[dcache.scala 171:42]
  wire  _GEN_2714 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2586 : _GEN_2074; // @[dcache.scala 171:42]
  wire  _GEN_2715 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2587 : _GEN_2075; // @[dcache.scala 171:42]
  wire  _GEN_2716 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2588 : _GEN_2076; // @[dcache.scala 171:42]
  wire  _GEN_2717 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2589 : _GEN_2077; // @[dcache.scala 171:42]
  wire  _GEN_2718 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2590 : _GEN_2078; // @[dcache.scala 171:42]
  wire  _GEN_2719 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2591 : _GEN_2079; // @[dcache.scala 171:42]
  wire  _GEN_2720 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2592 : _GEN_2080; // @[dcache.scala 171:42]
  wire  _GEN_2721 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2593 : _GEN_2081; // @[dcache.scala 171:42]
  wire  _GEN_2722 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2594 : _GEN_2082; // @[dcache.scala 171:42]
  wire  _GEN_2723 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2595 : _GEN_2083; // @[dcache.scala 171:42]
  wire  _GEN_2724 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2596 : _GEN_2084; // @[dcache.scala 171:42]
  wire  _GEN_2725 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2597 : _GEN_2085; // @[dcache.scala 171:42]
  wire  _GEN_2726 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2598 : _GEN_2086; // @[dcache.scala 171:42]
  wire  _GEN_2727 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2599 : _GEN_2087; // @[dcache.scala 171:42]
  wire  _GEN_2728 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2600 : _GEN_2088; // @[dcache.scala 171:42]
  wire  _GEN_2729 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2601 : _GEN_2089; // @[dcache.scala 171:42]
  wire  _GEN_2730 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2602 : _GEN_2090; // @[dcache.scala 171:42]
  wire  _GEN_2731 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2603 : _GEN_2091; // @[dcache.scala 171:42]
  wire  _GEN_2732 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2604 : _GEN_2092; // @[dcache.scala 171:42]
  wire  _GEN_2733 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2605 : _GEN_2093; // @[dcache.scala 171:42]
  wire  _GEN_2734 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2606 : _GEN_2094; // @[dcache.scala 171:42]
  wire  _GEN_2735 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2607 : _GEN_2095; // @[dcache.scala 171:42]
  wire  _GEN_2736 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2608 : _GEN_2096; // @[dcache.scala 171:42]
  wire  _GEN_2737 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2609 : _GEN_2097; // @[dcache.scala 171:42]
  wire  _GEN_2738 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2610 : _GEN_2098; // @[dcache.scala 171:42]
  wire  _GEN_2739 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2611 : _GEN_2099; // @[dcache.scala 171:42]
  wire  _GEN_2740 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2612 : _GEN_2100; // @[dcache.scala 171:42]
  wire  _GEN_2741 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2613 : _GEN_2101; // @[dcache.scala 171:42]
  wire  _GEN_2742 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2614 : _GEN_2102; // @[dcache.scala 171:42]
  wire  _GEN_2743 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2615 : _GEN_2103; // @[dcache.scala 171:42]
  wire  _GEN_2744 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2616 : _GEN_2104; // @[dcache.scala 171:42]
  wire  _GEN_2745 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2617 : _GEN_2105; // @[dcache.scala 171:42]
  wire  _GEN_2746 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2618 : _GEN_2106; // @[dcache.scala 171:42]
  wire  _GEN_2747 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2619 : _GEN_2107; // @[dcache.scala 171:42]
  wire  _GEN_2748 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2620 : _GEN_2108; // @[dcache.scala 171:42]
  wire  _GEN_2749 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2621 : _GEN_2109; // @[dcache.scala 171:42]
  wire  _GEN_2750 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2622 : _GEN_2110; // @[dcache.scala 171:42]
  wire  _GEN_2751 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2623 : _GEN_2111; // @[dcache.scala 171:42]
  wire  _GEN_2752 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2624 : _GEN_2112; // @[dcache.scala 171:42]
  wire  _GEN_2753 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2625 : _GEN_2113; // @[dcache.scala 171:42]
  wire  _GEN_2754 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2626 : _GEN_2114; // @[dcache.scala 171:42]
  wire  _GEN_2755 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2627 : _GEN_2115; // @[dcache.scala 171:42]
  wire  _GEN_2756 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2628 : _GEN_2116; // @[dcache.scala 171:42]
  wire  _GEN_2757 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2629 : _GEN_2117; // @[dcache.scala 171:42]
  wire  _GEN_2758 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2630 : _GEN_2118; // @[dcache.scala 171:42]
  wire  _GEN_2759 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2631 : _GEN_2119; // @[dcache.scala 171:42]
  wire  _GEN_2760 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2632 : _GEN_2120; // @[dcache.scala 171:42]
  wire  _GEN_2761 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2633 : _GEN_2121; // @[dcache.scala 171:42]
  wire  _GEN_2762 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2634 : _GEN_2122; // @[dcache.scala 171:42]
  wire  _GEN_2763 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2635 : _GEN_2123; // @[dcache.scala 171:42]
  wire  _GEN_2764 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2636 : _GEN_2124; // @[dcache.scala 171:42]
  wire  _GEN_2765 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2637 : _GEN_2125; // @[dcache.scala 171:42]
  wire  _GEN_2766 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2638 : _GEN_2126; // @[dcache.scala 171:42]
  wire  _GEN_2767 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2639 : _GEN_2127; // @[dcache.scala 171:42]
  wire  _GEN_2768 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2640 : _GEN_2128; // @[dcache.scala 171:42]
  wire  _GEN_2769 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2641 : _GEN_2129; // @[dcache.scala 171:42]
  wire  _GEN_2770 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2642 : _GEN_2130; // @[dcache.scala 171:42]
  wire  _GEN_2771 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2643 : _GEN_2131; // @[dcache.scala 171:42]
  wire  _GEN_2772 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2644 : _GEN_2132; // @[dcache.scala 171:42]
  wire  _GEN_2773 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2645 : _GEN_2133; // @[dcache.scala 171:42]
  wire  _GEN_2774 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2646 : _GEN_2134; // @[dcache.scala 171:42]
  wire  _GEN_2775 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2647 : _GEN_2135; // @[dcache.scala 171:42]
  wire  _GEN_2776 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2648 : _GEN_2136; // @[dcache.scala 171:42]
  wire  _GEN_2777 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2649 : _GEN_2137; // @[dcache.scala 171:42]
  wire  _GEN_2778 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2650 : _GEN_2138; // @[dcache.scala 171:42]
  wire  _GEN_2779 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2651 : _GEN_2139; // @[dcache.scala 171:42]
  wire  _GEN_2780 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2652 : _GEN_2140; // @[dcache.scala 171:42]
  wire  _GEN_2781 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2653 : _GEN_2141; // @[dcache.scala 171:42]
  wire  _GEN_2782 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2654 : _GEN_2142; // @[dcache.scala 171:42]
  wire  _GEN_2783 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2655 : _GEN_2143; // @[dcache.scala 171:42]
  wire  _GEN_2784 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2656 : _GEN_2144; // @[dcache.scala 171:42]
  wire  _GEN_2785 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2657 : _GEN_2145; // @[dcache.scala 171:42]
  wire  _GEN_2786 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2658 : _GEN_2146; // @[dcache.scala 171:42]
  wire  _GEN_2787 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2659 : _GEN_2147; // @[dcache.scala 171:42]
  wire  _GEN_2788 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2660 : _GEN_2148; // @[dcache.scala 171:42]
  wire  _GEN_2789 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2661 : _GEN_2149; // @[dcache.scala 171:42]
  wire  _GEN_2790 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2662 : _GEN_2150; // @[dcache.scala 171:42]
  wire  _GEN_2791 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2663 : _GEN_2151; // @[dcache.scala 171:42]
  wire  _GEN_2792 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2664 : _GEN_2152; // @[dcache.scala 171:42]
  wire  _GEN_2793 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2665 : _GEN_2153; // @[dcache.scala 171:42]
  wire  _GEN_2794 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2666 : _GEN_2154; // @[dcache.scala 171:42]
  wire  _GEN_2795 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2667 : _GEN_2155; // @[dcache.scala 171:42]
  wire  _GEN_2796 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2668 : _GEN_2156; // @[dcache.scala 171:42]
  wire  _GEN_2797 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2669 : _GEN_2157; // @[dcache.scala 171:42]
  wire  _GEN_2798 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2670 : _GEN_2158; // @[dcache.scala 171:42]
  wire  _GEN_2799 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2671 : _GEN_2159; // @[dcache.scala 171:42]
  wire  _GEN_2800 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2672 : _GEN_2160; // @[dcache.scala 171:42]
  wire  _GEN_2801 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2673 : _GEN_2161; // @[dcache.scala 171:42]
  wire  _GEN_2802 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2674 : _GEN_2162; // @[dcache.scala 171:42]
  wire  _GEN_2803 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2675 : _GEN_2163; // @[dcache.scala 171:42]
  wire  _GEN_2804 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2676 : _GEN_2164; // @[dcache.scala 171:42]
  wire  _GEN_2805 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2677 : _GEN_2165; // @[dcache.scala 171:42]
  wire  _GEN_2806 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2678 : _GEN_2166; // @[dcache.scala 171:42]
  wire  _GEN_2807 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2679 : _GEN_2167; // @[dcache.scala 171:42]
  wire  _GEN_2808 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2680 : _GEN_2168; // @[dcache.scala 171:42]
  wire  _GEN_2809 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2681 : _GEN_2169; // @[dcache.scala 171:42]
  wire  _GEN_2810 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2682 : _GEN_2170; // @[dcache.scala 171:42]
  wire  _GEN_2811 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2683 : _GEN_2171; // @[dcache.scala 171:42]
  wire  _GEN_2812 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2684 : _GEN_2172; // @[dcache.scala 171:42]
  wire  _GEN_2813 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2685 : _GEN_2173; // @[dcache.scala 171:42]
  wire  _GEN_2814 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2686 : _GEN_2174; // @[dcache.scala 171:42]
  wire  _GEN_2815 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2687 : _GEN_2175; // @[dcache.scala 171:42]
  wire  _GEN_2816 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2688 : _GEN_2176; // @[dcache.scala 171:42]
  wire  _GEN_2817 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2689 : _GEN_2177; // @[dcache.scala 171:42]
  wire  _GEN_2818 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2690 : _GEN_2178; // @[dcache.scala 171:42]
  wire  _GEN_2819 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2691 : _GEN_2179; // @[dcache.scala 171:42]
  wire  _GEN_2820 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2692 : _GEN_2180; // @[dcache.scala 171:42]
  wire  _GEN_2821 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2693 : _GEN_2181; // @[dcache.scala 171:42]
  wire  _GEN_2822 = cpu_mem_Mwout & hit_bank_1 ? _GEN_2694 : _GEN_2182; // @[dcache.scala 171:42]
  wire  _next_write_state_T = write_state == 3'h0; // @[dcache.scala 196:18]
  wire  _next_write_state_T_1 = write_state == 3'h2; // @[dcache.scala 197:18]
  wire  _next_write_state_T_2 = write_state == 3'h2 & io_mem_master_writeAddr_ready; // @[dcache.scala 197:33]
  wire  _next_write_state_T_3 = write_state == 3'h3; // @[dcache.scala 198:18]
  wire  _next_write_state_T_4 = write_state == 3'h3 & io_mem_master_writeData_ready; // @[dcache.scala 198:33]
  wire  _next_write_state_T_6 = write_state == 3'h4 & io_mem_master_writeResp_valid; // @[dcache.scala 199:33]
  wire  _next_write_state_T_9 = _io_cpu_mem_data_valid_T_6 & _io_cpu_mem_data_valid_T; // @[dcache.scala 200:30]
  wire  _next_write_state_T_14 = _io_cpu_mem_data_valid_T_6 & _next_state_T_2 & cpu_mem_Mwout; // @[dcache.scala 201:38]
  wire  _next_write_state_T_16 = _io_cpu_mem_data_valid_T_6 & should_write_back; // @[dcache.scala 202:30]
  wire [2:0] _next_write_state_T_17 = _next_write_state_T_16 ? 3'h2 : write_state; // @[Mux.scala 101:16]
  wire [2:0] _next_write_state_T_18 = _next_write_state_T_14 ? 3'h2 : _next_write_state_T_17; // @[Mux.scala 101:16]
  wire [2:0] _next_write_state_T_19 = _next_write_state_T_9 ? 3'h1 : _next_write_state_T_18; // @[Mux.scala 101:16]
  wire [2:0] _next_write_state_T_20 = _next_write_state_T_6 ? 3'h1 : _next_write_state_T_19; // @[Mux.scala 101:16]
  wire [2:0] _next_write_state_T_21 = _next_write_state_T_4 ? 3'h4 : _next_write_state_T_20; // @[Mux.scala 101:16]
  wire [2:0] _next_write_state_T_22 = _next_write_state_T_2 ? 3'h3 : _next_write_state_T_21; // @[Mux.scala 101:16]
  wire [2:0] next_write_state = _next_write_state_T ? 3'h1 : _next_write_state_T_22; // @[Mux.scala 101:16]
  wire  _T_23 = _write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1; // @[dcache.scala 174:51]
  wire  _GEN_2823 = _GEN_3336 | _GEN_2439; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2824 = _GEN_3337 | _GEN_2440; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2825 = _GEN_3338 | _GEN_2441; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2826 = _GEN_3339 | _GEN_2442; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2827 = _GEN_3340 | _GEN_2443; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2828 = _GEN_3341 | _GEN_2444; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2829 = _GEN_3342 | _GEN_2445; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2830 = _GEN_3343 | _GEN_2446; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2831 = _GEN_3344 | _GEN_2447; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2832 = _GEN_3345 | _GEN_2448; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2833 = _GEN_3346 | _GEN_2449; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2834 = _GEN_3347 | _GEN_2450; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2835 = _GEN_3348 | _GEN_2451; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2836 = _GEN_3349 | _GEN_2452; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2837 = _GEN_3350 | _GEN_2453; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2838 = _GEN_3351 | _GEN_2454; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2839 = _GEN_3352 | _GEN_2455; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2840 = _GEN_3353 | _GEN_2456; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2841 = _GEN_3354 | _GEN_2457; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2842 = _GEN_3355 | _GEN_2458; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2843 = _GEN_3356 | _GEN_2459; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2844 = _GEN_3357 | _GEN_2460; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2845 = _GEN_3358 | _GEN_2461; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2846 = _GEN_3359 | _GEN_2462; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2847 = _GEN_3360 | _GEN_2463; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2848 = _GEN_3361 | _GEN_2464; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2849 = _GEN_3362 | _GEN_2465; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2850 = _GEN_3363 | _GEN_2466; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2851 = _GEN_3364 | _GEN_2467; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2852 = _GEN_3365 | _GEN_2468; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2853 = _GEN_3366 | _GEN_2469; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2854 = _GEN_3367 | _GEN_2470; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2855 = _GEN_3368 | _GEN_2471; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2856 = _GEN_3369 | _GEN_2472; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2857 = _GEN_3370 | _GEN_2473; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2858 = _GEN_3371 | _GEN_2474; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2859 = _GEN_3372 | _GEN_2475; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2860 = _GEN_3373 | _GEN_2476; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2861 = _GEN_3374 | _GEN_2477; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2862 = _GEN_3375 | _GEN_2478; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2863 = _GEN_3376 | _GEN_2479; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2864 = _GEN_3377 | _GEN_2480; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2865 = _GEN_3378 | _GEN_2481; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2866 = _GEN_3379 | _GEN_2482; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2867 = _GEN_3380 | _GEN_2483; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2868 = _GEN_3381 | _GEN_2484; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2869 = _GEN_3382 | _GEN_2485; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2870 = _GEN_3383 | _GEN_2486; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2871 = _GEN_3384 | _GEN_2487; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2872 = _GEN_3385 | _GEN_2488; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2873 = _GEN_3386 | _GEN_2489; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2874 = _GEN_3387 | _GEN_2490; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2875 = _GEN_3388 | _GEN_2491; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2876 = _GEN_3389 | _GEN_2492; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2877 = _GEN_3390 | _GEN_2493; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2878 = _GEN_3391 | _GEN_2494; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2879 = _GEN_3392 | _GEN_2495; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2880 = _GEN_3393 | _GEN_2496; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2881 = _GEN_3394 | _GEN_2497; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2882 = _GEN_3395 | _GEN_2498; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2883 = _GEN_3396 | _GEN_2499; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2884 = _GEN_3397 | _GEN_2500; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2885 = _GEN_3398 | _GEN_2501; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2886 = _GEN_3399 | _GEN_2502; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2887 = _GEN_3400 | _GEN_2503; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2888 = _GEN_3401 | _GEN_2504; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2889 = _GEN_3402 | _GEN_2505; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2890 = _GEN_3403 | _GEN_2506; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2891 = _GEN_3404 | _GEN_2507; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2892 = _GEN_3405 | _GEN_2508; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2893 = _GEN_3406 | _GEN_2509; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2894 = _GEN_3407 | _GEN_2510; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2895 = _GEN_3408 | _GEN_2511; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2896 = _GEN_3409 | _GEN_2512; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2897 = _GEN_3410 | _GEN_2513; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2898 = _GEN_3411 | _GEN_2514; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2899 = _GEN_3412 | _GEN_2515; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2900 = _GEN_3413 | _GEN_2516; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2901 = _GEN_3414 | _GEN_2517; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2902 = _GEN_3415 | _GEN_2518; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2903 = _GEN_3416 | _GEN_2519; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2904 = _GEN_3417 | _GEN_2520; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2905 = _GEN_3418 | _GEN_2521; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2906 = _GEN_3419 | _GEN_2522; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2907 = _GEN_3420 | _GEN_2523; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2908 = _GEN_3421 | _GEN_2524; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2909 = _GEN_3422 | _GEN_2525; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2910 = _GEN_3423 | _GEN_2526; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2911 = _GEN_3424 | _GEN_2527; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2912 = _GEN_3425 | _GEN_2528; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2913 = _GEN_3426 | _GEN_2529; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2914 = _GEN_3427 | _GEN_2530; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2915 = _GEN_3428 | _GEN_2531; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2916 = _GEN_3429 | _GEN_2532; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2917 = _GEN_3430 | _GEN_2533; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2918 = _GEN_3431 | _GEN_2534; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2919 = _GEN_3432 | _GEN_2535; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2920 = _GEN_3433 | _GEN_2536; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2921 = _GEN_3434 | _GEN_2537; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2922 = _GEN_3435 | _GEN_2538; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2923 = _GEN_3436 | _GEN_2539; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2924 = _GEN_3437 | _GEN_2540; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2925 = _GEN_3438 | _GEN_2541; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2926 = _GEN_3439 | _GEN_2542; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2927 = _GEN_3440 | _GEN_2543; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2928 = _GEN_3441 | _GEN_2544; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2929 = _GEN_3442 | _GEN_2545; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2930 = _GEN_3443 | _GEN_2546; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2931 = _GEN_3444 | _GEN_2547; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2932 = _GEN_3445 | _GEN_2548; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2933 = _GEN_3446 | _GEN_2549; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2934 = _GEN_3447 | _GEN_2550; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2935 = _GEN_3448 | _GEN_2551; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2936 = _GEN_3449 | _GEN_2552; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2937 = _GEN_3450 | _GEN_2553; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2938 = _GEN_3451 | _GEN_2554; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2939 = _GEN_3452 | _GEN_2555; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2940 = _GEN_3453 | _GEN_2556; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2941 = _GEN_3454 | _GEN_2557; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2942 = _GEN_3455 | _GEN_2558; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2943 = _GEN_3456 | _GEN_2559; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2944 = _GEN_3457 | _GEN_2560; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2945 = _GEN_3458 | _GEN_2561; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2946 = _GEN_3459 | _GEN_2562; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2947 = _GEN_3460 | _GEN_2563; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2948 = _GEN_3461 | _GEN_2564; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2949 = _GEN_3462 | _GEN_2565; // @[dcache.scala 175:{19,19}]
  wire  _GEN_2950 = _GEN_3463 | _GEN_2566; // @[dcache.scala 175:{19,19}]
  wire  _GEN_3079 = _GEN_3336 | _GEN_2695; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3080 = _GEN_3337 | _GEN_2696; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3081 = _GEN_3338 | _GEN_2697; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3082 = _GEN_3339 | _GEN_2698; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3083 = _GEN_3340 | _GEN_2699; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3084 = _GEN_3341 | _GEN_2700; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3085 = _GEN_3342 | _GEN_2701; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3086 = _GEN_3343 | _GEN_2702; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3087 = _GEN_3344 | _GEN_2703; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3088 = _GEN_3345 | _GEN_2704; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3089 = _GEN_3346 | _GEN_2705; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3090 = _GEN_3347 | _GEN_2706; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3091 = _GEN_3348 | _GEN_2707; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3092 = _GEN_3349 | _GEN_2708; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3093 = _GEN_3350 | _GEN_2709; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3094 = _GEN_3351 | _GEN_2710; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3095 = _GEN_3352 | _GEN_2711; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3096 = _GEN_3353 | _GEN_2712; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3097 = _GEN_3354 | _GEN_2713; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3098 = _GEN_3355 | _GEN_2714; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3099 = _GEN_3356 | _GEN_2715; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3100 = _GEN_3357 | _GEN_2716; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3101 = _GEN_3358 | _GEN_2717; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3102 = _GEN_3359 | _GEN_2718; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3103 = _GEN_3360 | _GEN_2719; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3104 = _GEN_3361 | _GEN_2720; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3105 = _GEN_3362 | _GEN_2721; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3106 = _GEN_3363 | _GEN_2722; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3107 = _GEN_3364 | _GEN_2723; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3108 = _GEN_3365 | _GEN_2724; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3109 = _GEN_3366 | _GEN_2725; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3110 = _GEN_3367 | _GEN_2726; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3111 = _GEN_3368 | _GEN_2727; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3112 = _GEN_3369 | _GEN_2728; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3113 = _GEN_3370 | _GEN_2729; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3114 = _GEN_3371 | _GEN_2730; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3115 = _GEN_3372 | _GEN_2731; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3116 = _GEN_3373 | _GEN_2732; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3117 = _GEN_3374 | _GEN_2733; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3118 = _GEN_3375 | _GEN_2734; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3119 = _GEN_3376 | _GEN_2735; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3120 = _GEN_3377 | _GEN_2736; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3121 = _GEN_3378 | _GEN_2737; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3122 = _GEN_3379 | _GEN_2738; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3123 = _GEN_3380 | _GEN_2739; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3124 = _GEN_3381 | _GEN_2740; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3125 = _GEN_3382 | _GEN_2741; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3126 = _GEN_3383 | _GEN_2742; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3127 = _GEN_3384 | _GEN_2743; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3128 = _GEN_3385 | _GEN_2744; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3129 = _GEN_3386 | _GEN_2745; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3130 = _GEN_3387 | _GEN_2746; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3131 = _GEN_3388 | _GEN_2747; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3132 = _GEN_3389 | _GEN_2748; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3133 = _GEN_3390 | _GEN_2749; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3134 = _GEN_3391 | _GEN_2750; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3135 = _GEN_3392 | _GEN_2751; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3136 = _GEN_3393 | _GEN_2752; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3137 = _GEN_3394 | _GEN_2753; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3138 = _GEN_3395 | _GEN_2754; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3139 = _GEN_3396 | _GEN_2755; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3140 = _GEN_3397 | _GEN_2756; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3141 = _GEN_3398 | _GEN_2757; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3142 = _GEN_3399 | _GEN_2758; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3143 = _GEN_3400 | _GEN_2759; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3144 = _GEN_3401 | _GEN_2760; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3145 = _GEN_3402 | _GEN_2761; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3146 = _GEN_3403 | _GEN_2762; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3147 = _GEN_3404 | _GEN_2763; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3148 = _GEN_3405 | _GEN_2764; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3149 = _GEN_3406 | _GEN_2765; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3150 = _GEN_3407 | _GEN_2766; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3151 = _GEN_3408 | _GEN_2767; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3152 = _GEN_3409 | _GEN_2768; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3153 = _GEN_3410 | _GEN_2769; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3154 = _GEN_3411 | _GEN_2770; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3155 = _GEN_3412 | _GEN_2771; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3156 = _GEN_3413 | _GEN_2772; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3157 = _GEN_3414 | _GEN_2773; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3158 = _GEN_3415 | _GEN_2774; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3159 = _GEN_3416 | _GEN_2775; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3160 = _GEN_3417 | _GEN_2776; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3161 = _GEN_3418 | _GEN_2777; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3162 = _GEN_3419 | _GEN_2778; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3163 = _GEN_3420 | _GEN_2779; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3164 = _GEN_3421 | _GEN_2780; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3165 = _GEN_3422 | _GEN_2781; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3166 = _GEN_3423 | _GEN_2782; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3167 = _GEN_3424 | _GEN_2783; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3168 = _GEN_3425 | _GEN_2784; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3169 = _GEN_3426 | _GEN_2785; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3170 = _GEN_3427 | _GEN_2786; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3171 = _GEN_3428 | _GEN_2787; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3172 = _GEN_3429 | _GEN_2788; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3173 = _GEN_3430 | _GEN_2789; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3174 = _GEN_3431 | _GEN_2790; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3175 = _GEN_3432 | _GEN_2791; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3176 = _GEN_3433 | _GEN_2792; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3177 = _GEN_3434 | _GEN_2793; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3178 = _GEN_3435 | _GEN_2794; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3179 = _GEN_3436 | _GEN_2795; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3180 = _GEN_3437 | _GEN_2796; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3181 = _GEN_3438 | _GEN_2797; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3182 = _GEN_3439 | _GEN_2798; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3183 = _GEN_3440 | _GEN_2799; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3184 = _GEN_3441 | _GEN_2800; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3185 = _GEN_3442 | _GEN_2801; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3186 = _GEN_3443 | _GEN_2802; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3187 = _GEN_3444 | _GEN_2803; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3188 = _GEN_3445 | _GEN_2804; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3189 = _GEN_3446 | _GEN_2805; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3190 = _GEN_3447 | _GEN_2806; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3191 = _GEN_3448 | _GEN_2807; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3192 = _GEN_3449 | _GEN_2808; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3193 = _GEN_3450 | _GEN_2809; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3194 = _GEN_3451 | _GEN_2810; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3195 = _GEN_3452 | _GEN_2811; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3196 = _GEN_3453 | _GEN_2812; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3197 = _GEN_3454 | _GEN_2813; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3198 = _GEN_3455 | _GEN_2814; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3199 = _GEN_3456 | _GEN_2815; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3200 = _GEN_3457 | _GEN_2816; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3201 = _GEN_3458 | _GEN_2817; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3202 = _GEN_3459 | _GEN_2818; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3203 = _GEN_3460 | _GEN_2819; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3204 = _GEN_3461 | _GEN_2820; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3205 = _GEN_3462 | _GEN_2821; // @[dcache.scala 178:{19,19}]
  wire  _GEN_3206 = _GEN_3463 | _GEN_2822; // @[dcache.scala 178:{19,19}]
  wire [63:0] _io_mem_master_writeAddr_bits_addr_T_3 = {_GEN_646,index,4'h0}; // @[Cat.scala 33:92]
  wire [63:0] _io_mem_master_writeAddr_bits_addr_T_4 = {_GEN_774,index,4'h0}; // @[Cat.scala 33:92]
  wire [63:0] _io_mem_master_writeAddr_bits_addr_T_5 = _data_array_0_io_i_wen_T_9 ?
    _io_mem_master_writeAddr_bits_addr_T_3 : _io_mem_master_writeAddr_bits_addr_T_4; // @[dcache.scala 210:60]
  wire [127:0] _io_mem_master_writeData_bits_data_T_2 = victim ? data_array_1_io_o_rdata : data_array_0_io_o_rdata; // @[dcache.scala 212:61]
  Data_Array data_array_0 ( // @[dcache.scala 52:36]
    .clock(data_array_0_clock),
    .reset(data_array_0_reset),
    .io_i_wen(data_array_0_io_i_wen),
    .io_i_wstrb(data_array_0_io_i_wstrb),
    .io_i_addr(data_array_0_io_i_addr),
    .io_i_wdata(data_array_0_io_i_wdata),
    .io_o_rdata(data_array_0_io_o_rdata)
  );
  Data_Array data_array_1 ( // @[dcache.scala 52:36]
    .clock(data_array_1_clock),
    .reset(data_array_1_reset),
    .io_i_wen(data_array_1_io_i_wen),
    .io_i_wstrb(data_array_1_io_i_wstrb),
    .io_i_addr(data_array_1_io_i_addr),
    .io_i_wdata(data_array_1_io_i_wdata),
    .io_o_rdata(data_array_1_io_o_rdata)
  );
  assign io_cpu_mem_data_valid = next_state != 2'h2 & ~new_req & cpu_mem_Men & _write_back_is_finishing_T & write_state
     == 3'h1; // @[dcache.scala 111:94]
  assign io_cpu_mem_addr_ready = state == 2'h1; // @[dcache.scala 112:32]
  assign io_cpu_mem_MdataIn = _io_cpu_mem_MdataIn_T_2[63:0]; // @[dcache.scala 100:20]
  assign io_mem_master_readAddr_valid = _should_write_back_T & _write_back_is_finishing_T & cpu_mem_Men &
    _io_cpu_mem_data_valid_T_6; // @[dcache.scala 205:88]
  assign io_mem_master_readAddr_bits_addr = {cpu_mem_Maddr[63:4],4'h0}; // @[Cat.scala 33:92]
  assign io_mem_master_readData_ready = _should_write_back_T & _io_cpu_mem_data_valid_T_6; // @[dcache.scala 207:51]
  assign io_mem_master_writeAddr_valid = _next_write_state_T_1 | _next_write_state_T_3; // @[dcache.scala 209:62]
  assign io_mem_master_writeAddr_bits_addr = _write_back_is_finishing_T ? _io_mem_master_writeAddr_bits_addr_T_5 :
    cpu_mem_Maddr; // @[dcache.scala 210:41]
  assign io_mem_master_writeData_valid = _next_write_state_T_1 | _next_write_state_T_3; // @[dcache.scala 211:62]
  assign io_mem_master_writeData_bits_data = _write_back_is_finishing_T ? _io_mem_master_writeData_bits_data_T_2 : {{64
    'd0}, cpu_mem_MdataOut}; // @[dcache.scala 212:41]
  assign io_mem_master_writeData_bits_strb = _write_back_is_finishing_T ? 16'hffff : strb; // @[dcache.scala 213:41]
  assign io_mem_master_writeResp_ready = write_state == 3'h4; // @[dcache.scala 214:47]
  assign data_array_0_clock = clock;
  assign data_array_0_reset = reset;
  assign data_array_0_io_i_wen = cpu_mem_Mwout & cpu_mem_Men & hit_bank_0 | _write_back_is_finishing_T &
    _should_write_back_T & _T & ~victim; // @[dcache.scala 152:83]
  assign data_array_0_io_i_wstrb = hit ? strb_aligned : 16'hffff; // @[dcache.scala 153:36]
  assign data_array_0_io_i_addr = cpu_mem_Maddr[10:4]; // @[dcache.scala 115:23]
  assign data_array_0_io_i_wdata = _data_array_0_io_i_wdata_T_4[127:0]; // @[dcache.scala 155:30]
  assign data_array_1_clock = clock;
  assign data_array_1_reset = reset;
  assign data_array_1_io_i_wen = cpu_mem_Mwout & cpu_mem_Men & hit_bank_1 | _write_back_is_finishing_T &
    _should_write_back_T & _T & victim; // @[dcache.scala 152:83]
  assign data_array_1_io_i_wstrb = hit ? strb_aligned : 16'hffff; // @[dcache.scala 153:36]
  assign data_array_1_io_i_addr = cpu_mem_Maddr[10:4]; // @[dcache.scala 115:23]
  assign data_array_1_io_i_wdata = _data_array_0_io_i_wdata_T_4[127:0]; // @[dcache.scala 155:30]
  always @(posedge clock) begin
    if (reset) begin // @[dcache.scala 35:22]
      cpu_mem_Mwout <= 1'h0; // @[dcache.scala 35:22]
    end else if (next_state == 2'h1) begin // @[dcache.scala 88:26]
      cpu_mem_Mwout <= io_cpu_mem_Mwout; // @[dcache.scala 89:11]
    end
    if (reset) begin // @[dcache.scala 35:22]
      cpu_mem_Maddr <= 64'h0; // @[dcache.scala 35:22]
    end else if (next_state == 2'h1) begin // @[dcache.scala 88:26]
      cpu_mem_Maddr <= io_cpu_mem_Maddr; // @[dcache.scala 89:11]
    end
    if (reset) begin // @[dcache.scala 35:22]
      cpu_mem_Men <= 1'h0; // @[dcache.scala 35:22]
    end else if (next_state == 2'h1) begin // @[dcache.scala 88:26]
      cpu_mem_Men <= io_cpu_mem_Men; // @[dcache.scala 89:11]
    end
    if (reset) begin // @[dcache.scala 35:22]
      cpu_mem_Mlen <= 32'h0; // @[dcache.scala 35:22]
    end else if (next_state == 2'h1) begin // @[dcache.scala 88:26]
      cpu_mem_Mlen <= io_cpu_mem_Mlen; // @[dcache.scala 89:11]
    end
    if (reset) begin // @[dcache.scala 35:22]
      cpu_mem_MdataOut <= 64'h0; // @[dcache.scala 35:22]
    end else if (next_state == 2'h1) begin // @[dcache.scala 88:26]
      cpu_mem_MdataOut <= io_cpu_mem_MdataOut; // @[dcache.scala 89:11]
    end
    if (reset) begin // @[dcache.scala 36:23]
      last_req_Mwout <= 1'h0; // @[dcache.scala 36:23]
    end else begin
      last_req_Mwout <= cpu_mem_Mwout; // @[dcache.scala 37:10]
    end
    if (reset) begin // @[dcache.scala 36:23]
      last_req_Maddr <= 64'h0; // @[dcache.scala 36:23]
    end else begin
      last_req_Maddr <= cpu_mem_Maddr; // @[dcache.scala 37:10]
    end
    if (reset) begin // @[dcache.scala 36:23]
      last_req_Men <= 1'h0; // @[dcache.scala 36:23]
    end else begin
      last_req_Men <= cpu_mem_Men; // @[dcache.scala 37:10]
    end
    if (reset) begin // @[dcache.scala 36:23]
      last_req_Mlen <= 32'h0; // @[dcache.scala 36:23]
    end else begin
      last_req_Mlen <= cpu_mem_Mlen; // @[dcache.scala 37:10]
    end
    if (reset) begin // @[dcache.scala 36:23]
      last_req_MdataOut <= 64'h0; // @[dcache.scala 36:23]
    end else begin
      last_req_MdataOut <= cpu_mem_MdataOut; // @[dcache.scala 37:10]
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_0 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h0 == index) begin // @[dcache.scala 161:18]
        tags0_0 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_1 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1 == index) begin // @[dcache.scala 161:18]
        tags0_1 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_2 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2 == index) begin // @[dcache.scala 161:18]
        tags0_2 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_3 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3 == index) begin // @[dcache.scala 161:18]
        tags0_3 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_4 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4 == index) begin // @[dcache.scala 161:18]
        tags0_4 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_5 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5 == index) begin // @[dcache.scala 161:18]
        tags0_5 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_6 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6 == index) begin // @[dcache.scala 161:18]
        tags0_6 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_7 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7 == index) begin // @[dcache.scala 161:18]
        tags0_7 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_8 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h8 == index) begin // @[dcache.scala 161:18]
        tags0_8 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_9 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h9 == index) begin // @[dcache.scala 161:18]
        tags0_9 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_10 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'ha == index) begin // @[dcache.scala 161:18]
        tags0_10 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_11 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'hb == index) begin // @[dcache.scala 161:18]
        tags0_11 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_12 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'hc == index) begin // @[dcache.scala 161:18]
        tags0_12 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_13 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'hd == index) begin // @[dcache.scala 161:18]
        tags0_13 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_14 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'he == index) begin // @[dcache.scala 161:18]
        tags0_14 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_15 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'hf == index) begin // @[dcache.scala 161:18]
        tags0_15 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_16 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h10 == index) begin // @[dcache.scala 161:18]
        tags0_16 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_17 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h11 == index) begin // @[dcache.scala 161:18]
        tags0_17 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_18 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h12 == index) begin // @[dcache.scala 161:18]
        tags0_18 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_19 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h13 == index) begin // @[dcache.scala 161:18]
        tags0_19 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_20 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h14 == index) begin // @[dcache.scala 161:18]
        tags0_20 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_21 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h15 == index) begin // @[dcache.scala 161:18]
        tags0_21 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_22 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h16 == index) begin // @[dcache.scala 161:18]
        tags0_22 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_23 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h17 == index) begin // @[dcache.scala 161:18]
        tags0_23 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_24 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h18 == index) begin // @[dcache.scala 161:18]
        tags0_24 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_25 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h19 == index) begin // @[dcache.scala 161:18]
        tags0_25 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_26 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1a == index) begin // @[dcache.scala 161:18]
        tags0_26 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_27 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1b == index) begin // @[dcache.scala 161:18]
        tags0_27 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_28 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1c == index) begin // @[dcache.scala 161:18]
        tags0_28 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_29 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1d == index) begin // @[dcache.scala 161:18]
        tags0_29 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_30 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1e == index) begin // @[dcache.scala 161:18]
        tags0_30 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_31 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h1f == index) begin // @[dcache.scala 161:18]
        tags0_31 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_32 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h20 == index) begin // @[dcache.scala 161:18]
        tags0_32 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_33 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h21 == index) begin // @[dcache.scala 161:18]
        tags0_33 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_34 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h22 == index) begin // @[dcache.scala 161:18]
        tags0_34 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_35 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h23 == index) begin // @[dcache.scala 161:18]
        tags0_35 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_36 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h24 == index) begin // @[dcache.scala 161:18]
        tags0_36 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_37 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h25 == index) begin // @[dcache.scala 161:18]
        tags0_37 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_38 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h26 == index) begin // @[dcache.scala 161:18]
        tags0_38 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_39 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h27 == index) begin // @[dcache.scala 161:18]
        tags0_39 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_40 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h28 == index) begin // @[dcache.scala 161:18]
        tags0_40 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_41 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h29 == index) begin // @[dcache.scala 161:18]
        tags0_41 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_42 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2a == index) begin // @[dcache.scala 161:18]
        tags0_42 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_43 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2b == index) begin // @[dcache.scala 161:18]
        tags0_43 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_44 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2c == index) begin // @[dcache.scala 161:18]
        tags0_44 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_45 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2d == index) begin // @[dcache.scala 161:18]
        tags0_45 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_46 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2e == index) begin // @[dcache.scala 161:18]
        tags0_46 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_47 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h2f == index) begin // @[dcache.scala 161:18]
        tags0_47 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_48 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h30 == index) begin // @[dcache.scala 161:18]
        tags0_48 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_49 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h31 == index) begin // @[dcache.scala 161:18]
        tags0_49 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_50 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h32 == index) begin // @[dcache.scala 161:18]
        tags0_50 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_51 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h33 == index) begin // @[dcache.scala 161:18]
        tags0_51 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_52 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h34 == index) begin // @[dcache.scala 161:18]
        tags0_52 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_53 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h35 == index) begin // @[dcache.scala 161:18]
        tags0_53 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_54 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h36 == index) begin // @[dcache.scala 161:18]
        tags0_54 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_55 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h37 == index) begin // @[dcache.scala 161:18]
        tags0_55 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_56 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h38 == index) begin // @[dcache.scala 161:18]
        tags0_56 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_57 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h39 == index) begin // @[dcache.scala 161:18]
        tags0_57 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_58 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3a == index) begin // @[dcache.scala 161:18]
        tags0_58 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_59 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3b == index) begin // @[dcache.scala 161:18]
        tags0_59 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_60 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3c == index) begin // @[dcache.scala 161:18]
        tags0_60 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_61 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3d == index) begin // @[dcache.scala 161:18]
        tags0_61 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_62 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3e == index) begin // @[dcache.scala 161:18]
        tags0_62 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_63 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h3f == index) begin // @[dcache.scala 161:18]
        tags0_63 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_64 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h40 == index) begin // @[dcache.scala 161:18]
        tags0_64 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_65 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h41 == index) begin // @[dcache.scala 161:18]
        tags0_65 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_66 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h42 == index) begin // @[dcache.scala 161:18]
        tags0_66 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_67 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h43 == index) begin // @[dcache.scala 161:18]
        tags0_67 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_68 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h44 == index) begin // @[dcache.scala 161:18]
        tags0_68 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_69 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h45 == index) begin // @[dcache.scala 161:18]
        tags0_69 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_70 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h46 == index) begin // @[dcache.scala 161:18]
        tags0_70 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_71 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h47 == index) begin // @[dcache.scala 161:18]
        tags0_71 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_72 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h48 == index) begin // @[dcache.scala 161:18]
        tags0_72 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_73 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h49 == index) begin // @[dcache.scala 161:18]
        tags0_73 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_74 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4a == index) begin // @[dcache.scala 161:18]
        tags0_74 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_75 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4b == index) begin // @[dcache.scala 161:18]
        tags0_75 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_76 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4c == index) begin // @[dcache.scala 161:18]
        tags0_76 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_77 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4d == index) begin // @[dcache.scala 161:18]
        tags0_77 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_78 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4e == index) begin // @[dcache.scala 161:18]
        tags0_78 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_79 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h4f == index) begin // @[dcache.scala 161:18]
        tags0_79 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_80 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h50 == index) begin // @[dcache.scala 161:18]
        tags0_80 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_81 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h51 == index) begin // @[dcache.scala 161:18]
        tags0_81 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_82 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h52 == index) begin // @[dcache.scala 161:18]
        tags0_82 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_83 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h53 == index) begin // @[dcache.scala 161:18]
        tags0_83 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_84 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h54 == index) begin // @[dcache.scala 161:18]
        tags0_84 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_85 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h55 == index) begin // @[dcache.scala 161:18]
        tags0_85 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_86 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h56 == index) begin // @[dcache.scala 161:18]
        tags0_86 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_87 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h57 == index) begin // @[dcache.scala 161:18]
        tags0_87 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_88 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h58 == index) begin // @[dcache.scala 161:18]
        tags0_88 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_89 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h59 == index) begin // @[dcache.scala 161:18]
        tags0_89 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_90 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5a == index) begin // @[dcache.scala 161:18]
        tags0_90 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_91 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5b == index) begin // @[dcache.scala 161:18]
        tags0_91 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_92 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5c == index) begin // @[dcache.scala 161:18]
        tags0_92 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_93 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5d == index) begin // @[dcache.scala 161:18]
        tags0_93 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_94 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5e == index) begin // @[dcache.scala 161:18]
        tags0_94 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_95 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h5f == index) begin // @[dcache.scala 161:18]
        tags0_95 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_96 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h60 == index) begin // @[dcache.scala 161:18]
        tags0_96 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_97 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h61 == index) begin // @[dcache.scala 161:18]
        tags0_97 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_98 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h62 == index) begin // @[dcache.scala 161:18]
        tags0_98 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_99 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h63 == index) begin // @[dcache.scala 161:18]
        tags0_99 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_100 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h64 == index) begin // @[dcache.scala 161:18]
        tags0_100 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_101 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h65 == index) begin // @[dcache.scala 161:18]
        tags0_101 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_102 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h66 == index) begin // @[dcache.scala 161:18]
        tags0_102 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_103 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h67 == index) begin // @[dcache.scala 161:18]
        tags0_103 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_104 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h68 == index) begin // @[dcache.scala 161:18]
        tags0_104 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_105 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h69 == index) begin // @[dcache.scala 161:18]
        tags0_105 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_106 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6a == index) begin // @[dcache.scala 161:18]
        tags0_106 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_107 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6b == index) begin // @[dcache.scala 161:18]
        tags0_107 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_108 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6c == index) begin // @[dcache.scala 161:18]
        tags0_108 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_109 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6d == index) begin // @[dcache.scala 161:18]
        tags0_109 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_110 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6e == index) begin // @[dcache.scala 161:18]
        tags0_110 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_111 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h6f == index) begin // @[dcache.scala 161:18]
        tags0_111 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_112 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h70 == index) begin // @[dcache.scala 161:18]
        tags0_112 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_113 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h71 == index) begin // @[dcache.scala 161:18]
        tags0_113 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_114 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h72 == index) begin // @[dcache.scala 161:18]
        tags0_114 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_115 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h73 == index) begin // @[dcache.scala 161:18]
        tags0_115 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_116 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h74 == index) begin // @[dcache.scala 161:18]
        tags0_116 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_117 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h75 == index) begin // @[dcache.scala 161:18]
        tags0_117 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_118 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h76 == index) begin // @[dcache.scala 161:18]
        tags0_118 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_119 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h77 == index) begin // @[dcache.scala 161:18]
        tags0_119 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_120 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h78 == index) begin // @[dcache.scala 161:18]
        tags0_120 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_121 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h79 == index) begin // @[dcache.scala 161:18]
        tags0_121 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_122 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7a == index) begin // @[dcache.scala 161:18]
        tags0_122 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_123 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7b == index) begin // @[dcache.scala 161:18]
        tags0_123 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_124 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7c == index) begin // @[dcache.scala 161:18]
        tags0_124 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_125 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7d == index) begin // @[dcache.scala 161:18]
        tags0_125 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_126 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7e == index) begin // @[dcache.scala 161:18]
        tags0_126 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 46:20]
      tags0_127 <= 53'h0; // @[dcache.scala 46:20]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      if (7'h7f == index) begin // @[dcache.scala 161:18]
        tags0_127 <= tag; // @[dcache.scala 161:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_0 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h0 == index) begin // @[dcache.scala 166:18]
        tags1_0 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_1 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1 == index) begin // @[dcache.scala 166:18]
        tags1_1 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_2 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2 == index) begin // @[dcache.scala 166:18]
        tags1_2 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_3 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3 == index) begin // @[dcache.scala 166:18]
        tags1_3 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_4 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4 == index) begin // @[dcache.scala 166:18]
        tags1_4 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_5 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5 == index) begin // @[dcache.scala 166:18]
        tags1_5 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_6 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6 == index) begin // @[dcache.scala 166:18]
        tags1_6 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_7 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7 == index) begin // @[dcache.scala 166:18]
        tags1_7 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_8 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h8 == index) begin // @[dcache.scala 166:18]
        tags1_8 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_9 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h9 == index) begin // @[dcache.scala 166:18]
        tags1_9 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_10 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'ha == index) begin // @[dcache.scala 166:18]
        tags1_10 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_11 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'hb == index) begin // @[dcache.scala 166:18]
        tags1_11 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_12 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'hc == index) begin // @[dcache.scala 166:18]
        tags1_12 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_13 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'hd == index) begin // @[dcache.scala 166:18]
        tags1_13 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_14 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'he == index) begin // @[dcache.scala 166:18]
        tags1_14 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_15 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'hf == index) begin // @[dcache.scala 166:18]
        tags1_15 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_16 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h10 == index) begin // @[dcache.scala 166:18]
        tags1_16 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_17 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h11 == index) begin // @[dcache.scala 166:18]
        tags1_17 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_18 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h12 == index) begin // @[dcache.scala 166:18]
        tags1_18 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_19 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h13 == index) begin // @[dcache.scala 166:18]
        tags1_19 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_20 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h14 == index) begin // @[dcache.scala 166:18]
        tags1_20 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_21 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h15 == index) begin // @[dcache.scala 166:18]
        tags1_21 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_22 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h16 == index) begin // @[dcache.scala 166:18]
        tags1_22 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_23 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h17 == index) begin // @[dcache.scala 166:18]
        tags1_23 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_24 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h18 == index) begin // @[dcache.scala 166:18]
        tags1_24 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_25 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h19 == index) begin // @[dcache.scala 166:18]
        tags1_25 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_26 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1a == index) begin // @[dcache.scala 166:18]
        tags1_26 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_27 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1b == index) begin // @[dcache.scala 166:18]
        tags1_27 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_28 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1c == index) begin // @[dcache.scala 166:18]
        tags1_28 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_29 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1d == index) begin // @[dcache.scala 166:18]
        tags1_29 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_30 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1e == index) begin // @[dcache.scala 166:18]
        tags1_30 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_31 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h1f == index) begin // @[dcache.scala 166:18]
        tags1_31 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_32 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h20 == index) begin // @[dcache.scala 166:18]
        tags1_32 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_33 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h21 == index) begin // @[dcache.scala 166:18]
        tags1_33 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_34 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h22 == index) begin // @[dcache.scala 166:18]
        tags1_34 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_35 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h23 == index) begin // @[dcache.scala 166:18]
        tags1_35 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_36 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h24 == index) begin // @[dcache.scala 166:18]
        tags1_36 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_37 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h25 == index) begin // @[dcache.scala 166:18]
        tags1_37 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_38 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h26 == index) begin // @[dcache.scala 166:18]
        tags1_38 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_39 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h27 == index) begin // @[dcache.scala 166:18]
        tags1_39 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_40 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h28 == index) begin // @[dcache.scala 166:18]
        tags1_40 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_41 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h29 == index) begin // @[dcache.scala 166:18]
        tags1_41 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_42 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2a == index) begin // @[dcache.scala 166:18]
        tags1_42 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_43 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2b == index) begin // @[dcache.scala 166:18]
        tags1_43 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_44 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2c == index) begin // @[dcache.scala 166:18]
        tags1_44 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_45 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2d == index) begin // @[dcache.scala 166:18]
        tags1_45 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_46 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2e == index) begin // @[dcache.scala 166:18]
        tags1_46 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_47 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h2f == index) begin // @[dcache.scala 166:18]
        tags1_47 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_48 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h30 == index) begin // @[dcache.scala 166:18]
        tags1_48 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_49 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h31 == index) begin // @[dcache.scala 166:18]
        tags1_49 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_50 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h32 == index) begin // @[dcache.scala 166:18]
        tags1_50 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_51 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h33 == index) begin // @[dcache.scala 166:18]
        tags1_51 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_52 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h34 == index) begin // @[dcache.scala 166:18]
        tags1_52 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_53 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h35 == index) begin // @[dcache.scala 166:18]
        tags1_53 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_54 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h36 == index) begin // @[dcache.scala 166:18]
        tags1_54 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_55 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h37 == index) begin // @[dcache.scala 166:18]
        tags1_55 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_56 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h38 == index) begin // @[dcache.scala 166:18]
        tags1_56 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_57 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h39 == index) begin // @[dcache.scala 166:18]
        tags1_57 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_58 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3a == index) begin // @[dcache.scala 166:18]
        tags1_58 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_59 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3b == index) begin // @[dcache.scala 166:18]
        tags1_59 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_60 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3c == index) begin // @[dcache.scala 166:18]
        tags1_60 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_61 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3d == index) begin // @[dcache.scala 166:18]
        tags1_61 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_62 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3e == index) begin // @[dcache.scala 166:18]
        tags1_62 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_63 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h3f == index) begin // @[dcache.scala 166:18]
        tags1_63 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_64 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h40 == index) begin // @[dcache.scala 166:18]
        tags1_64 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_65 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h41 == index) begin // @[dcache.scala 166:18]
        tags1_65 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_66 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h42 == index) begin // @[dcache.scala 166:18]
        tags1_66 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_67 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h43 == index) begin // @[dcache.scala 166:18]
        tags1_67 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_68 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h44 == index) begin // @[dcache.scala 166:18]
        tags1_68 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_69 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h45 == index) begin // @[dcache.scala 166:18]
        tags1_69 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_70 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h46 == index) begin // @[dcache.scala 166:18]
        tags1_70 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_71 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h47 == index) begin // @[dcache.scala 166:18]
        tags1_71 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_72 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h48 == index) begin // @[dcache.scala 166:18]
        tags1_72 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_73 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h49 == index) begin // @[dcache.scala 166:18]
        tags1_73 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_74 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4a == index) begin // @[dcache.scala 166:18]
        tags1_74 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_75 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4b == index) begin // @[dcache.scala 166:18]
        tags1_75 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_76 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4c == index) begin // @[dcache.scala 166:18]
        tags1_76 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_77 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4d == index) begin // @[dcache.scala 166:18]
        tags1_77 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_78 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4e == index) begin // @[dcache.scala 166:18]
        tags1_78 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_79 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h4f == index) begin // @[dcache.scala 166:18]
        tags1_79 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_80 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h50 == index) begin // @[dcache.scala 166:18]
        tags1_80 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_81 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h51 == index) begin // @[dcache.scala 166:18]
        tags1_81 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_82 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h52 == index) begin // @[dcache.scala 166:18]
        tags1_82 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_83 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h53 == index) begin // @[dcache.scala 166:18]
        tags1_83 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_84 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h54 == index) begin // @[dcache.scala 166:18]
        tags1_84 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_85 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h55 == index) begin // @[dcache.scala 166:18]
        tags1_85 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_86 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h56 == index) begin // @[dcache.scala 166:18]
        tags1_86 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_87 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h57 == index) begin // @[dcache.scala 166:18]
        tags1_87 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_88 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h58 == index) begin // @[dcache.scala 166:18]
        tags1_88 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_89 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h59 == index) begin // @[dcache.scala 166:18]
        tags1_89 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_90 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5a == index) begin // @[dcache.scala 166:18]
        tags1_90 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_91 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5b == index) begin // @[dcache.scala 166:18]
        tags1_91 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_92 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5c == index) begin // @[dcache.scala 166:18]
        tags1_92 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_93 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5d == index) begin // @[dcache.scala 166:18]
        tags1_93 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_94 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5e == index) begin // @[dcache.scala 166:18]
        tags1_94 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_95 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h5f == index) begin // @[dcache.scala 166:18]
        tags1_95 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_96 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h60 == index) begin // @[dcache.scala 166:18]
        tags1_96 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_97 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h61 == index) begin // @[dcache.scala 166:18]
        tags1_97 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_98 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h62 == index) begin // @[dcache.scala 166:18]
        tags1_98 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_99 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h63 == index) begin // @[dcache.scala 166:18]
        tags1_99 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_100 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h64 == index) begin // @[dcache.scala 166:18]
        tags1_100 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_101 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h65 == index) begin // @[dcache.scala 166:18]
        tags1_101 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_102 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h66 == index) begin // @[dcache.scala 166:18]
        tags1_102 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_103 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h67 == index) begin // @[dcache.scala 166:18]
        tags1_103 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_104 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h68 == index) begin // @[dcache.scala 166:18]
        tags1_104 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_105 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h69 == index) begin // @[dcache.scala 166:18]
        tags1_105 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_106 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6a == index) begin // @[dcache.scala 166:18]
        tags1_106 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_107 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6b == index) begin // @[dcache.scala 166:18]
        tags1_107 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_108 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6c == index) begin // @[dcache.scala 166:18]
        tags1_108 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_109 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6d == index) begin // @[dcache.scala 166:18]
        tags1_109 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_110 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6e == index) begin // @[dcache.scala 166:18]
        tags1_110 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_111 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h6f == index) begin // @[dcache.scala 166:18]
        tags1_111 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_112 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h70 == index) begin // @[dcache.scala 166:18]
        tags1_112 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_113 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h71 == index) begin // @[dcache.scala 166:18]
        tags1_113 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_114 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h72 == index) begin // @[dcache.scala 166:18]
        tags1_114 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_115 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h73 == index) begin // @[dcache.scala 166:18]
        tags1_115 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_116 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h74 == index) begin // @[dcache.scala 166:18]
        tags1_116 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_117 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h75 == index) begin // @[dcache.scala 166:18]
        tags1_117 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_118 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h76 == index) begin // @[dcache.scala 166:18]
        tags1_118 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_119 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h77 == index) begin // @[dcache.scala 166:18]
        tags1_119 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_120 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h78 == index) begin // @[dcache.scala 166:18]
        tags1_120 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_121 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h79 == index) begin // @[dcache.scala 166:18]
        tags1_121 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_122 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7a == index) begin // @[dcache.scala 166:18]
        tags1_122 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_123 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7b == index) begin // @[dcache.scala 166:18]
        tags1_123 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_124 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7c == index) begin // @[dcache.scala 166:18]
        tags1_124 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_125 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7d == index) begin // @[dcache.scala 166:18]
        tags1_125 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_126 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7e == index) begin // @[dcache.scala 166:18]
        tags1_126 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 47:20]
      tags1_127 <= 53'h0; // @[dcache.scala 47:20]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      if (7'h7f == index) begin // @[dcache.scala 166:18]
        tags1_127 <= tag; // @[dcache.scala 166:18]
      end
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_0 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_0 <= _GEN_775;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_1 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_1 <= _GEN_776;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_2 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_2 <= _GEN_777;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_3 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_3 <= _GEN_778;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_4 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_4 <= _GEN_779;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_5 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_5 <= _GEN_780;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_6 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_6 <= _GEN_781;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_7 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_7 <= _GEN_782;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_8 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_8 <= _GEN_783;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_9 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_9 <= _GEN_784;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_10 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_10 <= _GEN_785;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_11 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_11 <= _GEN_786;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_12 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_12 <= _GEN_787;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_13 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_13 <= _GEN_788;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_14 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_14 <= _GEN_789;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_15 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_15 <= _GEN_790;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_16 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_16 <= _GEN_791;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_17 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_17 <= _GEN_792;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_18 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_18 <= _GEN_793;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_19 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_19 <= _GEN_794;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_20 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_20 <= _GEN_795;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_21 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_21 <= _GEN_796;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_22 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_22 <= _GEN_797;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_23 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_23 <= _GEN_798;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_24 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_24 <= _GEN_799;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_25 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_25 <= _GEN_800;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_26 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_26 <= _GEN_801;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_27 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_27 <= _GEN_802;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_28 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_28 <= _GEN_803;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_29 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_29 <= _GEN_804;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_30 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_30 <= _GEN_805;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_31 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_31 <= _GEN_806;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_32 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_32 <= _GEN_807;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_33 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_33 <= _GEN_808;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_34 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_34 <= _GEN_809;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_35 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_35 <= _GEN_810;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_36 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_36 <= _GEN_811;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_37 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_37 <= _GEN_812;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_38 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_38 <= _GEN_813;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_39 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_39 <= _GEN_814;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_40 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_40 <= _GEN_815;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_41 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_41 <= _GEN_816;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_42 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_42 <= _GEN_817;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_43 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_43 <= _GEN_818;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_44 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_44 <= _GEN_819;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_45 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_45 <= _GEN_820;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_46 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_46 <= _GEN_821;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_47 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_47 <= _GEN_822;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_48 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_48 <= _GEN_823;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_49 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_49 <= _GEN_824;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_50 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_50 <= _GEN_825;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_51 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_51 <= _GEN_826;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_52 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_52 <= _GEN_827;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_53 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_53 <= _GEN_828;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_54 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_54 <= _GEN_829;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_55 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_55 <= _GEN_830;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_56 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_56 <= _GEN_831;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_57 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_57 <= _GEN_832;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_58 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_58 <= _GEN_833;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_59 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_59 <= _GEN_834;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_60 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_60 <= _GEN_835;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_61 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_61 <= _GEN_836;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_62 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_62 <= _GEN_837;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_63 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_63 <= _GEN_838;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_64 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_64 <= _GEN_839;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_65 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_65 <= _GEN_840;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_66 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_66 <= _GEN_841;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_67 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_67 <= _GEN_842;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_68 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_68 <= _GEN_843;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_69 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_69 <= _GEN_844;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_70 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_70 <= _GEN_845;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_71 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_71 <= _GEN_846;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_72 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_72 <= _GEN_847;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_73 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_73 <= _GEN_848;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_74 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_74 <= _GEN_849;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_75 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_75 <= _GEN_850;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_76 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_76 <= _GEN_851;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_77 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_77 <= _GEN_852;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_78 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_78 <= _GEN_853;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_79 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_79 <= _GEN_854;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_80 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_80 <= _GEN_855;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_81 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_81 <= _GEN_856;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_82 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_82 <= _GEN_857;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_83 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_83 <= _GEN_858;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_84 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_84 <= _GEN_859;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_85 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_85 <= _GEN_860;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_86 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_86 <= _GEN_861;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_87 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_87 <= _GEN_862;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_88 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_88 <= _GEN_863;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_89 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_89 <= _GEN_864;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_90 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_90 <= _GEN_865;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_91 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_91 <= _GEN_866;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_92 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_92 <= _GEN_867;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_93 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_93 <= _GEN_868;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_94 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_94 <= _GEN_869;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_95 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_95 <= _GEN_870;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_96 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_96 <= _GEN_871;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_97 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_97 <= _GEN_872;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_98 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_98 <= _GEN_873;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_99 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_99 <= _GEN_874;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_100 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_100 <= _GEN_875;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_101 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_101 <= _GEN_876;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_102 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_102 <= _GEN_877;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_103 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_103 <= _GEN_878;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_104 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_104 <= _GEN_879;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_105 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_105 <= _GEN_880;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_106 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_106 <= _GEN_881;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_107 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_107 <= _GEN_882;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_108 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_108 <= _GEN_883;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_109 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_109 <= _GEN_884;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_110 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_110 <= _GEN_885;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_111 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_111 <= _GEN_886;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_112 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_112 <= _GEN_887;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_113 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_113 <= _GEN_888;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_114 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_114 <= _GEN_889;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_115 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_115 <= _GEN_890;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_116 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_116 <= _GEN_891;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_117 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_117 <= _GEN_892;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_118 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_118 <= _GEN_893;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_119 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_119 <= _GEN_894;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_120 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_120 <= _GEN_895;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_121 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_121 <= _GEN_896;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_122 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_122 <= _GEN_897;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_123 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_123 <= _GEN_898;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_124 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_124 <= _GEN_899;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_125 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_125 <= _GEN_900;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_126 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_126 <= _GEN_901;
    end
    if (reset) begin // @[dcache.scala 48:21]
      valid0_127 <= 1'h0; // @[dcache.scala 48:21]
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      valid0_127 <= _GEN_902;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_0 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_0 <= _GEN_1543;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_1 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_1 <= _GEN_1544;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_2 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_2 <= _GEN_1545;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_3 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_3 <= _GEN_1546;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_4 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_4 <= _GEN_1547;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_5 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_5 <= _GEN_1548;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_6 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_6 <= _GEN_1549;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_7 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_7 <= _GEN_1550;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_8 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_8 <= _GEN_1551;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_9 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_9 <= _GEN_1552;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_10 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_10 <= _GEN_1553;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_11 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_11 <= _GEN_1554;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_12 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_12 <= _GEN_1555;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_13 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_13 <= _GEN_1556;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_14 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_14 <= _GEN_1557;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_15 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_15 <= _GEN_1558;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_16 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_16 <= _GEN_1559;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_17 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_17 <= _GEN_1560;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_18 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_18 <= _GEN_1561;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_19 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_19 <= _GEN_1562;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_20 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_20 <= _GEN_1563;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_21 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_21 <= _GEN_1564;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_22 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_22 <= _GEN_1565;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_23 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_23 <= _GEN_1566;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_24 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_24 <= _GEN_1567;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_25 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_25 <= _GEN_1568;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_26 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_26 <= _GEN_1569;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_27 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_27 <= _GEN_1570;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_28 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_28 <= _GEN_1571;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_29 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_29 <= _GEN_1572;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_30 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_30 <= _GEN_1573;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_31 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_31 <= _GEN_1574;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_32 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_32 <= _GEN_1575;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_33 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_33 <= _GEN_1576;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_34 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_34 <= _GEN_1577;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_35 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_35 <= _GEN_1578;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_36 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_36 <= _GEN_1579;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_37 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_37 <= _GEN_1580;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_38 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_38 <= _GEN_1581;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_39 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_39 <= _GEN_1582;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_40 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_40 <= _GEN_1583;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_41 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_41 <= _GEN_1584;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_42 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_42 <= _GEN_1585;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_43 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_43 <= _GEN_1586;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_44 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_44 <= _GEN_1587;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_45 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_45 <= _GEN_1588;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_46 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_46 <= _GEN_1589;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_47 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_47 <= _GEN_1590;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_48 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_48 <= _GEN_1591;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_49 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_49 <= _GEN_1592;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_50 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_50 <= _GEN_1593;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_51 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_51 <= _GEN_1594;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_52 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_52 <= _GEN_1595;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_53 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_53 <= _GEN_1596;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_54 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_54 <= _GEN_1597;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_55 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_55 <= _GEN_1598;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_56 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_56 <= _GEN_1599;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_57 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_57 <= _GEN_1600;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_58 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_58 <= _GEN_1601;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_59 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_59 <= _GEN_1602;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_60 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_60 <= _GEN_1603;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_61 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_61 <= _GEN_1604;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_62 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_62 <= _GEN_1605;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_63 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_63 <= _GEN_1606;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_64 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_64 <= _GEN_1607;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_65 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_65 <= _GEN_1608;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_66 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_66 <= _GEN_1609;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_67 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_67 <= _GEN_1610;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_68 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_68 <= _GEN_1611;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_69 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_69 <= _GEN_1612;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_70 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_70 <= _GEN_1613;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_71 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_71 <= _GEN_1614;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_72 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_72 <= _GEN_1615;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_73 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_73 <= _GEN_1616;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_74 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_74 <= _GEN_1617;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_75 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_75 <= _GEN_1618;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_76 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_76 <= _GEN_1619;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_77 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_77 <= _GEN_1620;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_78 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_78 <= _GEN_1621;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_79 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_79 <= _GEN_1622;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_80 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_80 <= _GEN_1623;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_81 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_81 <= _GEN_1624;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_82 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_82 <= _GEN_1625;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_83 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_83 <= _GEN_1626;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_84 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_84 <= _GEN_1627;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_85 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_85 <= _GEN_1628;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_86 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_86 <= _GEN_1629;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_87 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_87 <= _GEN_1630;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_88 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_88 <= _GEN_1631;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_89 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_89 <= _GEN_1632;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_90 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_90 <= _GEN_1633;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_91 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_91 <= _GEN_1634;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_92 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_92 <= _GEN_1635;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_93 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_93 <= _GEN_1636;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_94 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_94 <= _GEN_1637;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_95 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_95 <= _GEN_1638;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_96 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_96 <= _GEN_1639;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_97 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_97 <= _GEN_1640;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_98 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_98 <= _GEN_1641;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_99 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_99 <= _GEN_1642;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_100 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_100 <= _GEN_1643;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_101 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_101 <= _GEN_1644;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_102 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_102 <= _GEN_1645;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_103 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_103 <= _GEN_1646;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_104 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_104 <= _GEN_1647;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_105 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_105 <= _GEN_1648;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_106 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_106 <= _GEN_1649;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_107 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_107 <= _GEN_1650;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_108 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_108 <= _GEN_1651;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_109 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_109 <= _GEN_1652;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_110 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_110 <= _GEN_1653;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_111 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_111 <= _GEN_1654;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_112 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_112 <= _GEN_1655;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_113 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_113 <= _GEN_1656;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_114 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_114 <= _GEN_1657;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_115 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_115 <= _GEN_1658;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_116 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_116 <= _GEN_1659;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_117 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_117 <= _GEN_1660;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_118 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_118 <= _GEN_1661;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_119 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_119 <= _GEN_1662;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_120 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_120 <= _GEN_1663;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_121 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_121 <= _GEN_1664;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_122 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_122 <= _GEN_1665;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_123 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_123 <= _GEN_1666;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_124 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_124 <= _GEN_1667;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_125 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_125 <= _GEN_1668;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_126 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_126 <= _GEN_1669;
    end
    if (reset) begin // @[dcache.scala 49:21]
      valid1_127 <= 1'h0; // @[dcache.scala 49:21]
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      valid1_127 <= _GEN_1670;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_0 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_0 <= _GEN_2823;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_0 <= _GEN_2311;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_0 <= _GEN_903;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_1 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_1 <= _GEN_2824;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_1 <= _GEN_2312;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_1 <= _GEN_904;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_2 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_2 <= _GEN_2825;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_2 <= _GEN_2313;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_2 <= _GEN_905;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_3 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_3 <= _GEN_2826;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_3 <= _GEN_2314;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_3 <= _GEN_906;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_4 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_4 <= _GEN_2827;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_4 <= _GEN_2315;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_4 <= _GEN_907;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_5 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_5 <= _GEN_2828;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_5 <= _GEN_2316;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_5 <= _GEN_908;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_6 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_6 <= _GEN_2829;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_6 <= _GEN_2317;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_6 <= _GEN_909;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_7 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_7 <= _GEN_2830;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_7 <= _GEN_2318;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_7 <= _GEN_910;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_8 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_8 <= _GEN_2831;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_8 <= _GEN_2319;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_8 <= _GEN_911;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_9 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_9 <= _GEN_2832;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_9 <= _GEN_2320;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_9 <= _GEN_912;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_10 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_10 <= _GEN_2833;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_10 <= _GEN_2321;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_10 <= _GEN_913;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_11 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_11 <= _GEN_2834;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_11 <= _GEN_2322;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_11 <= _GEN_914;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_12 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_12 <= _GEN_2835;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_12 <= _GEN_2323;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_12 <= _GEN_915;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_13 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_13 <= _GEN_2836;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_13 <= _GEN_2324;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_13 <= _GEN_916;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_14 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_14 <= _GEN_2837;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_14 <= _GEN_2325;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_14 <= _GEN_917;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_15 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_15 <= _GEN_2838;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_15 <= _GEN_2326;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_15 <= _GEN_918;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_16 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_16 <= _GEN_2839;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_16 <= _GEN_2327;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_16 <= _GEN_919;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_17 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_17 <= _GEN_2840;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_17 <= _GEN_2328;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_17 <= _GEN_920;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_18 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_18 <= _GEN_2841;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_18 <= _GEN_2329;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_18 <= _GEN_921;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_19 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_19 <= _GEN_2842;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_19 <= _GEN_2330;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_19 <= _GEN_922;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_20 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_20 <= _GEN_2843;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_20 <= _GEN_2331;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_20 <= _GEN_923;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_21 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_21 <= _GEN_2844;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_21 <= _GEN_2332;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_21 <= _GEN_924;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_22 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_22 <= _GEN_2845;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_22 <= _GEN_2333;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_22 <= _GEN_925;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_23 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_23 <= _GEN_2846;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_23 <= _GEN_2334;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_23 <= _GEN_926;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_24 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_24 <= _GEN_2847;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_24 <= _GEN_2335;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_24 <= _GEN_927;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_25 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_25 <= _GEN_2848;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_25 <= _GEN_2336;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_25 <= _GEN_928;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_26 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_26 <= _GEN_2849;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_26 <= _GEN_2337;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_26 <= _GEN_929;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_27 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_27 <= _GEN_2850;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_27 <= _GEN_2338;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_27 <= _GEN_930;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_28 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_28 <= _GEN_2851;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_28 <= _GEN_2339;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_28 <= _GEN_931;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_29 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_29 <= _GEN_2852;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_29 <= _GEN_2340;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_29 <= _GEN_932;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_30 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_30 <= _GEN_2853;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_30 <= _GEN_2341;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_30 <= _GEN_933;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_31 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_31 <= _GEN_2854;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_31 <= _GEN_2342;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_31 <= _GEN_934;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_32 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_32 <= _GEN_2855;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_32 <= _GEN_2343;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_32 <= _GEN_935;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_33 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_33 <= _GEN_2856;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_33 <= _GEN_2344;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_33 <= _GEN_936;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_34 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_34 <= _GEN_2857;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_34 <= _GEN_2345;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_34 <= _GEN_937;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_35 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_35 <= _GEN_2858;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_35 <= _GEN_2346;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_35 <= _GEN_938;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_36 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_36 <= _GEN_2859;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_36 <= _GEN_2347;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_36 <= _GEN_939;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_37 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_37 <= _GEN_2860;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_37 <= _GEN_2348;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_37 <= _GEN_940;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_38 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_38 <= _GEN_2861;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_38 <= _GEN_2349;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_38 <= _GEN_941;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_39 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_39 <= _GEN_2862;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_39 <= _GEN_2350;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_39 <= _GEN_942;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_40 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_40 <= _GEN_2863;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_40 <= _GEN_2351;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_40 <= _GEN_943;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_41 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_41 <= _GEN_2864;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_41 <= _GEN_2352;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_41 <= _GEN_944;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_42 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_42 <= _GEN_2865;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_42 <= _GEN_2353;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_42 <= _GEN_945;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_43 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_43 <= _GEN_2866;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_43 <= _GEN_2354;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_43 <= _GEN_946;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_44 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_44 <= _GEN_2867;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_44 <= _GEN_2355;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_44 <= _GEN_947;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_45 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_45 <= _GEN_2868;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_45 <= _GEN_2356;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_45 <= _GEN_948;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_46 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_46 <= _GEN_2869;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_46 <= _GEN_2357;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_46 <= _GEN_949;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_47 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_47 <= _GEN_2870;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_47 <= _GEN_2358;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_47 <= _GEN_950;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_48 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_48 <= _GEN_2871;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_48 <= _GEN_2359;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_48 <= _GEN_951;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_49 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_49 <= _GEN_2872;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_49 <= _GEN_2360;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_49 <= _GEN_952;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_50 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_50 <= _GEN_2873;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_50 <= _GEN_2361;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_50 <= _GEN_953;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_51 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_51 <= _GEN_2874;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_51 <= _GEN_2362;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_51 <= _GEN_954;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_52 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_52 <= _GEN_2875;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_52 <= _GEN_2363;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_52 <= _GEN_955;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_53 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_53 <= _GEN_2876;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_53 <= _GEN_2364;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_53 <= _GEN_956;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_54 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_54 <= _GEN_2877;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_54 <= _GEN_2365;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_54 <= _GEN_957;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_55 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_55 <= _GEN_2878;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_55 <= _GEN_2366;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_55 <= _GEN_958;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_56 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_56 <= _GEN_2879;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_56 <= _GEN_2367;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_56 <= _GEN_959;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_57 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_57 <= _GEN_2880;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_57 <= _GEN_2368;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_57 <= _GEN_960;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_58 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_58 <= _GEN_2881;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_58 <= _GEN_2369;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_58 <= _GEN_961;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_59 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_59 <= _GEN_2882;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_59 <= _GEN_2370;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_59 <= _GEN_962;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_60 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_60 <= _GEN_2883;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_60 <= _GEN_2371;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_60 <= _GEN_963;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_61 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_61 <= _GEN_2884;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_61 <= _GEN_2372;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_61 <= _GEN_964;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_62 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_62 <= _GEN_2885;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_62 <= _GEN_2373;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_62 <= _GEN_965;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_63 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_63 <= _GEN_2886;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_63 <= _GEN_2374;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_63 <= _GEN_966;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_64 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_64 <= _GEN_2887;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_64 <= _GEN_2375;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_64 <= _GEN_967;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_65 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_65 <= _GEN_2888;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_65 <= _GEN_2376;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_65 <= _GEN_968;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_66 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_66 <= _GEN_2889;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_66 <= _GEN_2377;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_66 <= _GEN_969;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_67 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_67 <= _GEN_2890;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_67 <= _GEN_2378;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_67 <= _GEN_970;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_68 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_68 <= _GEN_2891;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_68 <= _GEN_2379;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_68 <= _GEN_971;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_69 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_69 <= _GEN_2892;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_69 <= _GEN_2380;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_69 <= _GEN_972;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_70 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_70 <= _GEN_2893;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_70 <= _GEN_2381;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_70 <= _GEN_973;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_71 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_71 <= _GEN_2894;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_71 <= _GEN_2382;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_71 <= _GEN_974;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_72 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_72 <= _GEN_2895;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_72 <= _GEN_2383;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_72 <= _GEN_975;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_73 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_73 <= _GEN_2896;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_73 <= _GEN_2384;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_73 <= _GEN_976;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_74 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_74 <= _GEN_2897;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_74 <= _GEN_2385;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_74 <= _GEN_977;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_75 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_75 <= _GEN_2898;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_75 <= _GEN_2386;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_75 <= _GEN_978;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_76 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_76 <= _GEN_2899;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_76 <= _GEN_2387;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_76 <= _GEN_979;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_77 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_77 <= _GEN_2900;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_77 <= _GEN_2388;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_77 <= _GEN_980;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_78 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_78 <= _GEN_2901;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_78 <= _GEN_2389;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_78 <= _GEN_981;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_79 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_79 <= _GEN_2902;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_79 <= _GEN_2390;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_79 <= _GEN_982;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_80 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_80 <= _GEN_2903;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_80 <= _GEN_2391;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_80 <= _GEN_983;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_81 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_81 <= _GEN_2904;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_81 <= _GEN_2392;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_81 <= _GEN_984;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_82 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_82 <= _GEN_2905;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_82 <= _GEN_2393;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_82 <= _GEN_985;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_83 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_83 <= _GEN_2906;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_83 <= _GEN_2394;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_83 <= _GEN_986;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_84 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_84 <= _GEN_2907;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_84 <= _GEN_2395;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_84 <= _GEN_987;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_85 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_85 <= _GEN_2908;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_85 <= _GEN_2396;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_85 <= _GEN_988;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_86 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_86 <= _GEN_2909;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_86 <= _GEN_2397;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_86 <= _GEN_989;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_87 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_87 <= _GEN_2910;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_87 <= _GEN_2398;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_87 <= _GEN_990;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_88 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_88 <= _GEN_2911;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_88 <= _GEN_2399;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_88 <= _GEN_991;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_89 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_89 <= _GEN_2912;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_89 <= _GEN_2400;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_89 <= _GEN_992;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_90 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_90 <= _GEN_2913;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_90 <= _GEN_2401;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_90 <= _GEN_993;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_91 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_91 <= _GEN_2914;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_91 <= _GEN_2402;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_91 <= _GEN_994;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_92 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_92 <= _GEN_2915;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_92 <= _GEN_2403;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_92 <= _GEN_995;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_93 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_93 <= _GEN_2916;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_93 <= _GEN_2404;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_93 <= _GEN_996;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_94 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_94 <= _GEN_2917;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_94 <= _GEN_2405;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_94 <= _GEN_997;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_95 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_95 <= _GEN_2918;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_95 <= _GEN_2406;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_95 <= _GEN_998;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_96 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_96 <= _GEN_2919;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_96 <= _GEN_2407;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_96 <= _GEN_999;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_97 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_97 <= _GEN_2920;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_97 <= _GEN_2408;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_97 <= _GEN_1000;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_98 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_98 <= _GEN_2921;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_98 <= _GEN_2409;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_98 <= _GEN_1001;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_99 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_99 <= _GEN_2922;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_99 <= _GEN_2410;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_99 <= _GEN_1002;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_100 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_100 <= _GEN_2923;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_100 <= _GEN_2411;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_100 <= _GEN_1003;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_101 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_101 <= _GEN_2924;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_101 <= _GEN_2412;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_101 <= _GEN_1004;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_102 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_102 <= _GEN_2925;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_102 <= _GEN_2413;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_102 <= _GEN_1005;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_103 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_103 <= _GEN_2926;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_103 <= _GEN_2414;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_103 <= _GEN_1006;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_104 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_104 <= _GEN_2927;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_104 <= _GEN_2415;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_104 <= _GEN_1007;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_105 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_105 <= _GEN_2928;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_105 <= _GEN_2416;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_105 <= _GEN_1008;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_106 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_106 <= _GEN_2929;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_106 <= _GEN_2417;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_106 <= _GEN_1009;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_107 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_107 <= _GEN_2930;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_107 <= _GEN_2418;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_107 <= _GEN_1010;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_108 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_108 <= _GEN_2931;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_108 <= _GEN_2419;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_108 <= _GEN_1011;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_109 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_109 <= _GEN_2932;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_109 <= _GEN_2420;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_109 <= _GEN_1012;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_110 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_110 <= _GEN_2933;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_110 <= _GEN_2421;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_110 <= _GEN_1013;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_111 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_111 <= _GEN_2934;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_111 <= _GEN_2422;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_111 <= _GEN_1014;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_112 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_112 <= _GEN_2935;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_112 <= _GEN_2423;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_112 <= _GEN_1015;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_113 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_113 <= _GEN_2936;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_113 <= _GEN_2424;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_113 <= _GEN_1016;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_114 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_114 <= _GEN_2937;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_114 <= _GEN_2425;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_114 <= _GEN_1017;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_115 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_115 <= _GEN_2938;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_115 <= _GEN_2426;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_115 <= _GEN_1018;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_116 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_116 <= _GEN_2939;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_116 <= _GEN_2427;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_116 <= _GEN_1019;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_117 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_117 <= _GEN_2940;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_117 <= _GEN_2428;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_117 <= _GEN_1020;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_118 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_118 <= _GEN_2941;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_118 <= _GEN_2429;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_118 <= _GEN_1021;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_119 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_119 <= _GEN_2942;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_119 <= _GEN_2430;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_119 <= _GEN_1022;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_120 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_120 <= _GEN_2943;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_120 <= _GEN_2431;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_120 <= _GEN_1023;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_121 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_121 <= _GEN_2944;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_121 <= _GEN_2432;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_121 <= _GEN_1024;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_122 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_122 <= _GEN_2945;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_122 <= _GEN_2433;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_122 <= _GEN_1025;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_123 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_123 <= _GEN_2946;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_123 <= _GEN_2434;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_123 <= _GEN_1026;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_124 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_124 <= _GEN_2947;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_124 <= _GEN_2435;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_124 <= _GEN_1027;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_125 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_125 <= _GEN_2948;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_125 <= _GEN_2436;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_125 <= _GEN_1028;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_126 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_126 <= _GEN_2949;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_126 <= _GEN_2437;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_126 <= _GEN_1029;
    end
    if (reset) begin // @[dcache.scala 50:21]
      dirty0_127 <= 1'h0; // @[dcache.scala 50:21]
    end else if (_write_back_is_finishing_T & next_write_state == 3'h1 & write_state != 3'h1 & hit_bank_0) begin // @[dcache.scala 174:91]
      dirty0_127 <= _GEN_2950;
    end else if (cpu_mem_Mwout & hit_bank_0) begin // @[dcache.scala 168:42]
      dirty0_127 <= _GEN_2438;
    end else if (_T & _should_write_back_T & _data_array_0_io_i_wen_T_9 & _write_back_is_finishing_T) begin // @[dcache.scala 158:91]
      dirty0_127 <= _GEN_1030;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_0 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_0 <= _GEN_3079;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_0 <= _GEN_2567;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_0 <= _GEN_1671;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_1 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_1 <= _GEN_3080;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_1 <= _GEN_2568;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_1 <= _GEN_1672;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_2 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_2 <= _GEN_3081;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_2 <= _GEN_2569;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_2 <= _GEN_1673;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_3 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_3 <= _GEN_3082;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_3 <= _GEN_2570;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_3 <= _GEN_1674;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_4 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_4 <= _GEN_3083;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_4 <= _GEN_2571;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_4 <= _GEN_1675;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_5 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_5 <= _GEN_3084;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_5 <= _GEN_2572;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_5 <= _GEN_1676;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_6 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_6 <= _GEN_3085;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_6 <= _GEN_2573;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_6 <= _GEN_1677;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_7 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_7 <= _GEN_3086;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_7 <= _GEN_2574;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_7 <= _GEN_1678;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_8 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_8 <= _GEN_3087;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_8 <= _GEN_2575;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_8 <= _GEN_1679;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_9 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_9 <= _GEN_3088;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_9 <= _GEN_2576;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_9 <= _GEN_1680;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_10 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_10 <= _GEN_3089;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_10 <= _GEN_2577;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_10 <= _GEN_1681;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_11 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_11 <= _GEN_3090;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_11 <= _GEN_2578;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_11 <= _GEN_1682;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_12 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_12 <= _GEN_3091;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_12 <= _GEN_2579;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_12 <= _GEN_1683;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_13 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_13 <= _GEN_3092;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_13 <= _GEN_2580;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_13 <= _GEN_1684;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_14 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_14 <= _GEN_3093;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_14 <= _GEN_2581;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_14 <= _GEN_1685;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_15 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_15 <= _GEN_3094;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_15 <= _GEN_2582;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_15 <= _GEN_1686;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_16 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_16 <= _GEN_3095;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_16 <= _GEN_2583;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_16 <= _GEN_1687;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_17 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_17 <= _GEN_3096;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_17 <= _GEN_2584;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_17 <= _GEN_1688;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_18 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_18 <= _GEN_3097;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_18 <= _GEN_2585;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_18 <= _GEN_1689;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_19 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_19 <= _GEN_3098;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_19 <= _GEN_2586;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_19 <= _GEN_1690;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_20 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_20 <= _GEN_3099;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_20 <= _GEN_2587;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_20 <= _GEN_1691;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_21 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_21 <= _GEN_3100;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_21 <= _GEN_2588;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_21 <= _GEN_1692;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_22 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_22 <= _GEN_3101;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_22 <= _GEN_2589;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_22 <= _GEN_1693;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_23 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_23 <= _GEN_3102;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_23 <= _GEN_2590;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_23 <= _GEN_1694;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_24 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_24 <= _GEN_3103;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_24 <= _GEN_2591;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_24 <= _GEN_1695;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_25 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_25 <= _GEN_3104;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_25 <= _GEN_2592;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_25 <= _GEN_1696;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_26 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_26 <= _GEN_3105;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_26 <= _GEN_2593;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_26 <= _GEN_1697;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_27 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_27 <= _GEN_3106;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_27 <= _GEN_2594;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_27 <= _GEN_1698;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_28 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_28 <= _GEN_3107;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_28 <= _GEN_2595;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_28 <= _GEN_1699;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_29 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_29 <= _GEN_3108;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_29 <= _GEN_2596;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_29 <= _GEN_1700;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_30 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_30 <= _GEN_3109;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_30 <= _GEN_2597;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_30 <= _GEN_1701;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_31 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_31 <= _GEN_3110;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_31 <= _GEN_2598;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_31 <= _GEN_1702;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_32 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_32 <= _GEN_3111;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_32 <= _GEN_2599;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_32 <= _GEN_1703;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_33 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_33 <= _GEN_3112;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_33 <= _GEN_2600;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_33 <= _GEN_1704;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_34 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_34 <= _GEN_3113;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_34 <= _GEN_2601;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_34 <= _GEN_1705;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_35 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_35 <= _GEN_3114;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_35 <= _GEN_2602;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_35 <= _GEN_1706;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_36 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_36 <= _GEN_3115;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_36 <= _GEN_2603;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_36 <= _GEN_1707;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_37 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_37 <= _GEN_3116;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_37 <= _GEN_2604;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_37 <= _GEN_1708;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_38 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_38 <= _GEN_3117;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_38 <= _GEN_2605;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_38 <= _GEN_1709;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_39 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_39 <= _GEN_3118;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_39 <= _GEN_2606;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_39 <= _GEN_1710;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_40 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_40 <= _GEN_3119;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_40 <= _GEN_2607;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_40 <= _GEN_1711;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_41 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_41 <= _GEN_3120;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_41 <= _GEN_2608;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_41 <= _GEN_1712;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_42 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_42 <= _GEN_3121;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_42 <= _GEN_2609;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_42 <= _GEN_1713;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_43 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_43 <= _GEN_3122;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_43 <= _GEN_2610;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_43 <= _GEN_1714;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_44 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_44 <= _GEN_3123;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_44 <= _GEN_2611;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_44 <= _GEN_1715;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_45 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_45 <= _GEN_3124;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_45 <= _GEN_2612;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_45 <= _GEN_1716;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_46 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_46 <= _GEN_3125;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_46 <= _GEN_2613;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_46 <= _GEN_1717;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_47 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_47 <= _GEN_3126;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_47 <= _GEN_2614;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_47 <= _GEN_1718;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_48 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_48 <= _GEN_3127;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_48 <= _GEN_2615;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_48 <= _GEN_1719;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_49 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_49 <= _GEN_3128;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_49 <= _GEN_2616;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_49 <= _GEN_1720;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_50 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_50 <= _GEN_3129;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_50 <= _GEN_2617;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_50 <= _GEN_1721;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_51 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_51 <= _GEN_3130;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_51 <= _GEN_2618;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_51 <= _GEN_1722;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_52 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_52 <= _GEN_3131;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_52 <= _GEN_2619;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_52 <= _GEN_1723;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_53 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_53 <= _GEN_3132;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_53 <= _GEN_2620;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_53 <= _GEN_1724;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_54 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_54 <= _GEN_3133;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_54 <= _GEN_2621;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_54 <= _GEN_1725;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_55 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_55 <= _GEN_3134;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_55 <= _GEN_2622;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_55 <= _GEN_1726;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_56 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_56 <= _GEN_3135;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_56 <= _GEN_2623;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_56 <= _GEN_1727;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_57 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_57 <= _GEN_3136;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_57 <= _GEN_2624;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_57 <= _GEN_1728;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_58 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_58 <= _GEN_3137;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_58 <= _GEN_2625;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_58 <= _GEN_1729;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_59 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_59 <= _GEN_3138;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_59 <= _GEN_2626;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_59 <= _GEN_1730;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_60 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_60 <= _GEN_3139;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_60 <= _GEN_2627;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_60 <= _GEN_1731;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_61 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_61 <= _GEN_3140;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_61 <= _GEN_2628;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_61 <= _GEN_1732;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_62 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_62 <= _GEN_3141;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_62 <= _GEN_2629;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_62 <= _GEN_1733;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_63 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_63 <= _GEN_3142;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_63 <= _GEN_2630;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_63 <= _GEN_1734;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_64 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_64 <= _GEN_3143;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_64 <= _GEN_2631;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_64 <= _GEN_1735;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_65 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_65 <= _GEN_3144;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_65 <= _GEN_2632;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_65 <= _GEN_1736;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_66 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_66 <= _GEN_3145;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_66 <= _GEN_2633;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_66 <= _GEN_1737;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_67 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_67 <= _GEN_3146;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_67 <= _GEN_2634;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_67 <= _GEN_1738;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_68 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_68 <= _GEN_3147;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_68 <= _GEN_2635;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_68 <= _GEN_1739;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_69 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_69 <= _GEN_3148;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_69 <= _GEN_2636;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_69 <= _GEN_1740;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_70 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_70 <= _GEN_3149;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_70 <= _GEN_2637;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_70 <= _GEN_1741;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_71 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_71 <= _GEN_3150;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_71 <= _GEN_2638;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_71 <= _GEN_1742;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_72 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_72 <= _GEN_3151;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_72 <= _GEN_2639;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_72 <= _GEN_1743;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_73 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_73 <= _GEN_3152;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_73 <= _GEN_2640;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_73 <= _GEN_1744;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_74 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_74 <= _GEN_3153;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_74 <= _GEN_2641;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_74 <= _GEN_1745;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_75 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_75 <= _GEN_3154;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_75 <= _GEN_2642;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_75 <= _GEN_1746;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_76 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_76 <= _GEN_3155;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_76 <= _GEN_2643;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_76 <= _GEN_1747;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_77 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_77 <= _GEN_3156;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_77 <= _GEN_2644;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_77 <= _GEN_1748;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_78 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_78 <= _GEN_3157;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_78 <= _GEN_2645;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_78 <= _GEN_1749;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_79 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_79 <= _GEN_3158;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_79 <= _GEN_2646;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_79 <= _GEN_1750;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_80 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_80 <= _GEN_3159;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_80 <= _GEN_2647;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_80 <= _GEN_1751;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_81 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_81 <= _GEN_3160;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_81 <= _GEN_2648;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_81 <= _GEN_1752;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_82 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_82 <= _GEN_3161;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_82 <= _GEN_2649;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_82 <= _GEN_1753;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_83 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_83 <= _GEN_3162;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_83 <= _GEN_2650;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_83 <= _GEN_1754;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_84 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_84 <= _GEN_3163;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_84 <= _GEN_2651;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_84 <= _GEN_1755;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_85 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_85 <= _GEN_3164;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_85 <= _GEN_2652;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_85 <= _GEN_1756;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_86 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_86 <= _GEN_3165;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_86 <= _GEN_2653;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_86 <= _GEN_1757;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_87 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_87 <= _GEN_3166;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_87 <= _GEN_2654;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_87 <= _GEN_1758;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_88 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_88 <= _GEN_3167;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_88 <= _GEN_2655;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_88 <= _GEN_1759;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_89 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_89 <= _GEN_3168;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_89 <= _GEN_2656;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_89 <= _GEN_1760;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_90 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_90 <= _GEN_3169;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_90 <= _GEN_2657;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_90 <= _GEN_1761;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_91 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_91 <= _GEN_3170;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_91 <= _GEN_2658;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_91 <= _GEN_1762;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_92 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_92 <= _GEN_3171;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_92 <= _GEN_2659;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_92 <= _GEN_1763;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_93 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_93 <= _GEN_3172;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_93 <= _GEN_2660;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_93 <= _GEN_1764;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_94 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_94 <= _GEN_3173;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_94 <= _GEN_2661;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_94 <= _GEN_1765;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_95 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_95 <= _GEN_3174;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_95 <= _GEN_2662;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_95 <= _GEN_1766;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_96 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_96 <= _GEN_3175;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_96 <= _GEN_2663;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_96 <= _GEN_1767;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_97 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_97 <= _GEN_3176;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_97 <= _GEN_2664;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_97 <= _GEN_1768;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_98 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_98 <= _GEN_3177;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_98 <= _GEN_2665;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_98 <= _GEN_1769;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_99 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_99 <= _GEN_3178;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_99 <= _GEN_2666;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_99 <= _GEN_1770;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_100 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_100 <= _GEN_3179;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_100 <= _GEN_2667;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_100 <= _GEN_1771;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_101 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_101 <= _GEN_3180;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_101 <= _GEN_2668;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_101 <= _GEN_1772;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_102 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_102 <= _GEN_3181;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_102 <= _GEN_2669;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_102 <= _GEN_1773;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_103 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_103 <= _GEN_3182;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_103 <= _GEN_2670;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_103 <= _GEN_1774;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_104 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_104 <= _GEN_3183;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_104 <= _GEN_2671;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_104 <= _GEN_1775;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_105 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_105 <= _GEN_3184;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_105 <= _GEN_2672;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_105 <= _GEN_1776;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_106 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_106 <= _GEN_3185;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_106 <= _GEN_2673;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_106 <= _GEN_1777;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_107 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_107 <= _GEN_3186;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_107 <= _GEN_2674;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_107 <= _GEN_1778;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_108 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_108 <= _GEN_3187;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_108 <= _GEN_2675;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_108 <= _GEN_1779;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_109 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_109 <= _GEN_3188;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_109 <= _GEN_2676;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_109 <= _GEN_1780;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_110 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_110 <= _GEN_3189;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_110 <= _GEN_2677;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_110 <= _GEN_1781;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_111 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_111 <= _GEN_3190;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_111 <= _GEN_2678;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_111 <= _GEN_1782;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_112 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_112 <= _GEN_3191;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_112 <= _GEN_2679;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_112 <= _GEN_1783;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_113 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_113 <= _GEN_3192;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_113 <= _GEN_2680;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_113 <= _GEN_1784;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_114 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_114 <= _GEN_3193;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_114 <= _GEN_2681;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_114 <= _GEN_1785;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_115 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_115 <= _GEN_3194;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_115 <= _GEN_2682;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_115 <= _GEN_1786;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_116 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_116 <= _GEN_3195;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_116 <= _GEN_2683;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_116 <= _GEN_1787;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_117 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_117 <= _GEN_3196;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_117 <= _GEN_2684;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_117 <= _GEN_1788;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_118 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_118 <= _GEN_3197;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_118 <= _GEN_2685;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_118 <= _GEN_1789;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_119 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_119 <= _GEN_3198;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_119 <= _GEN_2686;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_119 <= _GEN_1790;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_120 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_120 <= _GEN_3199;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_120 <= _GEN_2687;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_120 <= _GEN_1791;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_121 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_121 <= _GEN_3200;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_121 <= _GEN_2688;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_121 <= _GEN_1792;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_122 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_122 <= _GEN_3201;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_122 <= _GEN_2689;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_122 <= _GEN_1793;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_123 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_123 <= _GEN_3202;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_123 <= _GEN_2690;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_123 <= _GEN_1794;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_124 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_124 <= _GEN_3203;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_124 <= _GEN_2691;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_124 <= _GEN_1795;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_125 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_125 <= _GEN_3204;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_125 <= _GEN_2692;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_125 <= _GEN_1796;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_126 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_126 <= _GEN_3205;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_126 <= _GEN_2693;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_126 <= _GEN_1797;
    end
    if (reset) begin // @[dcache.scala 51:21]
      dirty1_127 <= 1'h0; // @[dcache.scala 51:21]
    end else if (_T_23 & hit_bank_1) begin // @[dcache.scala 177:91]
      dirty1_127 <= _GEN_3206;
    end else if (cpu_mem_Mwout & hit_bank_1) begin // @[dcache.scala 171:42]
      dirty1_127 <= _GEN_2694;
    end else if (_T_3 & victim & _write_back_is_finishing_T) begin // @[dcache.scala 163:91]
      dirty1_127 <= _GEN_1798;
    end
    if (_victim_T_1) begin // @[Mux.scala 101:16]
      victim <= 1'h0;
    end else begin
      victim <= _victim_T_5;
    end
    if (reset) begin // @[dcache.scala 61:32]
      read_from_mem_buf <= 128'h0; // @[dcache.scala 61:32]
    end else if (io_mem_master_readData_valid) begin // @[dcache.scala 85:25]
      read_from_mem_buf <= io_mem_master_readData_bits_data;
    end
    if (reset) begin // @[dcache.scala 68:26]
      write_state <= 3'h0; // @[dcache.scala 68:26]
    end else if (_next_write_state_T) begin // @[Mux.scala 101:16]
      write_state <= 3'h1;
    end else if (_next_write_state_T_2) begin // @[Mux.scala 101:16]
      write_state <= 3'h3;
    end else if (_next_write_state_T_4) begin // @[Mux.scala 101:16]
      write_state <= 3'h4;
    end else begin
      write_state <= _next_write_state_T_20;
    end
    if (reset) begin // @[dcache.scala 72:20]
      state <= 2'h0; // @[dcache.scala 72:20]
    end else if (_next_state_T) begin // @[Mux.scala 101:16]
      state <= 2'h1;
    end else if (_next_state_T_5) begin // @[Mux.scala 101:16]
      state <= 2'h2;
    end else if (_next_state_T_7) begin // @[Mux.scala 101:16]
      state <= 2'h1;
    end else begin
      state <= _next_state_T_16;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cpu_mem_Mwout = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  cpu_mem_Maddr = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  cpu_mem_Men = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cpu_mem_Mlen = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  cpu_mem_MdataOut = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  last_req_Mwout = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  last_req_Maddr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  last_req_Men = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  last_req_Mlen = _RAND_8[31:0];
  _RAND_9 = {2{`RANDOM}};
  last_req_MdataOut = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  tags0_0 = _RAND_10[52:0];
  _RAND_11 = {2{`RANDOM}};
  tags0_1 = _RAND_11[52:0];
  _RAND_12 = {2{`RANDOM}};
  tags0_2 = _RAND_12[52:0];
  _RAND_13 = {2{`RANDOM}};
  tags0_3 = _RAND_13[52:0];
  _RAND_14 = {2{`RANDOM}};
  tags0_4 = _RAND_14[52:0];
  _RAND_15 = {2{`RANDOM}};
  tags0_5 = _RAND_15[52:0];
  _RAND_16 = {2{`RANDOM}};
  tags0_6 = _RAND_16[52:0];
  _RAND_17 = {2{`RANDOM}};
  tags0_7 = _RAND_17[52:0];
  _RAND_18 = {2{`RANDOM}};
  tags0_8 = _RAND_18[52:0];
  _RAND_19 = {2{`RANDOM}};
  tags0_9 = _RAND_19[52:0];
  _RAND_20 = {2{`RANDOM}};
  tags0_10 = _RAND_20[52:0];
  _RAND_21 = {2{`RANDOM}};
  tags0_11 = _RAND_21[52:0];
  _RAND_22 = {2{`RANDOM}};
  tags0_12 = _RAND_22[52:0];
  _RAND_23 = {2{`RANDOM}};
  tags0_13 = _RAND_23[52:0];
  _RAND_24 = {2{`RANDOM}};
  tags0_14 = _RAND_24[52:0];
  _RAND_25 = {2{`RANDOM}};
  tags0_15 = _RAND_25[52:0];
  _RAND_26 = {2{`RANDOM}};
  tags0_16 = _RAND_26[52:0];
  _RAND_27 = {2{`RANDOM}};
  tags0_17 = _RAND_27[52:0];
  _RAND_28 = {2{`RANDOM}};
  tags0_18 = _RAND_28[52:0];
  _RAND_29 = {2{`RANDOM}};
  tags0_19 = _RAND_29[52:0];
  _RAND_30 = {2{`RANDOM}};
  tags0_20 = _RAND_30[52:0];
  _RAND_31 = {2{`RANDOM}};
  tags0_21 = _RAND_31[52:0];
  _RAND_32 = {2{`RANDOM}};
  tags0_22 = _RAND_32[52:0];
  _RAND_33 = {2{`RANDOM}};
  tags0_23 = _RAND_33[52:0];
  _RAND_34 = {2{`RANDOM}};
  tags0_24 = _RAND_34[52:0];
  _RAND_35 = {2{`RANDOM}};
  tags0_25 = _RAND_35[52:0];
  _RAND_36 = {2{`RANDOM}};
  tags0_26 = _RAND_36[52:0];
  _RAND_37 = {2{`RANDOM}};
  tags0_27 = _RAND_37[52:0];
  _RAND_38 = {2{`RANDOM}};
  tags0_28 = _RAND_38[52:0];
  _RAND_39 = {2{`RANDOM}};
  tags0_29 = _RAND_39[52:0];
  _RAND_40 = {2{`RANDOM}};
  tags0_30 = _RAND_40[52:0];
  _RAND_41 = {2{`RANDOM}};
  tags0_31 = _RAND_41[52:0];
  _RAND_42 = {2{`RANDOM}};
  tags0_32 = _RAND_42[52:0];
  _RAND_43 = {2{`RANDOM}};
  tags0_33 = _RAND_43[52:0];
  _RAND_44 = {2{`RANDOM}};
  tags0_34 = _RAND_44[52:0];
  _RAND_45 = {2{`RANDOM}};
  tags0_35 = _RAND_45[52:0];
  _RAND_46 = {2{`RANDOM}};
  tags0_36 = _RAND_46[52:0];
  _RAND_47 = {2{`RANDOM}};
  tags0_37 = _RAND_47[52:0];
  _RAND_48 = {2{`RANDOM}};
  tags0_38 = _RAND_48[52:0];
  _RAND_49 = {2{`RANDOM}};
  tags0_39 = _RAND_49[52:0];
  _RAND_50 = {2{`RANDOM}};
  tags0_40 = _RAND_50[52:0];
  _RAND_51 = {2{`RANDOM}};
  tags0_41 = _RAND_51[52:0];
  _RAND_52 = {2{`RANDOM}};
  tags0_42 = _RAND_52[52:0];
  _RAND_53 = {2{`RANDOM}};
  tags0_43 = _RAND_53[52:0];
  _RAND_54 = {2{`RANDOM}};
  tags0_44 = _RAND_54[52:0];
  _RAND_55 = {2{`RANDOM}};
  tags0_45 = _RAND_55[52:0];
  _RAND_56 = {2{`RANDOM}};
  tags0_46 = _RAND_56[52:0];
  _RAND_57 = {2{`RANDOM}};
  tags0_47 = _RAND_57[52:0];
  _RAND_58 = {2{`RANDOM}};
  tags0_48 = _RAND_58[52:0];
  _RAND_59 = {2{`RANDOM}};
  tags0_49 = _RAND_59[52:0];
  _RAND_60 = {2{`RANDOM}};
  tags0_50 = _RAND_60[52:0];
  _RAND_61 = {2{`RANDOM}};
  tags0_51 = _RAND_61[52:0];
  _RAND_62 = {2{`RANDOM}};
  tags0_52 = _RAND_62[52:0];
  _RAND_63 = {2{`RANDOM}};
  tags0_53 = _RAND_63[52:0];
  _RAND_64 = {2{`RANDOM}};
  tags0_54 = _RAND_64[52:0];
  _RAND_65 = {2{`RANDOM}};
  tags0_55 = _RAND_65[52:0];
  _RAND_66 = {2{`RANDOM}};
  tags0_56 = _RAND_66[52:0];
  _RAND_67 = {2{`RANDOM}};
  tags0_57 = _RAND_67[52:0];
  _RAND_68 = {2{`RANDOM}};
  tags0_58 = _RAND_68[52:0];
  _RAND_69 = {2{`RANDOM}};
  tags0_59 = _RAND_69[52:0];
  _RAND_70 = {2{`RANDOM}};
  tags0_60 = _RAND_70[52:0];
  _RAND_71 = {2{`RANDOM}};
  tags0_61 = _RAND_71[52:0];
  _RAND_72 = {2{`RANDOM}};
  tags0_62 = _RAND_72[52:0];
  _RAND_73 = {2{`RANDOM}};
  tags0_63 = _RAND_73[52:0];
  _RAND_74 = {2{`RANDOM}};
  tags0_64 = _RAND_74[52:0];
  _RAND_75 = {2{`RANDOM}};
  tags0_65 = _RAND_75[52:0];
  _RAND_76 = {2{`RANDOM}};
  tags0_66 = _RAND_76[52:0];
  _RAND_77 = {2{`RANDOM}};
  tags0_67 = _RAND_77[52:0];
  _RAND_78 = {2{`RANDOM}};
  tags0_68 = _RAND_78[52:0];
  _RAND_79 = {2{`RANDOM}};
  tags0_69 = _RAND_79[52:0];
  _RAND_80 = {2{`RANDOM}};
  tags0_70 = _RAND_80[52:0];
  _RAND_81 = {2{`RANDOM}};
  tags0_71 = _RAND_81[52:0];
  _RAND_82 = {2{`RANDOM}};
  tags0_72 = _RAND_82[52:0];
  _RAND_83 = {2{`RANDOM}};
  tags0_73 = _RAND_83[52:0];
  _RAND_84 = {2{`RANDOM}};
  tags0_74 = _RAND_84[52:0];
  _RAND_85 = {2{`RANDOM}};
  tags0_75 = _RAND_85[52:0];
  _RAND_86 = {2{`RANDOM}};
  tags0_76 = _RAND_86[52:0];
  _RAND_87 = {2{`RANDOM}};
  tags0_77 = _RAND_87[52:0];
  _RAND_88 = {2{`RANDOM}};
  tags0_78 = _RAND_88[52:0];
  _RAND_89 = {2{`RANDOM}};
  tags0_79 = _RAND_89[52:0];
  _RAND_90 = {2{`RANDOM}};
  tags0_80 = _RAND_90[52:0];
  _RAND_91 = {2{`RANDOM}};
  tags0_81 = _RAND_91[52:0];
  _RAND_92 = {2{`RANDOM}};
  tags0_82 = _RAND_92[52:0];
  _RAND_93 = {2{`RANDOM}};
  tags0_83 = _RAND_93[52:0];
  _RAND_94 = {2{`RANDOM}};
  tags0_84 = _RAND_94[52:0];
  _RAND_95 = {2{`RANDOM}};
  tags0_85 = _RAND_95[52:0];
  _RAND_96 = {2{`RANDOM}};
  tags0_86 = _RAND_96[52:0];
  _RAND_97 = {2{`RANDOM}};
  tags0_87 = _RAND_97[52:0];
  _RAND_98 = {2{`RANDOM}};
  tags0_88 = _RAND_98[52:0];
  _RAND_99 = {2{`RANDOM}};
  tags0_89 = _RAND_99[52:0];
  _RAND_100 = {2{`RANDOM}};
  tags0_90 = _RAND_100[52:0];
  _RAND_101 = {2{`RANDOM}};
  tags0_91 = _RAND_101[52:0];
  _RAND_102 = {2{`RANDOM}};
  tags0_92 = _RAND_102[52:0];
  _RAND_103 = {2{`RANDOM}};
  tags0_93 = _RAND_103[52:0];
  _RAND_104 = {2{`RANDOM}};
  tags0_94 = _RAND_104[52:0];
  _RAND_105 = {2{`RANDOM}};
  tags0_95 = _RAND_105[52:0];
  _RAND_106 = {2{`RANDOM}};
  tags0_96 = _RAND_106[52:0];
  _RAND_107 = {2{`RANDOM}};
  tags0_97 = _RAND_107[52:0];
  _RAND_108 = {2{`RANDOM}};
  tags0_98 = _RAND_108[52:0];
  _RAND_109 = {2{`RANDOM}};
  tags0_99 = _RAND_109[52:0];
  _RAND_110 = {2{`RANDOM}};
  tags0_100 = _RAND_110[52:0];
  _RAND_111 = {2{`RANDOM}};
  tags0_101 = _RAND_111[52:0];
  _RAND_112 = {2{`RANDOM}};
  tags0_102 = _RAND_112[52:0];
  _RAND_113 = {2{`RANDOM}};
  tags0_103 = _RAND_113[52:0];
  _RAND_114 = {2{`RANDOM}};
  tags0_104 = _RAND_114[52:0];
  _RAND_115 = {2{`RANDOM}};
  tags0_105 = _RAND_115[52:0];
  _RAND_116 = {2{`RANDOM}};
  tags0_106 = _RAND_116[52:0];
  _RAND_117 = {2{`RANDOM}};
  tags0_107 = _RAND_117[52:0];
  _RAND_118 = {2{`RANDOM}};
  tags0_108 = _RAND_118[52:0];
  _RAND_119 = {2{`RANDOM}};
  tags0_109 = _RAND_119[52:0];
  _RAND_120 = {2{`RANDOM}};
  tags0_110 = _RAND_120[52:0];
  _RAND_121 = {2{`RANDOM}};
  tags0_111 = _RAND_121[52:0];
  _RAND_122 = {2{`RANDOM}};
  tags0_112 = _RAND_122[52:0];
  _RAND_123 = {2{`RANDOM}};
  tags0_113 = _RAND_123[52:0];
  _RAND_124 = {2{`RANDOM}};
  tags0_114 = _RAND_124[52:0];
  _RAND_125 = {2{`RANDOM}};
  tags0_115 = _RAND_125[52:0];
  _RAND_126 = {2{`RANDOM}};
  tags0_116 = _RAND_126[52:0];
  _RAND_127 = {2{`RANDOM}};
  tags0_117 = _RAND_127[52:0];
  _RAND_128 = {2{`RANDOM}};
  tags0_118 = _RAND_128[52:0];
  _RAND_129 = {2{`RANDOM}};
  tags0_119 = _RAND_129[52:0];
  _RAND_130 = {2{`RANDOM}};
  tags0_120 = _RAND_130[52:0];
  _RAND_131 = {2{`RANDOM}};
  tags0_121 = _RAND_131[52:0];
  _RAND_132 = {2{`RANDOM}};
  tags0_122 = _RAND_132[52:0];
  _RAND_133 = {2{`RANDOM}};
  tags0_123 = _RAND_133[52:0];
  _RAND_134 = {2{`RANDOM}};
  tags0_124 = _RAND_134[52:0];
  _RAND_135 = {2{`RANDOM}};
  tags0_125 = _RAND_135[52:0];
  _RAND_136 = {2{`RANDOM}};
  tags0_126 = _RAND_136[52:0];
  _RAND_137 = {2{`RANDOM}};
  tags0_127 = _RAND_137[52:0];
  _RAND_138 = {2{`RANDOM}};
  tags1_0 = _RAND_138[52:0];
  _RAND_139 = {2{`RANDOM}};
  tags1_1 = _RAND_139[52:0];
  _RAND_140 = {2{`RANDOM}};
  tags1_2 = _RAND_140[52:0];
  _RAND_141 = {2{`RANDOM}};
  tags1_3 = _RAND_141[52:0];
  _RAND_142 = {2{`RANDOM}};
  tags1_4 = _RAND_142[52:0];
  _RAND_143 = {2{`RANDOM}};
  tags1_5 = _RAND_143[52:0];
  _RAND_144 = {2{`RANDOM}};
  tags1_6 = _RAND_144[52:0];
  _RAND_145 = {2{`RANDOM}};
  tags1_7 = _RAND_145[52:0];
  _RAND_146 = {2{`RANDOM}};
  tags1_8 = _RAND_146[52:0];
  _RAND_147 = {2{`RANDOM}};
  tags1_9 = _RAND_147[52:0];
  _RAND_148 = {2{`RANDOM}};
  tags1_10 = _RAND_148[52:0];
  _RAND_149 = {2{`RANDOM}};
  tags1_11 = _RAND_149[52:0];
  _RAND_150 = {2{`RANDOM}};
  tags1_12 = _RAND_150[52:0];
  _RAND_151 = {2{`RANDOM}};
  tags1_13 = _RAND_151[52:0];
  _RAND_152 = {2{`RANDOM}};
  tags1_14 = _RAND_152[52:0];
  _RAND_153 = {2{`RANDOM}};
  tags1_15 = _RAND_153[52:0];
  _RAND_154 = {2{`RANDOM}};
  tags1_16 = _RAND_154[52:0];
  _RAND_155 = {2{`RANDOM}};
  tags1_17 = _RAND_155[52:0];
  _RAND_156 = {2{`RANDOM}};
  tags1_18 = _RAND_156[52:0];
  _RAND_157 = {2{`RANDOM}};
  tags1_19 = _RAND_157[52:0];
  _RAND_158 = {2{`RANDOM}};
  tags1_20 = _RAND_158[52:0];
  _RAND_159 = {2{`RANDOM}};
  tags1_21 = _RAND_159[52:0];
  _RAND_160 = {2{`RANDOM}};
  tags1_22 = _RAND_160[52:0];
  _RAND_161 = {2{`RANDOM}};
  tags1_23 = _RAND_161[52:0];
  _RAND_162 = {2{`RANDOM}};
  tags1_24 = _RAND_162[52:0];
  _RAND_163 = {2{`RANDOM}};
  tags1_25 = _RAND_163[52:0];
  _RAND_164 = {2{`RANDOM}};
  tags1_26 = _RAND_164[52:0];
  _RAND_165 = {2{`RANDOM}};
  tags1_27 = _RAND_165[52:0];
  _RAND_166 = {2{`RANDOM}};
  tags1_28 = _RAND_166[52:0];
  _RAND_167 = {2{`RANDOM}};
  tags1_29 = _RAND_167[52:0];
  _RAND_168 = {2{`RANDOM}};
  tags1_30 = _RAND_168[52:0];
  _RAND_169 = {2{`RANDOM}};
  tags1_31 = _RAND_169[52:0];
  _RAND_170 = {2{`RANDOM}};
  tags1_32 = _RAND_170[52:0];
  _RAND_171 = {2{`RANDOM}};
  tags1_33 = _RAND_171[52:0];
  _RAND_172 = {2{`RANDOM}};
  tags1_34 = _RAND_172[52:0];
  _RAND_173 = {2{`RANDOM}};
  tags1_35 = _RAND_173[52:0];
  _RAND_174 = {2{`RANDOM}};
  tags1_36 = _RAND_174[52:0];
  _RAND_175 = {2{`RANDOM}};
  tags1_37 = _RAND_175[52:0];
  _RAND_176 = {2{`RANDOM}};
  tags1_38 = _RAND_176[52:0];
  _RAND_177 = {2{`RANDOM}};
  tags1_39 = _RAND_177[52:0];
  _RAND_178 = {2{`RANDOM}};
  tags1_40 = _RAND_178[52:0];
  _RAND_179 = {2{`RANDOM}};
  tags1_41 = _RAND_179[52:0];
  _RAND_180 = {2{`RANDOM}};
  tags1_42 = _RAND_180[52:0];
  _RAND_181 = {2{`RANDOM}};
  tags1_43 = _RAND_181[52:0];
  _RAND_182 = {2{`RANDOM}};
  tags1_44 = _RAND_182[52:0];
  _RAND_183 = {2{`RANDOM}};
  tags1_45 = _RAND_183[52:0];
  _RAND_184 = {2{`RANDOM}};
  tags1_46 = _RAND_184[52:0];
  _RAND_185 = {2{`RANDOM}};
  tags1_47 = _RAND_185[52:0];
  _RAND_186 = {2{`RANDOM}};
  tags1_48 = _RAND_186[52:0];
  _RAND_187 = {2{`RANDOM}};
  tags1_49 = _RAND_187[52:0];
  _RAND_188 = {2{`RANDOM}};
  tags1_50 = _RAND_188[52:0];
  _RAND_189 = {2{`RANDOM}};
  tags1_51 = _RAND_189[52:0];
  _RAND_190 = {2{`RANDOM}};
  tags1_52 = _RAND_190[52:0];
  _RAND_191 = {2{`RANDOM}};
  tags1_53 = _RAND_191[52:0];
  _RAND_192 = {2{`RANDOM}};
  tags1_54 = _RAND_192[52:0];
  _RAND_193 = {2{`RANDOM}};
  tags1_55 = _RAND_193[52:0];
  _RAND_194 = {2{`RANDOM}};
  tags1_56 = _RAND_194[52:0];
  _RAND_195 = {2{`RANDOM}};
  tags1_57 = _RAND_195[52:0];
  _RAND_196 = {2{`RANDOM}};
  tags1_58 = _RAND_196[52:0];
  _RAND_197 = {2{`RANDOM}};
  tags1_59 = _RAND_197[52:0];
  _RAND_198 = {2{`RANDOM}};
  tags1_60 = _RAND_198[52:0];
  _RAND_199 = {2{`RANDOM}};
  tags1_61 = _RAND_199[52:0];
  _RAND_200 = {2{`RANDOM}};
  tags1_62 = _RAND_200[52:0];
  _RAND_201 = {2{`RANDOM}};
  tags1_63 = _RAND_201[52:0];
  _RAND_202 = {2{`RANDOM}};
  tags1_64 = _RAND_202[52:0];
  _RAND_203 = {2{`RANDOM}};
  tags1_65 = _RAND_203[52:0];
  _RAND_204 = {2{`RANDOM}};
  tags1_66 = _RAND_204[52:0];
  _RAND_205 = {2{`RANDOM}};
  tags1_67 = _RAND_205[52:0];
  _RAND_206 = {2{`RANDOM}};
  tags1_68 = _RAND_206[52:0];
  _RAND_207 = {2{`RANDOM}};
  tags1_69 = _RAND_207[52:0];
  _RAND_208 = {2{`RANDOM}};
  tags1_70 = _RAND_208[52:0];
  _RAND_209 = {2{`RANDOM}};
  tags1_71 = _RAND_209[52:0];
  _RAND_210 = {2{`RANDOM}};
  tags1_72 = _RAND_210[52:0];
  _RAND_211 = {2{`RANDOM}};
  tags1_73 = _RAND_211[52:0];
  _RAND_212 = {2{`RANDOM}};
  tags1_74 = _RAND_212[52:0];
  _RAND_213 = {2{`RANDOM}};
  tags1_75 = _RAND_213[52:0];
  _RAND_214 = {2{`RANDOM}};
  tags1_76 = _RAND_214[52:0];
  _RAND_215 = {2{`RANDOM}};
  tags1_77 = _RAND_215[52:0];
  _RAND_216 = {2{`RANDOM}};
  tags1_78 = _RAND_216[52:0];
  _RAND_217 = {2{`RANDOM}};
  tags1_79 = _RAND_217[52:0];
  _RAND_218 = {2{`RANDOM}};
  tags1_80 = _RAND_218[52:0];
  _RAND_219 = {2{`RANDOM}};
  tags1_81 = _RAND_219[52:0];
  _RAND_220 = {2{`RANDOM}};
  tags1_82 = _RAND_220[52:0];
  _RAND_221 = {2{`RANDOM}};
  tags1_83 = _RAND_221[52:0];
  _RAND_222 = {2{`RANDOM}};
  tags1_84 = _RAND_222[52:0];
  _RAND_223 = {2{`RANDOM}};
  tags1_85 = _RAND_223[52:0];
  _RAND_224 = {2{`RANDOM}};
  tags1_86 = _RAND_224[52:0];
  _RAND_225 = {2{`RANDOM}};
  tags1_87 = _RAND_225[52:0];
  _RAND_226 = {2{`RANDOM}};
  tags1_88 = _RAND_226[52:0];
  _RAND_227 = {2{`RANDOM}};
  tags1_89 = _RAND_227[52:0];
  _RAND_228 = {2{`RANDOM}};
  tags1_90 = _RAND_228[52:0];
  _RAND_229 = {2{`RANDOM}};
  tags1_91 = _RAND_229[52:0];
  _RAND_230 = {2{`RANDOM}};
  tags1_92 = _RAND_230[52:0];
  _RAND_231 = {2{`RANDOM}};
  tags1_93 = _RAND_231[52:0];
  _RAND_232 = {2{`RANDOM}};
  tags1_94 = _RAND_232[52:0];
  _RAND_233 = {2{`RANDOM}};
  tags1_95 = _RAND_233[52:0];
  _RAND_234 = {2{`RANDOM}};
  tags1_96 = _RAND_234[52:0];
  _RAND_235 = {2{`RANDOM}};
  tags1_97 = _RAND_235[52:0];
  _RAND_236 = {2{`RANDOM}};
  tags1_98 = _RAND_236[52:0];
  _RAND_237 = {2{`RANDOM}};
  tags1_99 = _RAND_237[52:0];
  _RAND_238 = {2{`RANDOM}};
  tags1_100 = _RAND_238[52:0];
  _RAND_239 = {2{`RANDOM}};
  tags1_101 = _RAND_239[52:0];
  _RAND_240 = {2{`RANDOM}};
  tags1_102 = _RAND_240[52:0];
  _RAND_241 = {2{`RANDOM}};
  tags1_103 = _RAND_241[52:0];
  _RAND_242 = {2{`RANDOM}};
  tags1_104 = _RAND_242[52:0];
  _RAND_243 = {2{`RANDOM}};
  tags1_105 = _RAND_243[52:0];
  _RAND_244 = {2{`RANDOM}};
  tags1_106 = _RAND_244[52:0];
  _RAND_245 = {2{`RANDOM}};
  tags1_107 = _RAND_245[52:0];
  _RAND_246 = {2{`RANDOM}};
  tags1_108 = _RAND_246[52:0];
  _RAND_247 = {2{`RANDOM}};
  tags1_109 = _RAND_247[52:0];
  _RAND_248 = {2{`RANDOM}};
  tags1_110 = _RAND_248[52:0];
  _RAND_249 = {2{`RANDOM}};
  tags1_111 = _RAND_249[52:0];
  _RAND_250 = {2{`RANDOM}};
  tags1_112 = _RAND_250[52:0];
  _RAND_251 = {2{`RANDOM}};
  tags1_113 = _RAND_251[52:0];
  _RAND_252 = {2{`RANDOM}};
  tags1_114 = _RAND_252[52:0];
  _RAND_253 = {2{`RANDOM}};
  tags1_115 = _RAND_253[52:0];
  _RAND_254 = {2{`RANDOM}};
  tags1_116 = _RAND_254[52:0];
  _RAND_255 = {2{`RANDOM}};
  tags1_117 = _RAND_255[52:0];
  _RAND_256 = {2{`RANDOM}};
  tags1_118 = _RAND_256[52:0];
  _RAND_257 = {2{`RANDOM}};
  tags1_119 = _RAND_257[52:0];
  _RAND_258 = {2{`RANDOM}};
  tags1_120 = _RAND_258[52:0];
  _RAND_259 = {2{`RANDOM}};
  tags1_121 = _RAND_259[52:0];
  _RAND_260 = {2{`RANDOM}};
  tags1_122 = _RAND_260[52:0];
  _RAND_261 = {2{`RANDOM}};
  tags1_123 = _RAND_261[52:0];
  _RAND_262 = {2{`RANDOM}};
  tags1_124 = _RAND_262[52:0];
  _RAND_263 = {2{`RANDOM}};
  tags1_125 = _RAND_263[52:0];
  _RAND_264 = {2{`RANDOM}};
  tags1_126 = _RAND_264[52:0];
  _RAND_265 = {2{`RANDOM}};
  tags1_127 = _RAND_265[52:0];
  _RAND_266 = {1{`RANDOM}};
  valid0_0 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid0_1 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid0_2 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid0_3 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid0_4 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid0_5 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid0_6 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid0_7 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid0_8 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid0_9 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid0_10 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid0_11 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid0_12 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid0_13 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid0_14 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid0_15 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid0_16 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid0_17 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid0_18 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid0_19 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid0_20 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid0_21 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid0_22 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid0_23 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid0_24 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid0_25 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid0_26 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid0_27 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid0_28 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid0_29 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid0_30 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid0_31 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid0_32 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid0_33 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid0_34 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid0_35 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid0_36 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid0_37 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid0_38 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid0_39 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid0_40 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid0_41 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid0_42 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid0_43 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid0_44 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid0_45 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid0_46 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid0_47 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid0_48 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid0_49 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid0_50 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid0_51 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid0_52 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid0_53 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid0_54 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid0_55 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid0_56 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid0_57 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid0_58 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid0_59 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid0_60 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid0_61 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid0_62 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid0_63 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid0_64 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid0_65 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid0_66 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid0_67 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid0_68 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid0_69 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid0_70 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid0_71 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid0_72 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid0_73 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid0_74 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid0_75 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid0_76 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid0_77 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid0_78 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid0_79 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid0_80 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid0_81 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid0_82 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid0_83 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid0_84 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid0_85 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid0_86 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid0_87 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid0_88 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid0_89 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid0_90 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid0_91 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid0_92 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid0_93 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid0_94 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid0_95 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid0_96 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid0_97 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid0_98 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid0_99 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid0_100 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid0_101 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid0_102 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid0_103 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid0_104 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid0_105 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid0_106 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid0_107 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid0_108 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid0_109 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid0_110 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid0_111 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid0_112 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid0_113 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid0_114 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid0_115 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid0_116 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid0_117 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid0_118 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid0_119 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid0_120 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid0_121 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid0_122 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid0_123 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid0_124 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid0_125 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid0_126 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid0_127 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid1_0 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid1_1 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid1_2 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid1_3 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid1_4 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid1_5 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid1_6 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid1_7 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid1_8 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid1_9 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid1_10 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid1_11 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid1_12 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid1_13 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid1_14 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid1_15 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid1_16 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid1_17 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid1_18 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid1_19 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid1_20 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid1_21 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid1_22 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid1_23 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid1_24 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid1_25 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid1_26 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid1_27 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid1_28 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid1_29 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid1_30 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid1_31 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid1_32 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid1_33 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid1_34 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid1_35 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid1_36 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid1_37 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid1_38 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid1_39 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid1_40 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid1_41 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid1_42 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid1_43 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid1_44 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid1_45 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid1_46 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid1_47 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid1_48 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid1_49 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid1_50 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid1_51 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid1_52 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid1_53 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid1_54 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid1_55 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid1_56 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid1_57 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid1_58 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid1_59 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid1_60 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid1_61 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid1_62 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid1_63 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid1_64 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid1_65 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid1_66 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid1_67 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid1_68 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid1_69 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid1_70 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid1_71 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid1_72 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid1_73 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid1_74 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid1_75 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid1_76 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid1_77 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid1_78 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid1_79 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid1_80 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid1_81 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid1_82 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid1_83 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid1_84 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid1_85 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid1_86 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid1_87 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid1_88 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid1_89 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid1_90 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid1_91 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid1_92 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid1_93 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid1_94 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid1_95 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid1_96 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid1_97 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid1_98 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid1_99 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid1_100 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid1_101 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid1_102 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid1_103 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid1_104 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid1_105 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid1_106 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid1_107 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid1_108 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid1_109 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid1_110 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid1_111 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid1_112 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid1_113 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid1_114 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid1_115 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid1_116 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid1_117 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid1_118 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid1_119 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  valid1_120 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  valid1_121 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  valid1_122 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  valid1_123 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  valid1_124 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  valid1_125 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  valid1_126 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  valid1_127 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  dirty0_0 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  dirty0_1 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  dirty0_2 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  dirty0_3 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  dirty0_4 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  dirty0_5 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  dirty0_6 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  dirty0_7 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  dirty0_8 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  dirty0_9 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  dirty0_10 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  dirty0_11 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  dirty0_12 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  dirty0_13 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  dirty0_14 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  dirty0_15 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  dirty0_16 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  dirty0_17 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  dirty0_18 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  dirty0_19 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  dirty0_20 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  dirty0_21 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  dirty0_22 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  dirty0_23 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  dirty0_24 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  dirty0_25 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  dirty0_26 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  dirty0_27 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  dirty0_28 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  dirty0_29 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  dirty0_30 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  dirty0_31 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  dirty0_32 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  dirty0_33 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  dirty0_34 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  dirty0_35 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  dirty0_36 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  dirty0_37 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  dirty0_38 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  dirty0_39 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  dirty0_40 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  dirty0_41 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  dirty0_42 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  dirty0_43 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  dirty0_44 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  dirty0_45 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  dirty0_46 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  dirty0_47 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  dirty0_48 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  dirty0_49 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  dirty0_50 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  dirty0_51 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  dirty0_52 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  dirty0_53 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  dirty0_54 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  dirty0_55 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  dirty0_56 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  dirty0_57 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  dirty0_58 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  dirty0_59 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  dirty0_60 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  dirty0_61 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  dirty0_62 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  dirty0_63 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  dirty0_64 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  dirty0_65 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  dirty0_66 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  dirty0_67 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  dirty0_68 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  dirty0_69 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  dirty0_70 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  dirty0_71 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  dirty0_72 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  dirty0_73 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  dirty0_74 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  dirty0_75 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  dirty0_76 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  dirty0_77 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  dirty0_78 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  dirty0_79 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  dirty0_80 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  dirty0_81 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  dirty0_82 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  dirty0_83 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  dirty0_84 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  dirty0_85 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  dirty0_86 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  dirty0_87 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  dirty0_88 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  dirty0_89 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  dirty0_90 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  dirty0_91 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  dirty0_92 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  dirty0_93 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  dirty0_94 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  dirty0_95 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  dirty0_96 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  dirty0_97 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  dirty0_98 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  dirty0_99 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  dirty0_100 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  dirty0_101 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  dirty0_102 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  dirty0_103 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  dirty0_104 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  dirty0_105 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  dirty0_106 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  dirty0_107 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  dirty0_108 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  dirty0_109 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  dirty0_110 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  dirty0_111 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  dirty0_112 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  dirty0_113 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  dirty0_114 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  dirty0_115 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  dirty0_116 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  dirty0_117 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  dirty0_118 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  dirty0_119 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  dirty0_120 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  dirty0_121 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  dirty0_122 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  dirty0_123 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  dirty0_124 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  dirty0_125 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  dirty0_126 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  dirty0_127 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  dirty1_0 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  dirty1_1 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  dirty1_2 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  dirty1_3 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  dirty1_4 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  dirty1_5 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  dirty1_6 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  dirty1_7 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  dirty1_8 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  dirty1_9 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  dirty1_10 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  dirty1_11 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  dirty1_12 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  dirty1_13 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  dirty1_14 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  dirty1_15 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  dirty1_16 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  dirty1_17 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  dirty1_18 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  dirty1_19 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  dirty1_20 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  dirty1_21 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  dirty1_22 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  dirty1_23 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  dirty1_24 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  dirty1_25 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  dirty1_26 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  dirty1_27 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  dirty1_28 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  dirty1_29 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  dirty1_30 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  dirty1_31 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  dirty1_32 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  dirty1_33 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  dirty1_34 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  dirty1_35 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  dirty1_36 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  dirty1_37 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  dirty1_38 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  dirty1_39 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  dirty1_40 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  dirty1_41 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  dirty1_42 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  dirty1_43 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  dirty1_44 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  dirty1_45 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  dirty1_46 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  dirty1_47 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  dirty1_48 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  dirty1_49 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  dirty1_50 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  dirty1_51 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  dirty1_52 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  dirty1_53 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  dirty1_54 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  dirty1_55 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  dirty1_56 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  dirty1_57 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  dirty1_58 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  dirty1_59 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  dirty1_60 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  dirty1_61 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  dirty1_62 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  dirty1_63 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  dirty1_64 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  dirty1_65 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  dirty1_66 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  dirty1_67 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  dirty1_68 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  dirty1_69 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  dirty1_70 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  dirty1_71 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  dirty1_72 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  dirty1_73 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  dirty1_74 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  dirty1_75 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  dirty1_76 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  dirty1_77 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  dirty1_78 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  dirty1_79 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  dirty1_80 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  dirty1_81 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  dirty1_82 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  dirty1_83 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  dirty1_84 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  dirty1_85 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  dirty1_86 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  dirty1_87 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  dirty1_88 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  dirty1_89 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  dirty1_90 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  dirty1_91 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  dirty1_92 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  dirty1_93 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  dirty1_94 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  dirty1_95 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  dirty1_96 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  dirty1_97 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  dirty1_98 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  dirty1_99 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  dirty1_100 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  dirty1_101 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  dirty1_102 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  dirty1_103 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  dirty1_104 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  dirty1_105 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  dirty1_106 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  dirty1_107 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  dirty1_108 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  dirty1_109 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  dirty1_110 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  dirty1_111 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  dirty1_112 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  dirty1_113 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  dirty1_114 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  dirty1_115 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  dirty1_116 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  dirty1_117 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  dirty1_118 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  dirty1_119 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  dirty1_120 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  dirty1_121 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  dirty1_122 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  dirty1_123 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  dirty1_124 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  dirty1_125 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  dirty1_126 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  dirty1_127 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  victim = _RAND_778[0:0];
  _RAND_779 = {4{`RANDOM}};
  read_from_mem_buf = _RAND_779[127:0];
  _RAND_780 = {1{`RANDOM}};
  write_state = _RAND_780[2:0];
  _RAND_781 = {1{`RANDOM}};
  state = _RAND_781[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

module Icache(
  input          clock,
  input          reset,
  input          io_cpu_if_o_wen,
  input  [63:0]  io_cpu_if_o_addr,
  output [63:0]  io_cpu_if_i_data,
  output         io_cpu_if_i_addr_ready,
  input          io_cpu_if_o_addr_valid,
  output         io_cpu_if_i_data_valid,
  input          io_cpu_if_o_stall1,
  input          io_cpu_if_o_stall2,
  input          io_mem_master_readAddr_ready,
  output         io_mem_master_readAddr_valid,
  output [63:0]  io_mem_master_readAddr_bits_addr,
  output [2:0]   io_mem_master_readAddr_bits_prot,
  output         io_mem_master_readData_ready,
  input          io_mem_master_readData_valid,
  input  [127:0] io_mem_master_readData_bits_data,
  input  [1:0]   io_mem_master_readData_bits_resp,
  input          io_mem_master_writeAddr_ready,
  output         io_mem_master_writeAddr_valid,
  output [63:0]  io_mem_master_writeAddr_bits_addr,
  output [2:0]   io_mem_master_writeAddr_bits_prot,
  input          io_mem_master_writeData_ready,
  output         io_mem_master_writeData_valid,
  output [127:0] io_mem_master_writeData_bits_data,
  output [15:0]  io_mem_master_writeData_bits_strb,
  output         io_mem_master_writeResp_ready,
  input          io_mem_master_writeResp_valid,
  input  [1:0]   io_mem_master_writeResp_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [63:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [63:0] _RAND_152;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [63:0] _RAND_155;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [63:0] _RAND_188;
  reg [63:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [63:0] _RAND_192;
  reg [63:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [63:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [63:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [63:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [63:0] _RAND_203;
  reg [63:0] _RAND_204;
  reg [63:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [63:0] _RAND_207;
  reg [63:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [63:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [63:0] _RAND_215;
  reg [63:0] _RAND_216;
  reg [63:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [63:0] _RAND_219;
  reg [63:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [63:0] _RAND_223;
  reg [63:0] _RAND_224;
  reg [63:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [63:0] _RAND_227;
  reg [63:0] _RAND_228;
  reg [63:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [63:0] _RAND_232;
  reg [63:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [63:0] _RAND_236;
  reg [63:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [63:0] _RAND_239;
  reg [63:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [63:0] _RAND_243;
  reg [63:0] _RAND_244;
  reg [63:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [63:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [63:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [63:0] _RAND_252;
  reg [63:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [63:0] _RAND_255;
  reg [63:0] _RAND_256;
  reg [63:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [127:0] _RAND_516;
`endif // RANDOMIZE_REG_INIT
  wire  data_array_0_clock; // @[icache.scala 32:36]
  wire  data_array_0_reset; // @[icache.scala 32:36]
  wire  data_array_0_io_i_wen; // @[icache.scala 32:36]
  wire [15:0] data_array_0_io_i_wstrb; // @[icache.scala 32:36]
  wire [6:0] data_array_0_io_i_addr; // @[icache.scala 32:36]
  wire [127:0] data_array_0_io_i_wdata; // @[icache.scala 32:36]
  wire [127:0] data_array_0_io_o_rdata; // @[icache.scala 32:36]
  wire  data_array_1_clock; // @[icache.scala 32:36]
  wire  data_array_1_reset; // @[icache.scala 32:36]
  wire  data_array_1_io_i_wen; // @[icache.scala 32:36]
  wire [15:0] data_array_1_io_i_wstrb; // @[icache.scala 32:36]
  wire [6:0] data_array_1_io_i_addr; // @[icache.scala 32:36]
  wire [127:0] data_array_1_io_i_wdata; // @[icache.scala 32:36]
  wire [127:0] data_array_1_io_o_rdata; // @[icache.scala 32:36]
  reg [63:0] cpu_if1_o_addr; // @[icache.scala 24:22]
  reg [63:0] cpu_if2_o_addr; // @[icache.scala 25:22]
  reg [52:0] tags0_0; // @[icache.scala 28:20]
  reg [52:0] tags0_1; // @[icache.scala 28:20]
  reg [52:0] tags0_2; // @[icache.scala 28:20]
  reg [52:0] tags0_3; // @[icache.scala 28:20]
  reg [52:0] tags0_4; // @[icache.scala 28:20]
  reg [52:0] tags0_5; // @[icache.scala 28:20]
  reg [52:0] tags0_6; // @[icache.scala 28:20]
  reg [52:0] tags0_7; // @[icache.scala 28:20]
  reg [52:0] tags0_8; // @[icache.scala 28:20]
  reg [52:0] tags0_9; // @[icache.scala 28:20]
  reg [52:0] tags0_10; // @[icache.scala 28:20]
  reg [52:0] tags0_11; // @[icache.scala 28:20]
  reg [52:0] tags0_12; // @[icache.scala 28:20]
  reg [52:0] tags0_13; // @[icache.scala 28:20]
  reg [52:0] tags0_14; // @[icache.scala 28:20]
  reg [52:0] tags0_15; // @[icache.scala 28:20]
  reg [52:0] tags0_16; // @[icache.scala 28:20]
  reg [52:0] tags0_17; // @[icache.scala 28:20]
  reg [52:0] tags0_18; // @[icache.scala 28:20]
  reg [52:0] tags0_19; // @[icache.scala 28:20]
  reg [52:0] tags0_20; // @[icache.scala 28:20]
  reg [52:0] tags0_21; // @[icache.scala 28:20]
  reg [52:0] tags0_22; // @[icache.scala 28:20]
  reg [52:0] tags0_23; // @[icache.scala 28:20]
  reg [52:0] tags0_24; // @[icache.scala 28:20]
  reg [52:0] tags0_25; // @[icache.scala 28:20]
  reg [52:0] tags0_26; // @[icache.scala 28:20]
  reg [52:0] tags0_27; // @[icache.scala 28:20]
  reg [52:0] tags0_28; // @[icache.scala 28:20]
  reg [52:0] tags0_29; // @[icache.scala 28:20]
  reg [52:0] tags0_30; // @[icache.scala 28:20]
  reg [52:0] tags0_31; // @[icache.scala 28:20]
  reg [52:0] tags0_32; // @[icache.scala 28:20]
  reg [52:0] tags0_33; // @[icache.scala 28:20]
  reg [52:0] tags0_34; // @[icache.scala 28:20]
  reg [52:0] tags0_35; // @[icache.scala 28:20]
  reg [52:0] tags0_36; // @[icache.scala 28:20]
  reg [52:0] tags0_37; // @[icache.scala 28:20]
  reg [52:0] tags0_38; // @[icache.scala 28:20]
  reg [52:0] tags0_39; // @[icache.scala 28:20]
  reg [52:0] tags0_40; // @[icache.scala 28:20]
  reg [52:0] tags0_41; // @[icache.scala 28:20]
  reg [52:0] tags0_42; // @[icache.scala 28:20]
  reg [52:0] tags0_43; // @[icache.scala 28:20]
  reg [52:0] tags0_44; // @[icache.scala 28:20]
  reg [52:0] tags0_45; // @[icache.scala 28:20]
  reg [52:0] tags0_46; // @[icache.scala 28:20]
  reg [52:0] tags0_47; // @[icache.scala 28:20]
  reg [52:0] tags0_48; // @[icache.scala 28:20]
  reg [52:0] tags0_49; // @[icache.scala 28:20]
  reg [52:0] tags0_50; // @[icache.scala 28:20]
  reg [52:0] tags0_51; // @[icache.scala 28:20]
  reg [52:0] tags0_52; // @[icache.scala 28:20]
  reg [52:0] tags0_53; // @[icache.scala 28:20]
  reg [52:0] tags0_54; // @[icache.scala 28:20]
  reg [52:0] tags0_55; // @[icache.scala 28:20]
  reg [52:0] tags0_56; // @[icache.scala 28:20]
  reg [52:0] tags0_57; // @[icache.scala 28:20]
  reg [52:0] tags0_58; // @[icache.scala 28:20]
  reg [52:0] tags0_59; // @[icache.scala 28:20]
  reg [52:0] tags0_60; // @[icache.scala 28:20]
  reg [52:0] tags0_61; // @[icache.scala 28:20]
  reg [52:0] tags0_62; // @[icache.scala 28:20]
  reg [52:0] tags0_63; // @[icache.scala 28:20]
  reg [52:0] tags0_64; // @[icache.scala 28:20]
  reg [52:0] tags0_65; // @[icache.scala 28:20]
  reg [52:0] tags0_66; // @[icache.scala 28:20]
  reg [52:0] tags0_67; // @[icache.scala 28:20]
  reg [52:0] tags0_68; // @[icache.scala 28:20]
  reg [52:0] tags0_69; // @[icache.scala 28:20]
  reg [52:0] tags0_70; // @[icache.scala 28:20]
  reg [52:0] tags0_71; // @[icache.scala 28:20]
  reg [52:0] tags0_72; // @[icache.scala 28:20]
  reg [52:0] tags0_73; // @[icache.scala 28:20]
  reg [52:0] tags0_74; // @[icache.scala 28:20]
  reg [52:0] tags0_75; // @[icache.scala 28:20]
  reg [52:0] tags0_76; // @[icache.scala 28:20]
  reg [52:0] tags0_77; // @[icache.scala 28:20]
  reg [52:0] tags0_78; // @[icache.scala 28:20]
  reg [52:0] tags0_79; // @[icache.scala 28:20]
  reg [52:0] tags0_80; // @[icache.scala 28:20]
  reg [52:0] tags0_81; // @[icache.scala 28:20]
  reg [52:0] tags0_82; // @[icache.scala 28:20]
  reg [52:0] tags0_83; // @[icache.scala 28:20]
  reg [52:0] tags0_84; // @[icache.scala 28:20]
  reg [52:0] tags0_85; // @[icache.scala 28:20]
  reg [52:0] tags0_86; // @[icache.scala 28:20]
  reg [52:0] tags0_87; // @[icache.scala 28:20]
  reg [52:0] tags0_88; // @[icache.scala 28:20]
  reg [52:0] tags0_89; // @[icache.scala 28:20]
  reg [52:0] tags0_90; // @[icache.scala 28:20]
  reg [52:0] tags0_91; // @[icache.scala 28:20]
  reg [52:0] tags0_92; // @[icache.scala 28:20]
  reg [52:0] tags0_93; // @[icache.scala 28:20]
  reg [52:0] tags0_94; // @[icache.scala 28:20]
  reg [52:0] tags0_95; // @[icache.scala 28:20]
  reg [52:0] tags0_96; // @[icache.scala 28:20]
  reg [52:0] tags0_97; // @[icache.scala 28:20]
  reg [52:0] tags0_98; // @[icache.scala 28:20]
  reg [52:0] tags0_99; // @[icache.scala 28:20]
  reg [52:0] tags0_100; // @[icache.scala 28:20]
  reg [52:0] tags0_101; // @[icache.scala 28:20]
  reg [52:0] tags0_102; // @[icache.scala 28:20]
  reg [52:0] tags0_103; // @[icache.scala 28:20]
  reg [52:0] tags0_104; // @[icache.scala 28:20]
  reg [52:0] tags0_105; // @[icache.scala 28:20]
  reg [52:0] tags0_106; // @[icache.scala 28:20]
  reg [52:0] tags0_107; // @[icache.scala 28:20]
  reg [52:0] tags0_108; // @[icache.scala 28:20]
  reg [52:0] tags0_109; // @[icache.scala 28:20]
  reg [52:0] tags0_110; // @[icache.scala 28:20]
  reg [52:0] tags0_111; // @[icache.scala 28:20]
  reg [52:0] tags0_112; // @[icache.scala 28:20]
  reg [52:0] tags0_113; // @[icache.scala 28:20]
  reg [52:0] tags0_114; // @[icache.scala 28:20]
  reg [52:0] tags0_115; // @[icache.scala 28:20]
  reg [52:0] tags0_116; // @[icache.scala 28:20]
  reg [52:0] tags0_117; // @[icache.scala 28:20]
  reg [52:0] tags0_118; // @[icache.scala 28:20]
  reg [52:0] tags0_119; // @[icache.scala 28:20]
  reg [52:0] tags0_120; // @[icache.scala 28:20]
  reg [52:0] tags0_121; // @[icache.scala 28:20]
  reg [52:0] tags0_122; // @[icache.scala 28:20]
  reg [52:0] tags0_123; // @[icache.scala 28:20]
  reg [52:0] tags0_124; // @[icache.scala 28:20]
  reg [52:0] tags0_125; // @[icache.scala 28:20]
  reg [52:0] tags0_126; // @[icache.scala 28:20]
  reg [52:0] tags0_127; // @[icache.scala 28:20]
  reg [52:0] tags1_0; // @[icache.scala 29:20]
  reg [52:0] tags1_1; // @[icache.scala 29:20]
  reg [52:0] tags1_2; // @[icache.scala 29:20]
  reg [52:0] tags1_3; // @[icache.scala 29:20]
  reg [52:0] tags1_4; // @[icache.scala 29:20]
  reg [52:0] tags1_5; // @[icache.scala 29:20]
  reg [52:0] tags1_6; // @[icache.scala 29:20]
  reg [52:0] tags1_7; // @[icache.scala 29:20]
  reg [52:0] tags1_8; // @[icache.scala 29:20]
  reg [52:0] tags1_9; // @[icache.scala 29:20]
  reg [52:0] tags1_10; // @[icache.scala 29:20]
  reg [52:0] tags1_11; // @[icache.scala 29:20]
  reg [52:0] tags1_12; // @[icache.scala 29:20]
  reg [52:0] tags1_13; // @[icache.scala 29:20]
  reg [52:0] tags1_14; // @[icache.scala 29:20]
  reg [52:0] tags1_15; // @[icache.scala 29:20]
  reg [52:0] tags1_16; // @[icache.scala 29:20]
  reg [52:0] tags1_17; // @[icache.scala 29:20]
  reg [52:0] tags1_18; // @[icache.scala 29:20]
  reg [52:0] tags1_19; // @[icache.scala 29:20]
  reg [52:0] tags1_20; // @[icache.scala 29:20]
  reg [52:0] tags1_21; // @[icache.scala 29:20]
  reg [52:0] tags1_22; // @[icache.scala 29:20]
  reg [52:0] tags1_23; // @[icache.scala 29:20]
  reg [52:0] tags1_24; // @[icache.scala 29:20]
  reg [52:0] tags1_25; // @[icache.scala 29:20]
  reg [52:0] tags1_26; // @[icache.scala 29:20]
  reg [52:0] tags1_27; // @[icache.scala 29:20]
  reg [52:0] tags1_28; // @[icache.scala 29:20]
  reg [52:0] tags1_29; // @[icache.scala 29:20]
  reg [52:0] tags1_30; // @[icache.scala 29:20]
  reg [52:0] tags1_31; // @[icache.scala 29:20]
  reg [52:0] tags1_32; // @[icache.scala 29:20]
  reg [52:0] tags1_33; // @[icache.scala 29:20]
  reg [52:0] tags1_34; // @[icache.scala 29:20]
  reg [52:0] tags1_35; // @[icache.scala 29:20]
  reg [52:0] tags1_36; // @[icache.scala 29:20]
  reg [52:0] tags1_37; // @[icache.scala 29:20]
  reg [52:0] tags1_38; // @[icache.scala 29:20]
  reg [52:0] tags1_39; // @[icache.scala 29:20]
  reg [52:0] tags1_40; // @[icache.scala 29:20]
  reg [52:0] tags1_41; // @[icache.scala 29:20]
  reg [52:0] tags1_42; // @[icache.scala 29:20]
  reg [52:0] tags1_43; // @[icache.scala 29:20]
  reg [52:0] tags1_44; // @[icache.scala 29:20]
  reg [52:0] tags1_45; // @[icache.scala 29:20]
  reg [52:0] tags1_46; // @[icache.scala 29:20]
  reg [52:0] tags1_47; // @[icache.scala 29:20]
  reg [52:0] tags1_48; // @[icache.scala 29:20]
  reg [52:0] tags1_49; // @[icache.scala 29:20]
  reg [52:0] tags1_50; // @[icache.scala 29:20]
  reg [52:0] tags1_51; // @[icache.scala 29:20]
  reg [52:0] tags1_52; // @[icache.scala 29:20]
  reg [52:0] tags1_53; // @[icache.scala 29:20]
  reg [52:0] tags1_54; // @[icache.scala 29:20]
  reg [52:0] tags1_55; // @[icache.scala 29:20]
  reg [52:0] tags1_56; // @[icache.scala 29:20]
  reg [52:0] tags1_57; // @[icache.scala 29:20]
  reg [52:0] tags1_58; // @[icache.scala 29:20]
  reg [52:0] tags1_59; // @[icache.scala 29:20]
  reg [52:0] tags1_60; // @[icache.scala 29:20]
  reg [52:0] tags1_61; // @[icache.scala 29:20]
  reg [52:0] tags1_62; // @[icache.scala 29:20]
  reg [52:0] tags1_63; // @[icache.scala 29:20]
  reg [52:0] tags1_64; // @[icache.scala 29:20]
  reg [52:0] tags1_65; // @[icache.scala 29:20]
  reg [52:0] tags1_66; // @[icache.scala 29:20]
  reg [52:0] tags1_67; // @[icache.scala 29:20]
  reg [52:0] tags1_68; // @[icache.scala 29:20]
  reg [52:0] tags1_69; // @[icache.scala 29:20]
  reg [52:0] tags1_70; // @[icache.scala 29:20]
  reg [52:0] tags1_71; // @[icache.scala 29:20]
  reg [52:0] tags1_72; // @[icache.scala 29:20]
  reg [52:0] tags1_73; // @[icache.scala 29:20]
  reg [52:0] tags1_74; // @[icache.scala 29:20]
  reg [52:0] tags1_75; // @[icache.scala 29:20]
  reg [52:0] tags1_76; // @[icache.scala 29:20]
  reg [52:0] tags1_77; // @[icache.scala 29:20]
  reg [52:0] tags1_78; // @[icache.scala 29:20]
  reg [52:0] tags1_79; // @[icache.scala 29:20]
  reg [52:0] tags1_80; // @[icache.scala 29:20]
  reg [52:0] tags1_81; // @[icache.scala 29:20]
  reg [52:0] tags1_82; // @[icache.scala 29:20]
  reg [52:0] tags1_83; // @[icache.scala 29:20]
  reg [52:0] tags1_84; // @[icache.scala 29:20]
  reg [52:0] tags1_85; // @[icache.scala 29:20]
  reg [52:0] tags1_86; // @[icache.scala 29:20]
  reg [52:0] tags1_87; // @[icache.scala 29:20]
  reg [52:0] tags1_88; // @[icache.scala 29:20]
  reg [52:0] tags1_89; // @[icache.scala 29:20]
  reg [52:0] tags1_90; // @[icache.scala 29:20]
  reg [52:0] tags1_91; // @[icache.scala 29:20]
  reg [52:0] tags1_92; // @[icache.scala 29:20]
  reg [52:0] tags1_93; // @[icache.scala 29:20]
  reg [52:0] tags1_94; // @[icache.scala 29:20]
  reg [52:0] tags1_95; // @[icache.scala 29:20]
  reg [52:0] tags1_96; // @[icache.scala 29:20]
  reg [52:0] tags1_97; // @[icache.scala 29:20]
  reg [52:0] tags1_98; // @[icache.scala 29:20]
  reg [52:0] tags1_99; // @[icache.scala 29:20]
  reg [52:0] tags1_100; // @[icache.scala 29:20]
  reg [52:0] tags1_101; // @[icache.scala 29:20]
  reg [52:0] tags1_102; // @[icache.scala 29:20]
  reg [52:0] tags1_103; // @[icache.scala 29:20]
  reg [52:0] tags1_104; // @[icache.scala 29:20]
  reg [52:0] tags1_105; // @[icache.scala 29:20]
  reg [52:0] tags1_106; // @[icache.scala 29:20]
  reg [52:0] tags1_107; // @[icache.scala 29:20]
  reg [52:0] tags1_108; // @[icache.scala 29:20]
  reg [52:0] tags1_109; // @[icache.scala 29:20]
  reg [52:0] tags1_110; // @[icache.scala 29:20]
  reg [52:0] tags1_111; // @[icache.scala 29:20]
  reg [52:0] tags1_112; // @[icache.scala 29:20]
  reg [52:0] tags1_113; // @[icache.scala 29:20]
  reg [52:0] tags1_114; // @[icache.scala 29:20]
  reg [52:0] tags1_115; // @[icache.scala 29:20]
  reg [52:0] tags1_116; // @[icache.scala 29:20]
  reg [52:0] tags1_117; // @[icache.scala 29:20]
  reg [52:0] tags1_118; // @[icache.scala 29:20]
  reg [52:0] tags1_119; // @[icache.scala 29:20]
  reg [52:0] tags1_120; // @[icache.scala 29:20]
  reg [52:0] tags1_121; // @[icache.scala 29:20]
  reg [52:0] tags1_122; // @[icache.scala 29:20]
  reg [52:0] tags1_123; // @[icache.scala 29:20]
  reg [52:0] tags1_124; // @[icache.scala 29:20]
  reg [52:0] tags1_125; // @[icache.scala 29:20]
  reg [52:0] tags1_126; // @[icache.scala 29:20]
  reg [52:0] tags1_127; // @[icache.scala 29:20]
  reg  valid0_0; // @[icache.scala 30:21]
  reg  valid0_1; // @[icache.scala 30:21]
  reg  valid0_2; // @[icache.scala 30:21]
  reg  valid0_3; // @[icache.scala 30:21]
  reg  valid0_4; // @[icache.scala 30:21]
  reg  valid0_5; // @[icache.scala 30:21]
  reg  valid0_6; // @[icache.scala 30:21]
  reg  valid0_7; // @[icache.scala 30:21]
  reg  valid0_8; // @[icache.scala 30:21]
  reg  valid0_9; // @[icache.scala 30:21]
  reg  valid0_10; // @[icache.scala 30:21]
  reg  valid0_11; // @[icache.scala 30:21]
  reg  valid0_12; // @[icache.scala 30:21]
  reg  valid0_13; // @[icache.scala 30:21]
  reg  valid0_14; // @[icache.scala 30:21]
  reg  valid0_15; // @[icache.scala 30:21]
  reg  valid0_16; // @[icache.scala 30:21]
  reg  valid0_17; // @[icache.scala 30:21]
  reg  valid0_18; // @[icache.scala 30:21]
  reg  valid0_19; // @[icache.scala 30:21]
  reg  valid0_20; // @[icache.scala 30:21]
  reg  valid0_21; // @[icache.scala 30:21]
  reg  valid0_22; // @[icache.scala 30:21]
  reg  valid0_23; // @[icache.scala 30:21]
  reg  valid0_24; // @[icache.scala 30:21]
  reg  valid0_25; // @[icache.scala 30:21]
  reg  valid0_26; // @[icache.scala 30:21]
  reg  valid0_27; // @[icache.scala 30:21]
  reg  valid0_28; // @[icache.scala 30:21]
  reg  valid0_29; // @[icache.scala 30:21]
  reg  valid0_30; // @[icache.scala 30:21]
  reg  valid0_31; // @[icache.scala 30:21]
  reg  valid0_32; // @[icache.scala 30:21]
  reg  valid0_33; // @[icache.scala 30:21]
  reg  valid0_34; // @[icache.scala 30:21]
  reg  valid0_35; // @[icache.scala 30:21]
  reg  valid0_36; // @[icache.scala 30:21]
  reg  valid0_37; // @[icache.scala 30:21]
  reg  valid0_38; // @[icache.scala 30:21]
  reg  valid0_39; // @[icache.scala 30:21]
  reg  valid0_40; // @[icache.scala 30:21]
  reg  valid0_41; // @[icache.scala 30:21]
  reg  valid0_42; // @[icache.scala 30:21]
  reg  valid0_43; // @[icache.scala 30:21]
  reg  valid0_44; // @[icache.scala 30:21]
  reg  valid0_45; // @[icache.scala 30:21]
  reg  valid0_46; // @[icache.scala 30:21]
  reg  valid0_47; // @[icache.scala 30:21]
  reg  valid0_48; // @[icache.scala 30:21]
  reg  valid0_49; // @[icache.scala 30:21]
  reg  valid0_50; // @[icache.scala 30:21]
  reg  valid0_51; // @[icache.scala 30:21]
  reg  valid0_52; // @[icache.scala 30:21]
  reg  valid0_53; // @[icache.scala 30:21]
  reg  valid0_54; // @[icache.scala 30:21]
  reg  valid0_55; // @[icache.scala 30:21]
  reg  valid0_56; // @[icache.scala 30:21]
  reg  valid0_57; // @[icache.scala 30:21]
  reg  valid0_58; // @[icache.scala 30:21]
  reg  valid0_59; // @[icache.scala 30:21]
  reg  valid0_60; // @[icache.scala 30:21]
  reg  valid0_61; // @[icache.scala 30:21]
  reg  valid0_62; // @[icache.scala 30:21]
  reg  valid0_63; // @[icache.scala 30:21]
  reg  valid0_64; // @[icache.scala 30:21]
  reg  valid0_65; // @[icache.scala 30:21]
  reg  valid0_66; // @[icache.scala 30:21]
  reg  valid0_67; // @[icache.scala 30:21]
  reg  valid0_68; // @[icache.scala 30:21]
  reg  valid0_69; // @[icache.scala 30:21]
  reg  valid0_70; // @[icache.scala 30:21]
  reg  valid0_71; // @[icache.scala 30:21]
  reg  valid0_72; // @[icache.scala 30:21]
  reg  valid0_73; // @[icache.scala 30:21]
  reg  valid0_74; // @[icache.scala 30:21]
  reg  valid0_75; // @[icache.scala 30:21]
  reg  valid0_76; // @[icache.scala 30:21]
  reg  valid0_77; // @[icache.scala 30:21]
  reg  valid0_78; // @[icache.scala 30:21]
  reg  valid0_79; // @[icache.scala 30:21]
  reg  valid0_80; // @[icache.scala 30:21]
  reg  valid0_81; // @[icache.scala 30:21]
  reg  valid0_82; // @[icache.scala 30:21]
  reg  valid0_83; // @[icache.scala 30:21]
  reg  valid0_84; // @[icache.scala 30:21]
  reg  valid0_85; // @[icache.scala 30:21]
  reg  valid0_86; // @[icache.scala 30:21]
  reg  valid0_87; // @[icache.scala 30:21]
  reg  valid0_88; // @[icache.scala 30:21]
  reg  valid0_89; // @[icache.scala 30:21]
  reg  valid0_90; // @[icache.scala 30:21]
  reg  valid0_91; // @[icache.scala 30:21]
  reg  valid0_92; // @[icache.scala 30:21]
  reg  valid0_93; // @[icache.scala 30:21]
  reg  valid0_94; // @[icache.scala 30:21]
  reg  valid0_95; // @[icache.scala 30:21]
  reg  valid0_96; // @[icache.scala 30:21]
  reg  valid0_97; // @[icache.scala 30:21]
  reg  valid0_98; // @[icache.scala 30:21]
  reg  valid0_99; // @[icache.scala 30:21]
  reg  valid0_100; // @[icache.scala 30:21]
  reg  valid0_101; // @[icache.scala 30:21]
  reg  valid0_102; // @[icache.scala 30:21]
  reg  valid0_103; // @[icache.scala 30:21]
  reg  valid0_104; // @[icache.scala 30:21]
  reg  valid0_105; // @[icache.scala 30:21]
  reg  valid0_106; // @[icache.scala 30:21]
  reg  valid0_107; // @[icache.scala 30:21]
  reg  valid0_108; // @[icache.scala 30:21]
  reg  valid0_109; // @[icache.scala 30:21]
  reg  valid0_110; // @[icache.scala 30:21]
  reg  valid0_111; // @[icache.scala 30:21]
  reg  valid0_112; // @[icache.scala 30:21]
  reg  valid0_113; // @[icache.scala 30:21]
  reg  valid0_114; // @[icache.scala 30:21]
  reg  valid0_115; // @[icache.scala 30:21]
  reg  valid0_116; // @[icache.scala 30:21]
  reg  valid0_117; // @[icache.scala 30:21]
  reg  valid0_118; // @[icache.scala 30:21]
  reg  valid0_119; // @[icache.scala 30:21]
  reg  valid0_120; // @[icache.scala 30:21]
  reg  valid0_121; // @[icache.scala 30:21]
  reg  valid0_122; // @[icache.scala 30:21]
  reg  valid0_123; // @[icache.scala 30:21]
  reg  valid0_124; // @[icache.scala 30:21]
  reg  valid0_125; // @[icache.scala 30:21]
  reg  valid0_126; // @[icache.scala 30:21]
  reg  valid0_127; // @[icache.scala 30:21]
  reg  valid1_0; // @[icache.scala 31:21]
  reg  valid1_1; // @[icache.scala 31:21]
  reg  valid1_2; // @[icache.scala 31:21]
  reg  valid1_3; // @[icache.scala 31:21]
  reg  valid1_4; // @[icache.scala 31:21]
  reg  valid1_5; // @[icache.scala 31:21]
  reg  valid1_6; // @[icache.scala 31:21]
  reg  valid1_7; // @[icache.scala 31:21]
  reg  valid1_8; // @[icache.scala 31:21]
  reg  valid1_9; // @[icache.scala 31:21]
  reg  valid1_10; // @[icache.scala 31:21]
  reg  valid1_11; // @[icache.scala 31:21]
  reg  valid1_12; // @[icache.scala 31:21]
  reg  valid1_13; // @[icache.scala 31:21]
  reg  valid1_14; // @[icache.scala 31:21]
  reg  valid1_15; // @[icache.scala 31:21]
  reg  valid1_16; // @[icache.scala 31:21]
  reg  valid1_17; // @[icache.scala 31:21]
  reg  valid1_18; // @[icache.scala 31:21]
  reg  valid1_19; // @[icache.scala 31:21]
  reg  valid1_20; // @[icache.scala 31:21]
  reg  valid1_21; // @[icache.scala 31:21]
  reg  valid1_22; // @[icache.scala 31:21]
  reg  valid1_23; // @[icache.scala 31:21]
  reg  valid1_24; // @[icache.scala 31:21]
  reg  valid1_25; // @[icache.scala 31:21]
  reg  valid1_26; // @[icache.scala 31:21]
  reg  valid1_27; // @[icache.scala 31:21]
  reg  valid1_28; // @[icache.scala 31:21]
  reg  valid1_29; // @[icache.scala 31:21]
  reg  valid1_30; // @[icache.scala 31:21]
  reg  valid1_31; // @[icache.scala 31:21]
  reg  valid1_32; // @[icache.scala 31:21]
  reg  valid1_33; // @[icache.scala 31:21]
  reg  valid1_34; // @[icache.scala 31:21]
  reg  valid1_35; // @[icache.scala 31:21]
  reg  valid1_36; // @[icache.scala 31:21]
  reg  valid1_37; // @[icache.scala 31:21]
  reg  valid1_38; // @[icache.scala 31:21]
  reg  valid1_39; // @[icache.scala 31:21]
  reg  valid1_40; // @[icache.scala 31:21]
  reg  valid1_41; // @[icache.scala 31:21]
  reg  valid1_42; // @[icache.scala 31:21]
  reg  valid1_43; // @[icache.scala 31:21]
  reg  valid1_44; // @[icache.scala 31:21]
  reg  valid1_45; // @[icache.scala 31:21]
  reg  valid1_46; // @[icache.scala 31:21]
  reg  valid1_47; // @[icache.scala 31:21]
  reg  valid1_48; // @[icache.scala 31:21]
  reg  valid1_49; // @[icache.scala 31:21]
  reg  valid1_50; // @[icache.scala 31:21]
  reg  valid1_51; // @[icache.scala 31:21]
  reg  valid1_52; // @[icache.scala 31:21]
  reg  valid1_53; // @[icache.scala 31:21]
  reg  valid1_54; // @[icache.scala 31:21]
  reg  valid1_55; // @[icache.scala 31:21]
  reg  valid1_56; // @[icache.scala 31:21]
  reg  valid1_57; // @[icache.scala 31:21]
  reg  valid1_58; // @[icache.scala 31:21]
  reg  valid1_59; // @[icache.scala 31:21]
  reg  valid1_60; // @[icache.scala 31:21]
  reg  valid1_61; // @[icache.scala 31:21]
  reg  valid1_62; // @[icache.scala 31:21]
  reg  valid1_63; // @[icache.scala 31:21]
  reg  valid1_64; // @[icache.scala 31:21]
  reg  valid1_65; // @[icache.scala 31:21]
  reg  valid1_66; // @[icache.scala 31:21]
  reg  valid1_67; // @[icache.scala 31:21]
  reg  valid1_68; // @[icache.scala 31:21]
  reg  valid1_69; // @[icache.scala 31:21]
  reg  valid1_70; // @[icache.scala 31:21]
  reg  valid1_71; // @[icache.scala 31:21]
  reg  valid1_72; // @[icache.scala 31:21]
  reg  valid1_73; // @[icache.scala 31:21]
  reg  valid1_74; // @[icache.scala 31:21]
  reg  valid1_75; // @[icache.scala 31:21]
  reg  valid1_76; // @[icache.scala 31:21]
  reg  valid1_77; // @[icache.scala 31:21]
  reg  valid1_78; // @[icache.scala 31:21]
  reg  valid1_79; // @[icache.scala 31:21]
  reg  valid1_80; // @[icache.scala 31:21]
  reg  valid1_81; // @[icache.scala 31:21]
  reg  valid1_82; // @[icache.scala 31:21]
  reg  valid1_83; // @[icache.scala 31:21]
  reg  valid1_84; // @[icache.scala 31:21]
  reg  valid1_85; // @[icache.scala 31:21]
  reg  valid1_86; // @[icache.scala 31:21]
  reg  valid1_87; // @[icache.scala 31:21]
  reg  valid1_88; // @[icache.scala 31:21]
  reg  valid1_89; // @[icache.scala 31:21]
  reg  valid1_90; // @[icache.scala 31:21]
  reg  valid1_91; // @[icache.scala 31:21]
  reg  valid1_92; // @[icache.scala 31:21]
  reg  valid1_93; // @[icache.scala 31:21]
  reg  valid1_94; // @[icache.scala 31:21]
  reg  valid1_95; // @[icache.scala 31:21]
  reg  valid1_96; // @[icache.scala 31:21]
  reg  valid1_97; // @[icache.scala 31:21]
  reg  valid1_98; // @[icache.scala 31:21]
  reg  valid1_99; // @[icache.scala 31:21]
  reg  valid1_100; // @[icache.scala 31:21]
  reg  valid1_101; // @[icache.scala 31:21]
  reg  valid1_102; // @[icache.scala 31:21]
  reg  valid1_103; // @[icache.scala 31:21]
  reg  valid1_104; // @[icache.scala 31:21]
  reg  valid1_105; // @[icache.scala 31:21]
  reg  valid1_106; // @[icache.scala 31:21]
  reg  valid1_107; // @[icache.scala 31:21]
  reg  valid1_108; // @[icache.scala 31:21]
  reg  valid1_109; // @[icache.scala 31:21]
  reg  valid1_110; // @[icache.scala 31:21]
  reg  valid1_111; // @[icache.scala 31:21]
  reg  valid1_112; // @[icache.scala 31:21]
  reg  valid1_113; // @[icache.scala 31:21]
  reg  valid1_114; // @[icache.scala 31:21]
  reg  valid1_115; // @[icache.scala 31:21]
  reg  valid1_116; // @[icache.scala 31:21]
  reg  valid1_117; // @[icache.scala 31:21]
  reg  valid1_118; // @[icache.scala 31:21]
  reg  valid1_119; // @[icache.scala 31:21]
  reg  valid1_120; // @[icache.scala 31:21]
  reg  valid1_121; // @[icache.scala 31:21]
  reg  valid1_122; // @[icache.scala 31:21]
  reg  valid1_123; // @[icache.scala 31:21]
  reg  valid1_124; // @[icache.scala 31:21]
  reg  valid1_125; // @[icache.scala 31:21]
  reg  valid1_126; // @[icache.scala 31:21]
  reg  valid1_127; // @[icache.scala 31:21]
  reg [1:0] state; // @[icache.scala 43:20]
  reg  last_stall; // @[icache.scala 64:25]
  reg [127:0] out_reg; // @[icache.scala 65:22]
  wire [6:0] index2 = cpu_if2_o_addr[10:4]; // @[icache.scala 91:25]
  wire  _GEN_644 = 7'h1 == index2 ? valid0_1 : valid0_0; // @[icache.scala 80:{33,33}]
  wire  _GEN_645 = 7'h2 == index2 ? valid0_2 : _GEN_644; // @[icache.scala 80:{33,33}]
  wire  _GEN_646 = 7'h3 == index2 ? valid0_3 : _GEN_645; // @[icache.scala 80:{33,33}]
  wire  _GEN_647 = 7'h4 == index2 ? valid0_4 : _GEN_646; // @[icache.scala 80:{33,33}]
  wire  _GEN_648 = 7'h5 == index2 ? valid0_5 : _GEN_647; // @[icache.scala 80:{33,33}]
  wire  _GEN_649 = 7'h6 == index2 ? valid0_6 : _GEN_648; // @[icache.scala 80:{33,33}]
  wire  _GEN_650 = 7'h7 == index2 ? valid0_7 : _GEN_649; // @[icache.scala 80:{33,33}]
  wire  _GEN_651 = 7'h8 == index2 ? valid0_8 : _GEN_650; // @[icache.scala 80:{33,33}]
  wire  _GEN_652 = 7'h9 == index2 ? valid0_9 : _GEN_651; // @[icache.scala 80:{33,33}]
  wire  _GEN_653 = 7'ha == index2 ? valid0_10 : _GEN_652; // @[icache.scala 80:{33,33}]
  wire  _GEN_654 = 7'hb == index2 ? valid0_11 : _GEN_653; // @[icache.scala 80:{33,33}]
  wire  _GEN_655 = 7'hc == index2 ? valid0_12 : _GEN_654; // @[icache.scala 80:{33,33}]
  wire  _GEN_656 = 7'hd == index2 ? valid0_13 : _GEN_655; // @[icache.scala 80:{33,33}]
  wire  _GEN_657 = 7'he == index2 ? valid0_14 : _GEN_656; // @[icache.scala 80:{33,33}]
  wire  _GEN_658 = 7'hf == index2 ? valid0_15 : _GEN_657; // @[icache.scala 80:{33,33}]
  wire  _GEN_659 = 7'h10 == index2 ? valid0_16 : _GEN_658; // @[icache.scala 80:{33,33}]
  wire  _GEN_660 = 7'h11 == index2 ? valid0_17 : _GEN_659; // @[icache.scala 80:{33,33}]
  wire  _GEN_661 = 7'h12 == index2 ? valid0_18 : _GEN_660; // @[icache.scala 80:{33,33}]
  wire  _GEN_662 = 7'h13 == index2 ? valid0_19 : _GEN_661; // @[icache.scala 80:{33,33}]
  wire  _GEN_663 = 7'h14 == index2 ? valid0_20 : _GEN_662; // @[icache.scala 80:{33,33}]
  wire  _GEN_664 = 7'h15 == index2 ? valid0_21 : _GEN_663; // @[icache.scala 80:{33,33}]
  wire  _GEN_665 = 7'h16 == index2 ? valid0_22 : _GEN_664; // @[icache.scala 80:{33,33}]
  wire  _GEN_666 = 7'h17 == index2 ? valid0_23 : _GEN_665; // @[icache.scala 80:{33,33}]
  wire  _GEN_667 = 7'h18 == index2 ? valid0_24 : _GEN_666; // @[icache.scala 80:{33,33}]
  wire  _GEN_668 = 7'h19 == index2 ? valid0_25 : _GEN_667; // @[icache.scala 80:{33,33}]
  wire  _GEN_669 = 7'h1a == index2 ? valid0_26 : _GEN_668; // @[icache.scala 80:{33,33}]
  wire  _GEN_670 = 7'h1b == index2 ? valid0_27 : _GEN_669; // @[icache.scala 80:{33,33}]
  wire  _GEN_671 = 7'h1c == index2 ? valid0_28 : _GEN_670; // @[icache.scala 80:{33,33}]
  wire  _GEN_672 = 7'h1d == index2 ? valid0_29 : _GEN_671; // @[icache.scala 80:{33,33}]
  wire  _GEN_673 = 7'h1e == index2 ? valid0_30 : _GEN_672; // @[icache.scala 80:{33,33}]
  wire  _GEN_674 = 7'h1f == index2 ? valid0_31 : _GEN_673; // @[icache.scala 80:{33,33}]
  wire  _GEN_675 = 7'h20 == index2 ? valid0_32 : _GEN_674; // @[icache.scala 80:{33,33}]
  wire  _GEN_676 = 7'h21 == index2 ? valid0_33 : _GEN_675; // @[icache.scala 80:{33,33}]
  wire  _GEN_677 = 7'h22 == index2 ? valid0_34 : _GEN_676; // @[icache.scala 80:{33,33}]
  wire  _GEN_678 = 7'h23 == index2 ? valid0_35 : _GEN_677; // @[icache.scala 80:{33,33}]
  wire  _GEN_679 = 7'h24 == index2 ? valid0_36 : _GEN_678; // @[icache.scala 80:{33,33}]
  wire  _GEN_680 = 7'h25 == index2 ? valid0_37 : _GEN_679; // @[icache.scala 80:{33,33}]
  wire  _GEN_681 = 7'h26 == index2 ? valid0_38 : _GEN_680; // @[icache.scala 80:{33,33}]
  wire  _GEN_682 = 7'h27 == index2 ? valid0_39 : _GEN_681; // @[icache.scala 80:{33,33}]
  wire  _GEN_683 = 7'h28 == index2 ? valid0_40 : _GEN_682; // @[icache.scala 80:{33,33}]
  wire  _GEN_684 = 7'h29 == index2 ? valid0_41 : _GEN_683; // @[icache.scala 80:{33,33}]
  wire  _GEN_685 = 7'h2a == index2 ? valid0_42 : _GEN_684; // @[icache.scala 80:{33,33}]
  wire  _GEN_686 = 7'h2b == index2 ? valid0_43 : _GEN_685; // @[icache.scala 80:{33,33}]
  wire  _GEN_687 = 7'h2c == index2 ? valid0_44 : _GEN_686; // @[icache.scala 80:{33,33}]
  wire  _GEN_688 = 7'h2d == index2 ? valid0_45 : _GEN_687; // @[icache.scala 80:{33,33}]
  wire  _GEN_689 = 7'h2e == index2 ? valid0_46 : _GEN_688; // @[icache.scala 80:{33,33}]
  wire  _GEN_690 = 7'h2f == index2 ? valid0_47 : _GEN_689; // @[icache.scala 80:{33,33}]
  wire  _GEN_691 = 7'h30 == index2 ? valid0_48 : _GEN_690; // @[icache.scala 80:{33,33}]
  wire  _GEN_692 = 7'h31 == index2 ? valid0_49 : _GEN_691; // @[icache.scala 80:{33,33}]
  wire  _GEN_693 = 7'h32 == index2 ? valid0_50 : _GEN_692; // @[icache.scala 80:{33,33}]
  wire  _GEN_694 = 7'h33 == index2 ? valid0_51 : _GEN_693; // @[icache.scala 80:{33,33}]
  wire  _GEN_695 = 7'h34 == index2 ? valid0_52 : _GEN_694; // @[icache.scala 80:{33,33}]
  wire  _GEN_696 = 7'h35 == index2 ? valid0_53 : _GEN_695; // @[icache.scala 80:{33,33}]
  wire  _GEN_697 = 7'h36 == index2 ? valid0_54 : _GEN_696; // @[icache.scala 80:{33,33}]
  wire  _GEN_698 = 7'h37 == index2 ? valid0_55 : _GEN_697; // @[icache.scala 80:{33,33}]
  wire  _GEN_699 = 7'h38 == index2 ? valid0_56 : _GEN_698; // @[icache.scala 80:{33,33}]
  wire  _GEN_700 = 7'h39 == index2 ? valid0_57 : _GEN_699; // @[icache.scala 80:{33,33}]
  wire  _GEN_701 = 7'h3a == index2 ? valid0_58 : _GEN_700; // @[icache.scala 80:{33,33}]
  wire  _GEN_702 = 7'h3b == index2 ? valid0_59 : _GEN_701; // @[icache.scala 80:{33,33}]
  wire  _GEN_703 = 7'h3c == index2 ? valid0_60 : _GEN_702; // @[icache.scala 80:{33,33}]
  wire  _GEN_704 = 7'h3d == index2 ? valid0_61 : _GEN_703; // @[icache.scala 80:{33,33}]
  wire  _GEN_705 = 7'h3e == index2 ? valid0_62 : _GEN_704; // @[icache.scala 80:{33,33}]
  wire  _GEN_706 = 7'h3f == index2 ? valid0_63 : _GEN_705; // @[icache.scala 80:{33,33}]
  wire  _GEN_707 = 7'h40 == index2 ? valid0_64 : _GEN_706; // @[icache.scala 80:{33,33}]
  wire  _GEN_708 = 7'h41 == index2 ? valid0_65 : _GEN_707; // @[icache.scala 80:{33,33}]
  wire  _GEN_709 = 7'h42 == index2 ? valid0_66 : _GEN_708; // @[icache.scala 80:{33,33}]
  wire  _GEN_710 = 7'h43 == index2 ? valid0_67 : _GEN_709; // @[icache.scala 80:{33,33}]
  wire  _GEN_711 = 7'h44 == index2 ? valid0_68 : _GEN_710; // @[icache.scala 80:{33,33}]
  wire  _GEN_712 = 7'h45 == index2 ? valid0_69 : _GEN_711; // @[icache.scala 80:{33,33}]
  wire  _GEN_713 = 7'h46 == index2 ? valid0_70 : _GEN_712; // @[icache.scala 80:{33,33}]
  wire  _GEN_714 = 7'h47 == index2 ? valid0_71 : _GEN_713; // @[icache.scala 80:{33,33}]
  wire  _GEN_715 = 7'h48 == index2 ? valid0_72 : _GEN_714; // @[icache.scala 80:{33,33}]
  wire  _GEN_716 = 7'h49 == index2 ? valid0_73 : _GEN_715; // @[icache.scala 80:{33,33}]
  wire  _GEN_717 = 7'h4a == index2 ? valid0_74 : _GEN_716; // @[icache.scala 80:{33,33}]
  wire  _GEN_718 = 7'h4b == index2 ? valid0_75 : _GEN_717; // @[icache.scala 80:{33,33}]
  wire  _GEN_719 = 7'h4c == index2 ? valid0_76 : _GEN_718; // @[icache.scala 80:{33,33}]
  wire  _GEN_720 = 7'h4d == index2 ? valid0_77 : _GEN_719; // @[icache.scala 80:{33,33}]
  wire  _GEN_721 = 7'h4e == index2 ? valid0_78 : _GEN_720; // @[icache.scala 80:{33,33}]
  wire  _GEN_722 = 7'h4f == index2 ? valid0_79 : _GEN_721; // @[icache.scala 80:{33,33}]
  wire  _GEN_723 = 7'h50 == index2 ? valid0_80 : _GEN_722; // @[icache.scala 80:{33,33}]
  wire  _GEN_724 = 7'h51 == index2 ? valid0_81 : _GEN_723; // @[icache.scala 80:{33,33}]
  wire  _GEN_725 = 7'h52 == index2 ? valid0_82 : _GEN_724; // @[icache.scala 80:{33,33}]
  wire  _GEN_726 = 7'h53 == index2 ? valid0_83 : _GEN_725; // @[icache.scala 80:{33,33}]
  wire  _GEN_727 = 7'h54 == index2 ? valid0_84 : _GEN_726; // @[icache.scala 80:{33,33}]
  wire  _GEN_728 = 7'h55 == index2 ? valid0_85 : _GEN_727; // @[icache.scala 80:{33,33}]
  wire  _GEN_729 = 7'h56 == index2 ? valid0_86 : _GEN_728; // @[icache.scala 80:{33,33}]
  wire  _GEN_730 = 7'h57 == index2 ? valid0_87 : _GEN_729; // @[icache.scala 80:{33,33}]
  wire  _GEN_731 = 7'h58 == index2 ? valid0_88 : _GEN_730; // @[icache.scala 80:{33,33}]
  wire  _GEN_732 = 7'h59 == index2 ? valid0_89 : _GEN_731; // @[icache.scala 80:{33,33}]
  wire  _GEN_733 = 7'h5a == index2 ? valid0_90 : _GEN_732; // @[icache.scala 80:{33,33}]
  wire  _GEN_734 = 7'h5b == index2 ? valid0_91 : _GEN_733; // @[icache.scala 80:{33,33}]
  wire  _GEN_735 = 7'h5c == index2 ? valid0_92 : _GEN_734; // @[icache.scala 80:{33,33}]
  wire  _GEN_736 = 7'h5d == index2 ? valid0_93 : _GEN_735; // @[icache.scala 80:{33,33}]
  wire  _GEN_737 = 7'h5e == index2 ? valid0_94 : _GEN_736; // @[icache.scala 80:{33,33}]
  wire  _GEN_738 = 7'h5f == index2 ? valid0_95 : _GEN_737; // @[icache.scala 80:{33,33}]
  wire  _GEN_739 = 7'h60 == index2 ? valid0_96 : _GEN_738; // @[icache.scala 80:{33,33}]
  wire  _GEN_740 = 7'h61 == index2 ? valid0_97 : _GEN_739; // @[icache.scala 80:{33,33}]
  wire  _GEN_741 = 7'h62 == index2 ? valid0_98 : _GEN_740; // @[icache.scala 80:{33,33}]
  wire  _GEN_742 = 7'h63 == index2 ? valid0_99 : _GEN_741; // @[icache.scala 80:{33,33}]
  wire  _GEN_743 = 7'h64 == index2 ? valid0_100 : _GEN_742; // @[icache.scala 80:{33,33}]
  wire  _GEN_744 = 7'h65 == index2 ? valid0_101 : _GEN_743; // @[icache.scala 80:{33,33}]
  wire  _GEN_745 = 7'h66 == index2 ? valid0_102 : _GEN_744; // @[icache.scala 80:{33,33}]
  wire  _GEN_746 = 7'h67 == index2 ? valid0_103 : _GEN_745; // @[icache.scala 80:{33,33}]
  wire  _GEN_747 = 7'h68 == index2 ? valid0_104 : _GEN_746; // @[icache.scala 80:{33,33}]
  wire  _GEN_748 = 7'h69 == index2 ? valid0_105 : _GEN_747; // @[icache.scala 80:{33,33}]
  wire  _GEN_749 = 7'h6a == index2 ? valid0_106 : _GEN_748; // @[icache.scala 80:{33,33}]
  wire  _GEN_750 = 7'h6b == index2 ? valid0_107 : _GEN_749; // @[icache.scala 80:{33,33}]
  wire  _GEN_751 = 7'h6c == index2 ? valid0_108 : _GEN_750; // @[icache.scala 80:{33,33}]
  wire  _GEN_752 = 7'h6d == index2 ? valid0_109 : _GEN_751; // @[icache.scala 80:{33,33}]
  wire  _GEN_753 = 7'h6e == index2 ? valid0_110 : _GEN_752; // @[icache.scala 80:{33,33}]
  wire  _GEN_754 = 7'h6f == index2 ? valid0_111 : _GEN_753; // @[icache.scala 80:{33,33}]
  wire  _GEN_755 = 7'h70 == index2 ? valid0_112 : _GEN_754; // @[icache.scala 80:{33,33}]
  wire  _GEN_756 = 7'h71 == index2 ? valid0_113 : _GEN_755; // @[icache.scala 80:{33,33}]
  wire  _GEN_757 = 7'h72 == index2 ? valid0_114 : _GEN_756; // @[icache.scala 80:{33,33}]
  wire  _GEN_758 = 7'h73 == index2 ? valid0_115 : _GEN_757; // @[icache.scala 80:{33,33}]
  wire  _GEN_759 = 7'h74 == index2 ? valid0_116 : _GEN_758; // @[icache.scala 80:{33,33}]
  wire  _GEN_760 = 7'h75 == index2 ? valid0_117 : _GEN_759; // @[icache.scala 80:{33,33}]
  wire  _GEN_761 = 7'h76 == index2 ? valid0_118 : _GEN_760; // @[icache.scala 80:{33,33}]
  wire  _GEN_762 = 7'h77 == index2 ? valid0_119 : _GEN_761; // @[icache.scala 80:{33,33}]
  wire  _GEN_763 = 7'h78 == index2 ? valid0_120 : _GEN_762; // @[icache.scala 80:{33,33}]
  wire  _GEN_764 = 7'h79 == index2 ? valid0_121 : _GEN_763; // @[icache.scala 80:{33,33}]
  wire  _GEN_765 = 7'h7a == index2 ? valid0_122 : _GEN_764; // @[icache.scala 80:{33,33}]
  wire  _GEN_766 = 7'h7b == index2 ? valid0_123 : _GEN_765; // @[icache.scala 80:{33,33}]
  wire  _GEN_767 = 7'h7c == index2 ? valid0_124 : _GEN_766; // @[icache.scala 80:{33,33}]
  wire  _GEN_768 = 7'h7d == index2 ? valid0_125 : _GEN_767; // @[icache.scala 80:{33,33}]
  wire  _GEN_769 = 7'h7e == index2 ? valid0_126 : _GEN_768; // @[icache.scala 80:{33,33}]
  wire  _GEN_770 = 7'h7f == index2 ? valid0_127 : _GEN_769; // @[icache.scala 80:{33,33}]
  wire [52:0] _GEN_516 = 7'h1 == index2 ? tags0_1 : tags0_0; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_517 = 7'h2 == index2 ? tags0_2 : _GEN_516; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_518 = 7'h3 == index2 ? tags0_3 : _GEN_517; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_519 = 7'h4 == index2 ? tags0_4 : _GEN_518; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_520 = 7'h5 == index2 ? tags0_5 : _GEN_519; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_521 = 7'h6 == index2 ? tags0_6 : _GEN_520; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_522 = 7'h7 == index2 ? tags0_7 : _GEN_521; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_523 = 7'h8 == index2 ? tags0_8 : _GEN_522; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_524 = 7'h9 == index2 ? tags0_9 : _GEN_523; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_525 = 7'ha == index2 ? tags0_10 : _GEN_524; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_526 = 7'hb == index2 ? tags0_11 : _GEN_525; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_527 = 7'hc == index2 ? tags0_12 : _GEN_526; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_528 = 7'hd == index2 ? tags0_13 : _GEN_527; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_529 = 7'he == index2 ? tags0_14 : _GEN_528; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_530 = 7'hf == index2 ? tags0_15 : _GEN_529; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_531 = 7'h10 == index2 ? tags0_16 : _GEN_530; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_532 = 7'h11 == index2 ? tags0_17 : _GEN_531; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_533 = 7'h12 == index2 ? tags0_18 : _GEN_532; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_534 = 7'h13 == index2 ? tags0_19 : _GEN_533; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_535 = 7'h14 == index2 ? tags0_20 : _GEN_534; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_536 = 7'h15 == index2 ? tags0_21 : _GEN_535; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_537 = 7'h16 == index2 ? tags0_22 : _GEN_536; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_538 = 7'h17 == index2 ? tags0_23 : _GEN_537; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_539 = 7'h18 == index2 ? tags0_24 : _GEN_538; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_540 = 7'h19 == index2 ? tags0_25 : _GEN_539; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_541 = 7'h1a == index2 ? tags0_26 : _GEN_540; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_542 = 7'h1b == index2 ? tags0_27 : _GEN_541; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_543 = 7'h1c == index2 ? tags0_28 : _GEN_542; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_544 = 7'h1d == index2 ? tags0_29 : _GEN_543; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_545 = 7'h1e == index2 ? tags0_30 : _GEN_544; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_546 = 7'h1f == index2 ? tags0_31 : _GEN_545; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_547 = 7'h20 == index2 ? tags0_32 : _GEN_546; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_548 = 7'h21 == index2 ? tags0_33 : _GEN_547; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_549 = 7'h22 == index2 ? tags0_34 : _GEN_548; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_550 = 7'h23 == index2 ? tags0_35 : _GEN_549; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_551 = 7'h24 == index2 ? tags0_36 : _GEN_550; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_552 = 7'h25 == index2 ? tags0_37 : _GEN_551; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_553 = 7'h26 == index2 ? tags0_38 : _GEN_552; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_554 = 7'h27 == index2 ? tags0_39 : _GEN_553; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_555 = 7'h28 == index2 ? tags0_40 : _GEN_554; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_556 = 7'h29 == index2 ? tags0_41 : _GEN_555; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_557 = 7'h2a == index2 ? tags0_42 : _GEN_556; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_558 = 7'h2b == index2 ? tags0_43 : _GEN_557; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_559 = 7'h2c == index2 ? tags0_44 : _GEN_558; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_560 = 7'h2d == index2 ? tags0_45 : _GEN_559; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_561 = 7'h2e == index2 ? tags0_46 : _GEN_560; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_562 = 7'h2f == index2 ? tags0_47 : _GEN_561; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_563 = 7'h30 == index2 ? tags0_48 : _GEN_562; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_564 = 7'h31 == index2 ? tags0_49 : _GEN_563; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_565 = 7'h32 == index2 ? tags0_50 : _GEN_564; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_566 = 7'h33 == index2 ? tags0_51 : _GEN_565; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_567 = 7'h34 == index2 ? tags0_52 : _GEN_566; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_568 = 7'h35 == index2 ? tags0_53 : _GEN_567; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_569 = 7'h36 == index2 ? tags0_54 : _GEN_568; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_570 = 7'h37 == index2 ? tags0_55 : _GEN_569; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_571 = 7'h38 == index2 ? tags0_56 : _GEN_570; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_572 = 7'h39 == index2 ? tags0_57 : _GEN_571; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_573 = 7'h3a == index2 ? tags0_58 : _GEN_572; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_574 = 7'h3b == index2 ? tags0_59 : _GEN_573; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_575 = 7'h3c == index2 ? tags0_60 : _GEN_574; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_576 = 7'h3d == index2 ? tags0_61 : _GEN_575; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_577 = 7'h3e == index2 ? tags0_62 : _GEN_576; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_578 = 7'h3f == index2 ? tags0_63 : _GEN_577; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_579 = 7'h40 == index2 ? tags0_64 : _GEN_578; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_580 = 7'h41 == index2 ? tags0_65 : _GEN_579; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_581 = 7'h42 == index2 ? tags0_66 : _GEN_580; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_582 = 7'h43 == index2 ? tags0_67 : _GEN_581; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_583 = 7'h44 == index2 ? tags0_68 : _GEN_582; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_584 = 7'h45 == index2 ? tags0_69 : _GEN_583; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_585 = 7'h46 == index2 ? tags0_70 : _GEN_584; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_586 = 7'h47 == index2 ? tags0_71 : _GEN_585; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_587 = 7'h48 == index2 ? tags0_72 : _GEN_586; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_588 = 7'h49 == index2 ? tags0_73 : _GEN_587; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_589 = 7'h4a == index2 ? tags0_74 : _GEN_588; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_590 = 7'h4b == index2 ? tags0_75 : _GEN_589; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_591 = 7'h4c == index2 ? tags0_76 : _GEN_590; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_592 = 7'h4d == index2 ? tags0_77 : _GEN_591; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_593 = 7'h4e == index2 ? tags0_78 : _GEN_592; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_594 = 7'h4f == index2 ? tags0_79 : _GEN_593; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_595 = 7'h50 == index2 ? tags0_80 : _GEN_594; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_596 = 7'h51 == index2 ? tags0_81 : _GEN_595; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_597 = 7'h52 == index2 ? tags0_82 : _GEN_596; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_598 = 7'h53 == index2 ? tags0_83 : _GEN_597; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_599 = 7'h54 == index2 ? tags0_84 : _GEN_598; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_600 = 7'h55 == index2 ? tags0_85 : _GEN_599; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_601 = 7'h56 == index2 ? tags0_86 : _GEN_600; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_602 = 7'h57 == index2 ? tags0_87 : _GEN_601; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_603 = 7'h58 == index2 ? tags0_88 : _GEN_602; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_604 = 7'h59 == index2 ? tags0_89 : _GEN_603; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_605 = 7'h5a == index2 ? tags0_90 : _GEN_604; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_606 = 7'h5b == index2 ? tags0_91 : _GEN_605; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_607 = 7'h5c == index2 ? tags0_92 : _GEN_606; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_608 = 7'h5d == index2 ? tags0_93 : _GEN_607; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_609 = 7'h5e == index2 ? tags0_94 : _GEN_608; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_610 = 7'h5f == index2 ? tags0_95 : _GEN_609; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_611 = 7'h60 == index2 ? tags0_96 : _GEN_610; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_612 = 7'h61 == index2 ? tags0_97 : _GEN_611; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_613 = 7'h62 == index2 ? tags0_98 : _GEN_612; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_614 = 7'h63 == index2 ? tags0_99 : _GEN_613; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_615 = 7'h64 == index2 ? tags0_100 : _GEN_614; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_616 = 7'h65 == index2 ? tags0_101 : _GEN_615; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_617 = 7'h66 == index2 ? tags0_102 : _GEN_616; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_618 = 7'h67 == index2 ? tags0_103 : _GEN_617; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_619 = 7'h68 == index2 ? tags0_104 : _GEN_618; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_620 = 7'h69 == index2 ? tags0_105 : _GEN_619; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_621 = 7'h6a == index2 ? tags0_106 : _GEN_620; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_622 = 7'h6b == index2 ? tags0_107 : _GEN_621; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_623 = 7'h6c == index2 ? tags0_108 : _GEN_622; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_624 = 7'h6d == index2 ? tags0_109 : _GEN_623; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_625 = 7'h6e == index2 ? tags0_110 : _GEN_624; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_626 = 7'h6f == index2 ? tags0_111 : _GEN_625; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_627 = 7'h70 == index2 ? tags0_112 : _GEN_626; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_628 = 7'h71 == index2 ? tags0_113 : _GEN_627; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_629 = 7'h72 == index2 ? tags0_114 : _GEN_628; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_630 = 7'h73 == index2 ? tags0_115 : _GEN_629; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_631 = 7'h74 == index2 ? tags0_116 : _GEN_630; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_632 = 7'h75 == index2 ? tags0_117 : _GEN_631; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_633 = 7'h76 == index2 ? tags0_118 : _GEN_632; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_634 = 7'h77 == index2 ? tags0_119 : _GEN_633; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_635 = 7'h78 == index2 ? tags0_120 : _GEN_634; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_636 = 7'h79 == index2 ? tags0_121 : _GEN_635; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_637 = 7'h7a == index2 ? tags0_122 : _GEN_636; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_638 = 7'h7b == index2 ? tags0_123 : _GEN_637; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_639 = 7'h7c == index2 ? tags0_124 : _GEN_638; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_640 = 7'h7d == index2 ? tags0_125 : _GEN_639; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_641 = 7'h7e == index2 ? tags0_126 : _GEN_640; // @[icache.scala 80:{50,50}]
  wire [52:0] _GEN_642 = 7'h7f == index2 ? tags0_127 : _GEN_641; // @[icache.scala 80:{50,50}]
  wire [52:0] tag = cpu_if1_o_addr[63:11]; // @[icache.scala 75:22]
  wire  hit_bank2_0 = _GEN_770 & _GEN_642 == tag; // @[icache.scala 80:33]
  wire [127:0] dout = hit_bank2_0 ? data_array_0_io_o_rdata : data_array_1_io_o_rdata; // @[icache.scala 66:15]
  wire [127:0] dout2 = last_stall ? out_reg : dout; // @[icache.scala 67:16]
  wire  _out_reg_T = state == 2'h2; // @[icache.scala 70:21]
  wire [6:0] index = cpu_if1_o_addr[10:4]; // @[icache.scala 76:24]
  wire [52:0] _GEN_4 = 7'h1 == index ? tags0_1 : tags0_0; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_5 = 7'h2 == index ? tags0_2 : _GEN_4; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_6 = 7'h3 == index ? tags0_3 : _GEN_5; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_7 = 7'h4 == index ? tags0_4 : _GEN_6; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_8 = 7'h5 == index ? tags0_5 : _GEN_7; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_9 = 7'h6 == index ? tags0_6 : _GEN_8; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_10 = 7'h7 == index ? tags0_7 : _GEN_9; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_11 = 7'h8 == index ? tags0_8 : _GEN_10; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_12 = 7'h9 == index ? tags0_9 : _GEN_11; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_13 = 7'ha == index ? tags0_10 : _GEN_12; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_14 = 7'hb == index ? tags0_11 : _GEN_13; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_15 = 7'hc == index ? tags0_12 : _GEN_14; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_16 = 7'hd == index ? tags0_13 : _GEN_15; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_17 = 7'he == index ? tags0_14 : _GEN_16; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_18 = 7'hf == index ? tags0_15 : _GEN_17; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_19 = 7'h10 == index ? tags0_16 : _GEN_18; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_20 = 7'h11 == index ? tags0_17 : _GEN_19; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_21 = 7'h12 == index ? tags0_18 : _GEN_20; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_22 = 7'h13 == index ? tags0_19 : _GEN_21; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_23 = 7'h14 == index ? tags0_20 : _GEN_22; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_24 = 7'h15 == index ? tags0_21 : _GEN_23; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_25 = 7'h16 == index ? tags0_22 : _GEN_24; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_26 = 7'h17 == index ? tags0_23 : _GEN_25; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_27 = 7'h18 == index ? tags0_24 : _GEN_26; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_28 = 7'h19 == index ? tags0_25 : _GEN_27; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_29 = 7'h1a == index ? tags0_26 : _GEN_28; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_30 = 7'h1b == index ? tags0_27 : _GEN_29; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_31 = 7'h1c == index ? tags0_28 : _GEN_30; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_32 = 7'h1d == index ? tags0_29 : _GEN_31; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_33 = 7'h1e == index ? tags0_30 : _GEN_32; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_34 = 7'h1f == index ? tags0_31 : _GEN_33; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_35 = 7'h20 == index ? tags0_32 : _GEN_34; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_36 = 7'h21 == index ? tags0_33 : _GEN_35; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_37 = 7'h22 == index ? tags0_34 : _GEN_36; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_38 = 7'h23 == index ? tags0_35 : _GEN_37; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_39 = 7'h24 == index ? tags0_36 : _GEN_38; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_40 = 7'h25 == index ? tags0_37 : _GEN_39; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_41 = 7'h26 == index ? tags0_38 : _GEN_40; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_42 = 7'h27 == index ? tags0_39 : _GEN_41; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_43 = 7'h28 == index ? tags0_40 : _GEN_42; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_44 = 7'h29 == index ? tags0_41 : _GEN_43; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_45 = 7'h2a == index ? tags0_42 : _GEN_44; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_46 = 7'h2b == index ? tags0_43 : _GEN_45; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_47 = 7'h2c == index ? tags0_44 : _GEN_46; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_48 = 7'h2d == index ? tags0_45 : _GEN_47; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_49 = 7'h2e == index ? tags0_46 : _GEN_48; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_50 = 7'h2f == index ? tags0_47 : _GEN_49; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_51 = 7'h30 == index ? tags0_48 : _GEN_50; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_52 = 7'h31 == index ? tags0_49 : _GEN_51; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_53 = 7'h32 == index ? tags0_50 : _GEN_52; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_54 = 7'h33 == index ? tags0_51 : _GEN_53; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_55 = 7'h34 == index ? tags0_52 : _GEN_54; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_56 = 7'h35 == index ? tags0_53 : _GEN_55; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_57 = 7'h36 == index ? tags0_54 : _GEN_56; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_58 = 7'h37 == index ? tags0_55 : _GEN_57; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_59 = 7'h38 == index ? tags0_56 : _GEN_58; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_60 = 7'h39 == index ? tags0_57 : _GEN_59; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_61 = 7'h3a == index ? tags0_58 : _GEN_60; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_62 = 7'h3b == index ? tags0_59 : _GEN_61; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_63 = 7'h3c == index ? tags0_60 : _GEN_62; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_64 = 7'h3d == index ? tags0_61 : _GEN_63; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_65 = 7'h3e == index ? tags0_62 : _GEN_64; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_66 = 7'h3f == index ? tags0_63 : _GEN_65; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_67 = 7'h40 == index ? tags0_64 : _GEN_66; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_68 = 7'h41 == index ? tags0_65 : _GEN_67; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_69 = 7'h42 == index ? tags0_66 : _GEN_68; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_70 = 7'h43 == index ? tags0_67 : _GEN_69; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_71 = 7'h44 == index ? tags0_68 : _GEN_70; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_72 = 7'h45 == index ? tags0_69 : _GEN_71; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_73 = 7'h46 == index ? tags0_70 : _GEN_72; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_74 = 7'h47 == index ? tags0_71 : _GEN_73; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_75 = 7'h48 == index ? tags0_72 : _GEN_74; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_76 = 7'h49 == index ? tags0_73 : _GEN_75; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_77 = 7'h4a == index ? tags0_74 : _GEN_76; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_78 = 7'h4b == index ? tags0_75 : _GEN_77; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_79 = 7'h4c == index ? tags0_76 : _GEN_78; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_80 = 7'h4d == index ? tags0_77 : _GEN_79; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_81 = 7'h4e == index ? tags0_78 : _GEN_80; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_82 = 7'h4f == index ? tags0_79 : _GEN_81; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_83 = 7'h50 == index ? tags0_80 : _GEN_82; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_84 = 7'h51 == index ? tags0_81 : _GEN_83; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_85 = 7'h52 == index ? tags0_82 : _GEN_84; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_86 = 7'h53 == index ? tags0_83 : _GEN_85; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_87 = 7'h54 == index ? tags0_84 : _GEN_86; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_88 = 7'h55 == index ? tags0_85 : _GEN_87; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_89 = 7'h56 == index ? tags0_86 : _GEN_88; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_90 = 7'h57 == index ? tags0_87 : _GEN_89; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_91 = 7'h58 == index ? tags0_88 : _GEN_90; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_92 = 7'h59 == index ? tags0_89 : _GEN_91; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_93 = 7'h5a == index ? tags0_90 : _GEN_92; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_94 = 7'h5b == index ? tags0_91 : _GEN_93; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_95 = 7'h5c == index ? tags0_92 : _GEN_94; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_96 = 7'h5d == index ? tags0_93 : _GEN_95; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_97 = 7'h5e == index ? tags0_94 : _GEN_96; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_98 = 7'h5f == index ? tags0_95 : _GEN_97; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_99 = 7'h60 == index ? tags0_96 : _GEN_98; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_100 = 7'h61 == index ? tags0_97 : _GEN_99; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_101 = 7'h62 == index ? tags0_98 : _GEN_100; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_102 = 7'h63 == index ? tags0_99 : _GEN_101; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_103 = 7'h64 == index ? tags0_100 : _GEN_102; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_104 = 7'h65 == index ? tags0_101 : _GEN_103; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_105 = 7'h66 == index ? tags0_102 : _GEN_104; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_106 = 7'h67 == index ? tags0_103 : _GEN_105; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_107 = 7'h68 == index ? tags0_104 : _GEN_106; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_108 = 7'h69 == index ? tags0_105 : _GEN_107; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_109 = 7'h6a == index ? tags0_106 : _GEN_108; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_110 = 7'h6b == index ? tags0_107 : _GEN_109; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_111 = 7'h6c == index ? tags0_108 : _GEN_110; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_112 = 7'h6d == index ? tags0_109 : _GEN_111; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_113 = 7'h6e == index ? tags0_110 : _GEN_112; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_114 = 7'h6f == index ? tags0_111 : _GEN_113; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_115 = 7'h70 == index ? tags0_112 : _GEN_114; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_116 = 7'h71 == index ? tags0_113 : _GEN_115; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_117 = 7'h72 == index ? tags0_114 : _GEN_116; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_118 = 7'h73 == index ? tags0_115 : _GEN_117; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_119 = 7'h74 == index ? tags0_116 : _GEN_118; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_120 = 7'h75 == index ? tags0_117 : _GEN_119; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_121 = 7'h76 == index ? tags0_118 : _GEN_120; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_122 = 7'h77 == index ? tags0_119 : _GEN_121; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_123 = 7'h78 == index ? tags0_120 : _GEN_122; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_124 = 7'h79 == index ? tags0_121 : _GEN_123; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_125 = 7'h7a == index ? tags0_122 : _GEN_124; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_126 = 7'h7b == index ? tags0_123 : _GEN_125; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_127 = 7'h7c == index ? tags0_124 : _GEN_126; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_128 = 7'h7d == index ? tags0_125 : _GEN_127; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_129 = 7'h7e == index ? tags0_126 : _GEN_128; // @[icache.scala 78:{47,47}]
  wire [52:0] _GEN_130 = 7'h7f == index ? tags0_127 : _GEN_129; // @[icache.scala 78:{47,47}]
  wire  _GEN_132 = 7'h1 == index ? valid0_1 : valid0_0; // @[icache.scala 78:{31,31}]
  wire  _GEN_133 = 7'h2 == index ? valid0_2 : _GEN_132; // @[icache.scala 78:{31,31}]
  wire  _GEN_134 = 7'h3 == index ? valid0_3 : _GEN_133; // @[icache.scala 78:{31,31}]
  wire  _GEN_135 = 7'h4 == index ? valid0_4 : _GEN_134; // @[icache.scala 78:{31,31}]
  wire  _GEN_136 = 7'h5 == index ? valid0_5 : _GEN_135; // @[icache.scala 78:{31,31}]
  wire  _GEN_137 = 7'h6 == index ? valid0_6 : _GEN_136; // @[icache.scala 78:{31,31}]
  wire  _GEN_138 = 7'h7 == index ? valid0_7 : _GEN_137; // @[icache.scala 78:{31,31}]
  wire  _GEN_139 = 7'h8 == index ? valid0_8 : _GEN_138; // @[icache.scala 78:{31,31}]
  wire  _GEN_140 = 7'h9 == index ? valid0_9 : _GEN_139; // @[icache.scala 78:{31,31}]
  wire  _GEN_141 = 7'ha == index ? valid0_10 : _GEN_140; // @[icache.scala 78:{31,31}]
  wire  _GEN_142 = 7'hb == index ? valid0_11 : _GEN_141; // @[icache.scala 78:{31,31}]
  wire  _GEN_143 = 7'hc == index ? valid0_12 : _GEN_142; // @[icache.scala 78:{31,31}]
  wire  _GEN_144 = 7'hd == index ? valid0_13 : _GEN_143; // @[icache.scala 78:{31,31}]
  wire  _GEN_145 = 7'he == index ? valid0_14 : _GEN_144; // @[icache.scala 78:{31,31}]
  wire  _GEN_146 = 7'hf == index ? valid0_15 : _GEN_145; // @[icache.scala 78:{31,31}]
  wire  _GEN_147 = 7'h10 == index ? valid0_16 : _GEN_146; // @[icache.scala 78:{31,31}]
  wire  _GEN_148 = 7'h11 == index ? valid0_17 : _GEN_147; // @[icache.scala 78:{31,31}]
  wire  _GEN_149 = 7'h12 == index ? valid0_18 : _GEN_148; // @[icache.scala 78:{31,31}]
  wire  _GEN_150 = 7'h13 == index ? valid0_19 : _GEN_149; // @[icache.scala 78:{31,31}]
  wire  _GEN_151 = 7'h14 == index ? valid0_20 : _GEN_150; // @[icache.scala 78:{31,31}]
  wire  _GEN_152 = 7'h15 == index ? valid0_21 : _GEN_151; // @[icache.scala 78:{31,31}]
  wire  _GEN_153 = 7'h16 == index ? valid0_22 : _GEN_152; // @[icache.scala 78:{31,31}]
  wire  _GEN_154 = 7'h17 == index ? valid0_23 : _GEN_153; // @[icache.scala 78:{31,31}]
  wire  _GEN_155 = 7'h18 == index ? valid0_24 : _GEN_154; // @[icache.scala 78:{31,31}]
  wire  _GEN_156 = 7'h19 == index ? valid0_25 : _GEN_155; // @[icache.scala 78:{31,31}]
  wire  _GEN_157 = 7'h1a == index ? valid0_26 : _GEN_156; // @[icache.scala 78:{31,31}]
  wire  _GEN_158 = 7'h1b == index ? valid0_27 : _GEN_157; // @[icache.scala 78:{31,31}]
  wire  _GEN_159 = 7'h1c == index ? valid0_28 : _GEN_158; // @[icache.scala 78:{31,31}]
  wire  _GEN_160 = 7'h1d == index ? valid0_29 : _GEN_159; // @[icache.scala 78:{31,31}]
  wire  _GEN_161 = 7'h1e == index ? valid0_30 : _GEN_160; // @[icache.scala 78:{31,31}]
  wire  _GEN_162 = 7'h1f == index ? valid0_31 : _GEN_161; // @[icache.scala 78:{31,31}]
  wire  _GEN_163 = 7'h20 == index ? valid0_32 : _GEN_162; // @[icache.scala 78:{31,31}]
  wire  _GEN_164 = 7'h21 == index ? valid0_33 : _GEN_163; // @[icache.scala 78:{31,31}]
  wire  _GEN_165 = 7'h22 == index ? valid0_34 : _GEN_164; // @[icache.scala 78:{31,31}]
  wire  _GEN_166 = 7'h23 == index ? valid0_35 : _GEN_165; // @[icache.scala 78:{31,31}]
  wire  _GEN_167 = 7'h24 == index ? valid0_36 : _GEN_166; // @[icache.scala 78:{31,31}]
  wire  _GEN_168 = 7'h25 == index ? valid0_37 : _GEN_167; // @[icache.scala 78:{31,31}]
  wire  _GEN_169 = 7'h26 == index ? valid0_38 : _GEN_168; // @[icache.scala 78:{31,31}]
  wire  _GEN_170 = 7'h27 == index ? valid0_39 : _GEN_169; // @[icache.scala 78:{31,31}]
  wire  _GEN_171 = 7'h28 == index ? valid0_40 : _GEN_170; // @[icache.scala 78:{31,31}]
  wire  _GEN_172 = 7'h29 == index ? valid0_41 : _GEN_171; // @[icache.scala 78:{31,31}]
  wire  _GEN_173 = 7'h2a == index ? valid0_42 : _GEN_172; // @[icache.scala 78:{31,31}]
  wire  _GEN_174 = 7'h2b == index ? valid0_43 : _GEN_173; // @[icache.scala 78:{31,31}]
  wire  _GEN_175 = 7'h2c == index ? valid0_44 : _GEN_174; // @[icache.scala 78:{31,31}]
  wire  _GEN_176 = 7'h2d == index ? valid0_45 : _GEN_175; // @[icache.scala 78:{31,31}]
  wire  _GEN_177 = 7'h2e == index ? valid0_46 : _GEN_176; // @[icache.scala 78:{31,31}]
  wire  _GEN_178 = 7'h2f == index ? valid0_47 : _GEN_177; // @[icache.scala 78:{31,31}]
  wire  _GEN_179 = 7'h30 == index ? valid0_48 : _GEN_178; // @[icache.scala 78:{31,31}]
  wire  _GEN_180 = 7'h31 == index ? valid0_49 : _GEN_179; // @[icache.scala 78:{31,31}]
  wire  _GEN_181 = 7'h32 == index ? valid0_50 : _GEN_180; // @[icache.scala 78:{31,31}]
  wire  _GEN_182 = 7'h33 == index ? valid0_51 : _GEN_181; // @[icache.scala 78:{31,31}]
  wire  _GEN_183 = 7'h34 == index ? valid0_52 : _GEN_182; // @[icache.scala 78:{31,31}]
  wire  _GEN_184 = 7'h35 == index ? valid0_53 : _GEN_183; // @[icache.scala 78:{31,31}]
  wire  _GEN_185 = 7'h36 == index ? valid0_54 : _GEN_184; // @[icache.scala 78:{31,31}]
  wire  _GEN_186 = 7'h37 == index ? valid0_55 : _GEN_185; // @[icache.scala 78:{31,31}]
  wire  _GEN_187 = 7'h38 == index ? valid0_56 : _GEN_186; // @[icache.scala 78:{31,31}]
  wire  _GEN_188 = 7'h39 == index ? valid0_57 : _GEN_187; // @[icache.scala 78:{31,31}]
  wire  _GEN_189 = 7'h3a == index ? valid0_58 : _GEN_188; // @[icache.scala 78:{31,31}]
  wire  _GEN_190 = 7'h3b == index ? valid0_59 : _GEN_189; // @[icache.scala 78:{31,31}]
  wire  _GEN_191 = 7'h3c == index ? valid0_60 : _GEN_190; // @[icache.scala 78:{31,31}]
  wire  _GEN_192 = 7'h3d == index ? valid0_61 : _GEN_191; // @[icache.scala 78:{31,31}]
  wire  _GEN_193 = 7'h3e == index ? valid0_62 : _GEN_192; // @[icache.scala 78:{31,31}]
  wire  _GEN_194 = 7'h3f == index ? valid0_63 : _GEN_193; // @[icache.scala 78:{31,31}]
  wire  _GEN_195 = 7'h40 == index ? valid0_64 : _GEN_194; // @[icache.scala 78:{31,31}]
  wire  _GEN_196 = 7'h41 == index ? valid0_65 : _GEN_195; // @[icache.scala 78:{31,31}]
  wire  _GEN_197 = 7'h42 == index ? valid0_66 : _GEN_196; // @[icache.scala 78:{31,31}]
  wire  _GEN_198 = 7'h43 == index ? valid0_67 : _GEN_197; // @[icache.scala 78:{31,31}]
  wire  _GEN_199 = 7'h44 == index ? valid0_68 : _GEN_198; // @[icache.scala 78:{31,31}]
  wire  _GEN_200 = 7'h45 == index ? valid0_69 : _GEN_199; // @[icache.scala 78:{31,31}]
  wire  _GEN_201 = 7'h46 == index ? valid0_70 : _GEN_200; // @[icache.scala 78:{31,31}]
  wire  _GEN_202 = 7'h47 == index ? valid0_71 : _GEN_201; // @[icache.scala 78:{31,31}]
  wire  _GEN_203 = 7'h48 == index ? valid0_72 : _GEN_202; // @[icache.scala 78:{31,31}]
  wire  _GEN_204 = 7'h49 == index ? valid0_73 : _GEN_203; // @[icache.scala 78:{31,31}]
  wire  _GEN_205 = 7'h4a == index ? valid0_74 : _GEN_204; // @[icache.scala 78:{31,31}]
  wire  _GEN_206 = 7'h4b == index ? valid0_75 : _GEN_205; // @[icache.scala 78:{31,31}]
  wire  _GEN_207 = 7'h4c == index ? valid0_76 : _GEN_206; // @[icache.scala 78:{31,31}]
  wire  _GEN_208 = 7'h4d == index ? valid0_77 : _GEN_207; // @[icache.scala 78:{31,31}]
  wire  _GEN_209 = 7'h4e == index ? valid0_78 : _GEN_208; // @[icache.scala 78:{31,31}]
  wire  _GEN_210 = 7'h4f == index ? valid0_79 : _GEN_209; // @[icache.scala 78:{31,31}]
  wire  _GEN_211 = 7'h50 == index ? valid0_80 : _GEN_210; // @[icache.scala 78:{31,31}]
  wire  _GEN_212 = 7'h51 == index ? valid0_81 : _GEN_211; // @[icache.scala 78:{31,31}]
  wire  _GEN_213 = 7'h52 == index ? valid0_82 : _GEN_212; // @[icache.scala 78:{31,31}]
  wire  _GEN_214 = 7'h53 == index ? valid0_83 : _GEN_213; // @[icache.scala 78:{31,31}]
  wire  _GEN_215 = 7'h54 == index ? valid0_84 : _GEN_214; // @[icache.scala 78:{31,31}]
  wire  _GEN_216 = 7'h55 == index ? valid0_85 : _GEN_215; // @[icache.scala 78:{31,31}]
  wire  _GEN_217 = 7'h56 == index ? valid0_86 : _GEN_216; // @[icache.scala 78:{31,31}]
  wire  _GEN_218 = 7'h57 == index ? valid0_87 : _GEN_217; // @[icache.scala 78:{31,31}]
  wire  _GEN_219 = 7'h58 == index ? valid0_88 : _GEN_218; // @[icache.scala 78:{31,31}]
  wire  _GEN_220 = 7'h59 == index ? valid0_89 : _GEN_219; // @[icache.scala 78:{31,31}]
  wire  _GEN_221 = 7'h5a == index ? valid0_90 : _GEN_220; // @[icache.scala 78:{31,31}]
  wire  _GEN_222 = 7'h5b == index ? valid0_91 : _GEN_221; // @[icache.scala 78:{31,31}]
  wire  _GEN_223 = 7'h5c == index ? valid0_92 : _GEN_222; // @[icache.scala 78:{31,31}]
  wire  _GEN_224 = 7'h5d == index ? valid0_93 : _GEN_223; // @[icache.scala 78:{31,31}]
  wire  _GEN_225 = 7'h5e == index ? valid0_94 : _GEN_224; // @[icache.scala 78:{31,31}]
  wire  _GEN_226 = 7'h5f == index ? valid0_95 : _GEN_225; // @[icache.scala 78:{31,31}]
  wire  _GEN_227 = 7'h60 == index ? valid0_96 : _GEN_226; // @[icache.scala 78:{31,31}]
  wire  _GEN_228 = 7'h61 == index ? valid0_97 : _GEN_227; // @[icache.scala 78:{31,31}]
  wire  _GEN_229 = 7'h62 == index ? valid0_98 : _GEN_228; // @[icache.scala 78:{31,31}]
  wire  _GEN_230 = 7'h63 == index ? valid0_99 : _GEN_229; // @[icache.scala 78:{31,31}]
  wire  _GEN_231 = 7'h64 == index ? valid0_100 : _GEN_230; // @[icache.scala 78:{31,31}]
  wire  _GEN_232 = 7'h65 == index ? valid0_101 : _GEN_231; // @[icache.scala 78:{31,31}]
  wire  _GEN_233 = 7'h66 == index ? valid0_102 : _GEN_232; // @[icache.scala 78:{31,31}]
  wire  _GEN_234 = 7'h67 == index ? valid0_103 : _GEN_233; // @[icache.scala 78:{31,31}]
  wire  _GEN_235 = 7'h68 == index ? valid0_104 : _GEN_234; // @[icache.scala 78:{31,31}]
  wire  _GEN_236 = 7'h69 == index ? valid0_105 : _GEN_235; // @[icache.scala 78:{31,31}]
  wire  _GEN_237 = 7'h6a == index ? valid0_106 : _GEN_236; // @[icache.scala 78:{31,31}]
  wire  _GEN_238 = 7'h6b == index ? valid0_107 : _GEN_237; // @[icache.scala 78:{31,31}]
  wire  _GEN_239 = 7'h6c == index ? valid0_108 : _GEN_238; // @[icache.scala 78:{31,31}]
  wire  _GEN_240 = 7'h6d == index ? valid0_109 : _GEN_239; // @[icache.scala 78:{31,31}]
  wire  _GEN_241 = 7'h6e == index ? valid0_110 : _GEN_240; // @[icache.scala 78:{31,31}]
  wire  _GEN_242 = 7'h6f == index ? valid0_111 : _GEN_241; // @[icache.scala 78:{31,31}]
  wire  _GEN_243 = 7'h70 == index ? valid0_112 : _GEN_242; // @[icache.scala 78:{31,31}]
  wire  _GEN_244 = 7'h71 == index ? valid0_113 : _GEN_243; // @[icache.scala 78:{31,31}]
  wire  _GEN_245 = 7'h72 == index ? valid0_114 : _GEN_244; // @[icache.scala 78:{31,31}]
  wire  _GEN_246 = 7'h73 == index ? valid0_115 : _GEN_245; // @[icache.scala 78:{31,31}]
  wire  _GEN_247 = 7'h74 == index ? valid0_116 : _GEN_246; // @[icache.scala 78:{31,31}]
  wire  _GEN_248 = 7'h75 == index ? valid0_117 : _GEN_247; // @[icache.scala 78:{31,31}]
  wire  _GEN_249 = 7'h76 == index ? valid0_118 : _GEN_248; // @[icache.scala 78:{31,31}]
  wire  _GEN_250 = 7'h77 == index ? valid0_119 : _GEN_249; // @[icache.scala 78:{31,31}]
  wire  _GEN_251 = 7'h78 == index ? valid0_120 : _GEN_250; // @[icache.scala 78:{31,31}]
  wire  _GEN_252 = 7'h79 == index ? valid0_121 : _GEN_251; // @[icache.scala 78:{31,31}]
  wire  _GEN_253 = 7'h7a == index ? valid0_122 : _GEN_252; // @[icache.scala 78:{31,31}]
  wire  _GEN_254 = 7'h7b == index ? valid0_123 : _GEN_253; // @[icache.scala 78:{31,31}]
  wire  _GEN_255 = 7'h7c == index ? valid0_124 : _GEN_254; // @[icache.scala 78:{31,31}]
  wire  _GEN_256 = 7'h7d == index ? valid0_125 : _GEN_255; // @[icache.scala 78:{31,31}]
  wire  _GEN_257 = 7'h7e == index ? valid0_126 : _GEN_256; // @[icache.scala 78:{31,31}]
  wire  _GEN_258 = 7'h7f == index ? valid0_127 : _GEN_257; // @[icache.scala 78:{31,31}]
  wire  hit_bank_0 = _GEN_258 & _GEN_130 == tag; // @[icache.scala 78:31]
  wire [52:0] _GEN_260 = 7'h1 == index ? tags1_1 : tags1_0; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_261 = 7'h2 == index ? tags1_2 : _GEN_260; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_262 = 7'h3 == index ? tags1_3 : _GEN_261; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_263 = 7'h4 == index ? tags1_4 : _GEN_262; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_264 = 7'h5 == index ? tags1_5 : _GEN_263; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_265 = 7'h6 == index ? tags1_6 : _GEN_264; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_266 = 7'h7 == index ? tags1_7 : _GEN_265; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_267 = 7'h8 == index ? tags1_8 : _GEN_266; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_268 = 7'h9 == index ? tags1_9 : _GEN_267; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_269 = 7'ha == index ? tags1_10 : _GEN_268; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_270 = 7'hb == index ? tags1_11 : _GEN_269; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_271 = 7'hc == index ? tags1_12 : _GEN_270; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_272 = 7'hd == index ? tags1_13 : _GEN_271; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_273 = 7'he == index ? tags1_14 : _GEN_272; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_274 = 7'hf == index ? tags1_15 : _GEN_273; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_275 = 7'h10 == index ? tags1_16 : _GEN_274; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_276 = 7'h11 == index ? tags1_17 : _GEN_275; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_277 = 7'h12 == index ? tags1_18 : _GEN_276; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_278 = 7'h13 == index ? tags1_19 : _GEN_277; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_279 = 7'h14 == index ? tags1_20 : _GEN_278; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_280 = 7'h15 == index ? tags1_21 : _GEN_279; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_281 = 7'h16 == index ? tags1_22 : _GEN_280; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_282 = 7'h17 == index ? tags1_23 : _GEN_281; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_283 = 7'h18 == index ? tags1_24 : _GEN_282; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_284 = 7'h19 == index ? tags1_25 : _GEN_283; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_285 = 7'h1a == index ? tags1_26 : _GEN_284; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_286 = 7'h1b == index ? tags1_27 : _GEN_285; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_287 = 7'h1c == index ? tags1_28 : _GEN_286; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_288 = 7'h1d == index ? tags1_29 : _GEN_287; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_289 = 7'h1e == index ? tags1_30 : _GEN_288; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_290 = 7'h1f == index ? tags1_31 : _GEN_289; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_291 = 7'h20 == index ? tags1_32 : _GEN_290; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_292 = 7'h21 == index ? tags1_33 : _GEN_291; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_293 = 7'h22 == index ? tags1_34 : _GEN_292; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_294 = 7'h23 == index ? tags1_35 : _GEN_293; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_295 = 7'h24 == index ? tags1_36 : _GEN_294; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_296 = 7'h25 == index ? tags1_37 : _GEN_295; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_297 = 7'h26 == index ? tags1_38 : _GEN_296; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_298 = 7'h27 == index ? tags1_39 : _GEN_297; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_299 = 7'h28 == index ? tags1_40 : _GEN_298; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_300 = 7'h29 == index ? tags1_41 : _GEN_299; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_301 = 7'h2a == index ? tags1_42 : _GEN_300; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_302 = 7'h2b == index ? tags1_43 : _GEN_301; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_303 = 7'h2c == index ? tags1_44 : _GEN_302; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_304 = 7'h2d == index ? tags1_45 : _GEN_303; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_305 = 7'h2e == index ? tags1_46 : _GEN_304; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_306 = 7'h2f == index ? tags1_47 : _GEN_305; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_307 = 7'h30 == index ? tags1_48 : _GEN_306; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_308 = 7'h31 == index ? tags1_49 : _GEN_307; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_309 = 7'h32 == index ? tags1_50 : _GEN_308; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_310 = 7'h33 == index ? tags1_51 : _GEN_309; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_311 = 7'h34 == index ? tags1_52 : _GEN_310; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_312 = 7'h35 == index ? tags1_53 : _GEN_311; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_313 = 7'h36 == index ? tags1_54 : _GEN_312; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_314 = 7'h37 == index ? tags1_55 : _GEN_313; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_315 = 7'h38 == index ? tags1_56 : _GEN_314; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_316 = 7'h39 == index ? tags1_57 : _GEN_315; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_317 = 7'h3a == index ? tags1_58 : _GEN_316; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_318 = 7'h3b == index ? tags1_59 : _GEN_317; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_319 = 7'h3c == index ? tags1_60 : _GEN_318; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_320 = 7'h3d == index ? tags1_61 : _GEN_319; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_321 = 7'h3e == index ? tags1_62 : _GEN_320; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_322 = 7'h3f == index ? tags1_63 : _GEN_321; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_323 = 7'h40 == index ? tags1_64 : _GEN_322; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_324 = 7'h41 == index ? tags1_65 : _GEN_323; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_325 = 7'h42 == index ? tags1_66 : _GEN_324; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_326 = 7'h43 == index ? tags1_67 : _GEN_325; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_327 = 7'h44 == index ? tags1_68 : _GEN_326; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_328 = 7'h45 == index ? tags1_69 : _GEN_327; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_329 = 7'h46 == index ? tags1_70 : _GEN_328; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_330 = 7'h47 == index ? tags1_71 : _GEN_329; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_331 = 7'h48 == index ? tags1_72 : _GEN_330; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_332 = 7'h49 == index ? tags1_73 : _GEN_331; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_333 = 7'h4a == index ? tags1_74 : _GEN_332; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_334 = 7'h4b == index ? tags1_75 : _GEN_333; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_335 = 7'h4c == index ? tags1_76 : _GEN_334; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_336 = 7'h4d == index ? tags1_77 : _GEN_335; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_337 = 7'h4e == index ? tags1_78 : _GEN_336; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_338 = 7'h4f == index ? tags1_79 : _GEN_337; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_339 = 7'h50 == index ? tags1_80 : _GEN_338; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_340 = 7'h51 == index ? tags1_81 : _GEN_339; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_341 = 7'h52 == index ? tags1_82 : _GEN_340; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_342 = 7'h53 == index ? tags1_83 : _GEN_341; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_343 = 7'h54 == index ? tags1_84 : _GEN_342; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_344 = 7'h55 == index ? tags1_85 : _GEN_343; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_345 = 7'h56 == index ? tags1_86 : _GEN_344; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_346 = 7'h57 == index ? tags1_87 : _GEN_345; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_347 = 7'h58 == index ? tags1_88 : _GEN_346; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_348 = 7'h59 == index ? tags1_89 : _GEN_347; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_349 = 7'h5a == index ? tags1_90 : _GEN_348; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_350 = 7'h5b == index ? tags1_91 : _GEN_349; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_351 = 7'h5c == index ? tags1_92 : _GEN_350; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_352 = 7'h5d == index ? tags1_93 : _GEN_351; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_353 = 7'h5e == index ? tags1_94 : _GEN_352; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_354 = 7'h5f == index ? tags1_95 : _GEN_353; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_355 = 7'h60 == index ? tags1_96 : _GEN_354; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_356 = 7'h61 == index ? tags1_97 : _GEN_355; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_357 = 7'h62 == index ? tags1_98 : _GEN_356; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_358 = 7'h63 == index ? tags1_99 : _GEN_357; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_359 = 7'h64 == index ? tags1_100 : _GEN_358; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_360 = 7'h65 == index ? tags1_101 : _GEN_359; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_361 = 7'h66 == index ? tags1_102 : _GEN_360; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_362 = 7'h67 == index ? tags1_103 : _GEN_361; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_363 = 7'h68 == index ? tags1_104 : _GEN_362; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_364 = 7'h69 == index ? tags1_105 : _GEN_363; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_365 = 7'h6a == index ? tags1_106 : _GEN_364; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_366 = 7'h6b == index ? tags1_107 : _GEN_365; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_367 = 7'h6c == index ? tags1_108 : _GEN_366; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_368 = 7'h6d == index ? tags1_109 : _GEN_367; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_369 = 7'h6e == index ? tags1_110 : _GEN_368; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_370 = 7'h6f == index ? tags1_111 : _GEN_369; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_371 = 7'h70 == index ? tags1_112 : _GEN_370; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_372 = 7'h71 == index ? tags1_113 : _GEN_371; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_373 = 7'h72 == index ? tags1_114 : _GEN_372; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_374 = 7'h73 == index ? tags1_115 : _GEN_373; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_375 = 7'h74 == index ? tags1_116 : _GEN_374; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_376 = 7'h75 == index ? tags1_117 : _GEN_375; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_377 = 7'h76 == index ? tags1_118 : _GEN_376; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_378 = 7'h77 == index ? tags1_119 : _GEN_377; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_379 = 7'h78 == index ? tags1_120 : _GEN_378; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_380 = 7'h79 == index ? tags1_121 : _GEN_379; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_381 = 7'h7a == index ? tags1_122 : _GEN_380; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_382 = 7'h7b == index ? tags1_123 : _GEN_381; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_383 = 7'h7c == index ? tags1_124 : _GEN_382; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_384 = 7'h7d == index ? tags1_125 : _GEN_383; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_385 = 7'h7e == index ? tags1_126 : _GEN_384; // @[icache.scala 79:{47,47}]
  wire [52:0] _GEN_386 = 7'h7f == index ? tags1_127 : _GEN_385; // @[icache.scala 79:{47,47}]
  wire  _GEN_388 = 7'h1 == index ? valid1_1 : valid1_0; // @[icache.scala 79:{31,31}]
  wire  _GEN_389 = 7'h2 == index ? valid1_2 : _GEN_388; // @[icache.scala 79:{31,31}]
  wire  _GEN_390 = 7'h3 == index ? valid1_3 : _GEN_389; // @[icache.scala 79:{31,31}]
  wire  _GEN_391 = 7'h4 == index ? valid1_4 : _GEN_390; // @[icache.scala 79:{31,31}]
  wire  _GEN_392 = 7'h5 == index ? valid1_5 : _GEN_391; // @[icache.scala 79:{31,31}]
  wire  _GEN_393 = 7'h6 == index ? valid1_6 : _GEN_392; // @[icache.scala 79:{31,31}]
  wire  _GEN_394 = 7'h7 == index ? valid1_7 : _GEN_393; // @[icache.scala 79:{31,31}]
  wire  _GEN_395 = 7'h8 == index ? valid1_8 : _GEN_394; // @[icache.scala 79:{31,31}]
  wire  _GEN_396 = 7'h9 == index ? valid1_9 : _GEN_395; // @[icache.scala 79:{31,31}]
  wire  _GEN_397 = 7'ha == index ? valid1_10 : _GEN_396; // @[icache.scala 79:{31,31}]
  wire  _GEN_398 = 7'hb == index ? valid1_11 : _GEN_397; // @[icache.scala 79:{31,31}]
  wire  _GEN_399 = 7'hc == index ? valid1_12 : _GEN_398; // @[icache.scala 79:{31,31}]
  wire  _GEN_400 = 7'hd == index ? valid1_13 : _GEN_399; // @[icache.scala 79:{31,31}]
  wire  _GEN_401 = 7'he == index ? valid1_14 : _GEN_400; // @[icache.scala 79:{31,31}]
  wire  _GEN_402 = 7'hf == index ? valid1_15 : _GEN_401; // @[icache.scala 79:{31,31}]
  wire  _GEN_403 = 7'h10 == index ? valid1_16 : _GEN_402; // @[icache.scala 79:{31,31}]
  wire  _GEN_404 = 7'h11 == index ? valid1_17 : _GEN_403; // @[icache.scala 79:{31,31}]
  wire  _GEN_405 = 7'h12 == index ? valid1_18 : _GEN_404; // @[icache.scala 79:{31,31}]
  wire  _GEN_406 = 7'h13 == index ? valid1_19 : _GEN_405; // @[icache.scala 79:{31,31}]
  wire  _GEN_407 = 7'h14 == index ? valid1_20 : _GEN_406; // @[icache.scala 79:{31,31}]
  wire  _GEN_408 = 7'h15 == index ? valid1_21 : _GEN_407; // @[icache.scala 79:{31,31}]
  wire  _GEN_409 = 7'h16 == index ? valid1_22 : _GEN_408; // @[icache.scala 79:{31,31}]
  wire  _GEN_410 = 7'h17 == index ? valid1_23 : _GEN_409; // @[icache.scala 79:{31,31}]
  wire  _GEN_411 = 7'h18 == index ? valid1_24 : _GEN_410; // @[icache.scala 79:{31,31}]
  wire  _GEN_412 = 7'h19 == index ? valid1_25 : _GEN_411; // @[icache.scala 79:{31,31}]
  wire  _GEN_413 = 7'h1a == index ? valid1_26 : _GEN_412; // @[icache.scala 79:{31,31}]
  wire  _GEN_414 = 7'h1b == index ? valid1_27 : _GEN_413; // @[icache.scala 79:{31,31}]
  wire  _GEN_415 = 7'h1c == index ? valid1_28 : _GEN_414; // @[icache.scala 79:{31,31}]
  wire  _GEN_416 = 7'h1d == index ? valid1_29 : _GEN_415; // @[icache.scala 79:{31,31}]
  wire  _GEN_417 = 7'h1e == index ? valid1_30 : _GEN_416; // @[icache.scala 79:{31,31}]
  wire  _GEN_418 = 7'h1f == index ? valid1_31 : _GEN_417; // @[icache.scala 79:{31,31}]
  wire  _GEN_419 = 7'h20 == index ? valid1_32 : _GEN_418; // @[icache.scala 79:{31,31}]
  wire  _GEN_420 = 7'h21 == index ? valid1_33 : _GEN_419; // @[icache.scala 79:{31,31}]
  wire  _GEN_421 = 7'h22 == index ? valid1_34 : _GEN_420; // @[icache.scala 79:{31,31}]
  wire  _GEN_422 = 7'h23 == index ? valid1_35 : _GEN_421; // @[icache.scala 79:{31,31}]
  wire  _GEN_423 = 7'h24 == index ? valid1_36 : _GEN_422; // @[icache.scala 79:{31,31}]
  wire  _GEN_424 = 7'h25 == index ? valid1_37 : _GEN_423; // @[icache.scala 79:{31,31}]
  wire  _GEN_425 = 7'h26 == index ? valid1_38 : _GEN_424; // @[icache.scala 79:{31,31}]
  wire  _GEN_426 = 7'h27 == index ? valid1_39 : _GEN_425; // @[icache.scala 79:{31,31}]
  wire  _GEN_427 = 7'h28 == index ? valid1_40 : _GEN_426; // @[icache.scala 79:{31,31}]
  wire  _GEN_428 = 7'h29 == index ? valid1_41 : _GEN_427; // @[icache.scala 79:{31,31}]
  wire  _GEN_429 = 7'h2a == index ? valid1_42 : _GEN_428; // @[icache.scala 79:{31,31}]
  wire  _GEN_430 = 7'h2b == index ? valid1_43 : _GEN_429; // @[icache.scala 79:{31,31}]
  wire  _GEN_431 = 7'h2c == index ? valid1_44 : _GEN_430; // @[icache.scala 79:{31,31}]
  wire  _GEN_432 = 7'h2d == index ? valid1_45 : _GEN_431; // @[icache.scala 79:{31,31}]
  wire  _GEN_433 = 7'h2e == index ? valid1_46 : _GEN_432; // @[icache.scala 79:{31,31}]
  wire  _GEN_434 = 7'h2f == index ? valid1_47 : _GEN_433; // @[icache.scala 79:{31,31}]
  wire  _GEN_435 = 7'h30 == index ? valid1_48 : _GEN_434; // @[icache.scala 79:{31,31}]
  wire  _GEN_436 = 7'h31 == index ? valid1_49 : _GEN_435; // @[icache.scala 79:{31,31}]
  wire  _GEN_437 = 7'h32 == index ? valid1_50 : _GEN_436; // @[icache.scala 79:{31,31}]
  wire  _GEN_438 = 7'h33 == index ? valid1_51 : _GEN_437; // @[icache.scala 79:{31,31}]
  wire  _GEN_439 = 7'h34 == index ? valid1_52 : _GEN_438; // @[icache.scala 79:{31,31}]
  wire  _GEN_440 = 7'h35 == index ? valid1_53 : _GEN_439; // @[icache.scala 79:{31,31}]
  wire  _GEN_441 = 7'h36 == index ? valid1_54 : _GEN_440; // @[icache.scala 79:{31,31}]
  wire  _GEN_442 = 7'h37 == index ? valid1_55 : _GEN_441; // @[icache.scala 79:{31,31}]
  wire  _GEN_443 = 7'h38 == index ? valid1_56 : _GEN_442; // @[icache.scala 79:{31,31}]
  wire  _GEN_444 = 7'h39 == index ? valid1_57 : _GEN_443; // @[icache.scala 79:{31,31}]
  wire  _GEN_445 = 7'h3a == index ? valid1_58 : _GEN_444; // @[icache.scala 79:{31,31}]
  wire  _GEN_446 = 7'h3b == index ? valid1_59 : _GEN_445; // @[icache.scala 79:{31,31}]
  wire  _GEN_447 = 7'h3c == index ? valid1_60 : _GEN_446; // @[icache.scala 79:{31,31}]
  wire  _GEN_448 = 7'h3d == index ? valid1_61 : _GEN_447; // @[icache.scala 79:{31,31}]
  wire  _GEN_449 = 7'h3e == index ? valid1_62 : _GEN_448; // @[icache.scala 79:{31,31}]
  wire  _GEN_450 = 7'h3f == index ? valid1_63 : _GEN_449; // @[icache.scala 79:{31,31}]
  wire  _GEN_451 = 7'h40 == index ? valid1_64 : _GEN_450; // @[icache.scala 79:{31,31}]
  wire  _GEN_452 = 7'h41 == index ? valid1_65 : _GEN_451; // @[icache.scala 79:{31,31}]
  wire  _GEN_453 = 7'h42 == index ? valid1_66 : _GEN_452; // @[icache.scala 79:{31,31}]
  wire  _GEN_454 = 7'h43 == index ? valid1_67 : _GEN_453; // @[icache.scala 79:{31,31}]
  wire  _GEN_455 = 7'h44 == index ? valid1_68 : _GEN_454; // @[icache.scala 79:{31,31}]
  wire  _GEN_456 = 7'h45 == index ? valid1_69 : _GEN_455; // @[icache.scala 79:{31,31}]
  wire  _GEN_457 = 7'h46 == index ? valid1_70 : _GEN_456; // @[icache.scala 79:{31,31}]
  wire  _GEN_458 = 7'h47 == index ? valid1_71 : _GEN_457; // @[icache.scala 79:{31,31}]
  wire  _GEN_459 = 7'h48 == index ? valid1_72 : _GEN_458; // @[icache.scala 79:{31,31}]
  wire  _GEN_460 = 7'h49 == index ? valid1_73 : _GEN_459; // @[icache.scala 79:{31,31}]
  wire  _GEN_461 = 7'h4a == index ? valid1_74 : _GEN_460; // @[icache.scala 79:{31,31}]
  wire  _GEN_462 = 7'h4b == index ? valid1_75 : _GEN_461; // @[icache.scala 79:{31,31}]
  wire  _GEN_463 = 7'h4c == index ? valid1_76 : _GEN_462; // @[icache.scala 79:{31,31}]
  wire  _GEN_464 = 7'h4d == index ? valid1_77 : _GEN_463; // @[icache.scala 79:{31,31}]
  wire  _GEN_465 = 7'h4e == index ? valid1_78 : _GEN_464; // @[icache.scala 79:{31,31}]
  wire  _GEN_466 = 7'h4f == index ? valid1_79 : _GEN_465; // @[icache.scala 79:{31,31}]
  wire  _GEN_467 = 7'h50 == index ? valid1_80 : _GEN_466; // @[icache.scala 79:{31,31}]
  wire  _GEN_468 = 7'h51 == index ? valid1_81 : _GEN_467; // @[icache.scala 79:{31,31}]
  wire  _GEN_469 = 7'h52 == index ? valid1_82 : _GEN_468; // @[icache.scala 79:{31,31}]
  wire  _GEN_470 = 7'h53 == index ? valid1_83 : _GEN_469; // @[icache.scala 79:{31,31}]
  wire  _GEN_471 = 7'h54 == index ? valid1_84 : _GEN_470; // @[icache.scala 79:{31,31}]
  wire  _GEN_472 = 7'h55 == index ? valid1_85 : _GEN_471; // @[icache.scala 79:{31,31}]
  wire  _GEN_473 = 7'h56 == index ? valid1_86 : _GEN_472; // @[icache.scala 79:{31,31}]
  wire  _GEN_474 = 7'h57 == index ? valid1_87 : _GEN_473; // @[icache.scala 79:{31,31}]
  wire  _GEN_475 = 7'h58 == index ? valid1_88 : _GEN_474; // @[icache.scala 79:{31,31}]
  wire  _GEN_476 = 7'h59 == index ? valid1_89 : _GEN_475; // @[icache.scala 79:{31,31}]
  wire  _GEN_477 = 7'h5a == index ? valid1_90 : _GEN_476; // @[icache.scala 79:{31,31}]
  wire  _GEN_478 = 7'h5b == index ? valid1_91 : _GEN_477; // @[icache.scala 79:{31,31}]
  wire  _GEN_479 = 7'h5c == index ? valid1_92 : _GEN_478; // @[icache.scala 79:{31,31}]
  wire  _GEN_480 = 7'h5d == index ? valid1_93 : _GEN_479; // @[icache.scala 79:{31,31}]
  wire  _GEN_481 = 7'h5e == index ? valid1_94 : _GEN_480; // @[icache.scala 79:{31,31}]
  wire  _GEN_482 = 7'h5f == index ? valid1_95 : _GEN_481; // @[icache.scala 79:{31,31}]
  wire  _GEN_483 = 7'h60 == index ? valid1_96 : _GEN_482; // @[icache.scala 79:{31,31}]
  wire  _GEN_484 = 7'h61 == index ? valid1_97 : _GEN_483; // @[icache.scala 79:{31,31}]
  wire  _GEN_485 = 7'h62 == index ? valid1_98 : _GEN_484; // @[icache.scala 79:{31,31}]
  wire  _GEN_486 = 7'h63 == index ? valid1_99 : _GEN_485; // @[icache.scala 79:{31,31}]
  wire  _GEN_487 = 7'h64 == index ? valid1_100 : _GEN_486; // @[icache.scala 79:{31,31}]
  wire  _GEN_488 = 7'h65 == index ? valid1_101 : _GEN_487; // @[icache.scala 79:{31,31}]
  wire  _GEN_489 = 7'h66 == index ? valid1_102 : _GEN_488; // @[icache.scala 79:{31,31}]
  wire  _GEN_490 = 7'h67 == index ? valid1_103 : _GEN_489; // @[icache.scala 79:{31,31}]
  wire  _GEN_491 = 7'h68 == index ? valid1_104 : _GEN_490; // @[icache.scala 79:{31,31}]
  wire  _GEN_492 = 7'h69 == index ? valid1_105 : _GEN_491; // @[icache.scala 79:{31,31}]
  wire  _GEN_493 = 7'h6a == index ? valid1_106 : _GEN_492; // @[icache.scala 79:{31,31}]
  wire  _GEN_494 = 7'h6b == index ? valid1_107 : _GEN_493; // @[icache.scala 79:{31,31}]
  wire  _GEN_495 = 7'h6c == index ? valid1_108 : _GEN_494; // @[icache.scala 79:{31,31}]
  wire  _GEN_496 = 7'h6d == index ? valid1_109 : _GEN_495; // @[icache.scala 79:{31,31}]
  wire  _GEN_497 = 7'h6e == index ? valid1_110 : _GEN_496; // @[icache.scala 79:{31,31}]
  wire  _GEN_498 = 7'h6f == index ? valid1_111 : _GEN_497; // @[icache.scala 79:{31,31}]
  wire  _GEN_499 = 7'h70 == index ? valid1_112 : _GEN_498; // @[icache.scala 79:{31,31}]
  wire  _GEN_500 = 7'h71 == index ? valid1_113 : _GEN_499; // @[icache.scala 79:{31,31}]
  wire  _GEN_501 = 7'h72 == index ? valid1_114 : _GEN_500; // @[icache.scala 79:{31,31}]
  wire  _GEN_502 = 7'h73 == index ? valid1_115 : _GEN_501; // @[icache.scala 79:{31,31}]
  wire  _GEN_503 = 7'h74 == index ? valid1_116 : _GEN_502; // @[icache.scala 79:{31,31}]
  wire  _GEN_504 = 7'h75 == index ? valid1_117 : _GEN_503; // @[icache.scala 79:{31,31}]
  wire  _GEN_505 = 7'h76 == index ? valid1_118 : _GEN_504; // @[icache.scala 79:{31,31}]
  wire  _GEN_506 = 7'h77 == index ? valid1_119 : _GEN_505; // @[icache.scala 79:{31,31}]
  wire  _GEN_507 = 7'h78 == index ? valid1_120 : _GEN_506; // @[icache.scala 79:{31,31}]
  wire  _GEN_508 = 7'h79 == index ? valid1_121 : _GEN_507; // @[icache.scala 79:{31,31}]
  wire  _GEN_509 = 7'h7a == index ? valid1_122 : _GEN_508; // @[icache.scala 79:{31,31}]
  wire  _GEN_510 = 7'h7b == index ? valid1_123 : _GEN_509; // @[icache.scala 79:{31,31}]
  wire  _GEN_511 = 7'h7c == index ? valid1_124 : _GEN_510; // @[icache.scala 79:{31,31}]
  wire  _GEN_512 = 7'h7d == index ? valid1_125 : _GEN_511; // @[icache.scala 79:{31,31}]
  wire  _GEN_513 = 7'h7e == index ? valid1_126 : _GEN_512; // @[icache.scala 79:{31,31}]
  wire  _GEN_514 = 7'h7f == index ? valid1_127 : _GEN_513; // @[icache.scala 79:{31,31}]
  wire  hit_bank_1 = _GEN_514 & _GEN_386 == tag; // @[icache.scala 79:31]
  wire  _GEN_900 = 7'h1 == index2 ? valid1_1 : valid1_0; // @[icache.scala 81:{33,33}]
  wire  _GEN_901 = 7'h2 == index2 ? valid1_2 : _GEN_900; // @[icache.scala 81:{33,33}]
  wire  _GEN_902 = 7'h3 == index2 ? valid1_3 : _GEN_901; // @[icache.scala 81:{33,33}]
  wire  _GEN_903 = 7'h4 == index2 ? valid1_4 : _GEN_902; // @[icache.scala 81:{33,33}]
  wire  _GEN_904 = 7'h5 == index2 ? valid1_5 : _GEN_903; // @[icache.scala 81:{33,33}]
  wire  _GEN_905 = 7'h6 == index2 ? valid1_6 : _GEN_904; // @[icache.scala 81:{33,33}]
  wire  _GEN_906 = 7'h7 == index2 ? valid1_7 : _GEN_905; // @[icache.scala 81:{33,33}]
  wire  _GEN_907 = 7'h8 == index2 ? valid1_8 : _GEN_906; // @[icache.scala 81:{33,33}]
  wire  _GEN_908 = 7'h9 == index2 ? valid1_9 : _GEN_907; // @[icache.scala 81:{33,33}]
  wire  _GEN_909 = 7'ha == index2 ? valid1_10 : _GEN_908; // @[icache.scala 81:{33,33}]
  wire  _GEN_910 = 7'hb == index2 ? valid1_11 : _GEN_909; // @[icache.scala 81:{33,33}]
  wire  _GEN_911 = 7'hc == index2 ? valid1_12 : _GEN_910; // @[icache.scala 81:{33,33}]
  wire  _GEN_912 = 7'hd == index2 ? valid1_13 : _GEN_911; // @[icache.scala 81:{33,33}]
  wire  _GEN_913 = 7'he == index2 ? valid1_14 : _GEN_912; // @[icache.scala 81:{33,33}]
  wire  _GEN_914 = 7'hf == index2 ? valid1_15 : _GEN_913; // @[icache.scala 81:{33,33}]
  wire  _GEN_915 = 7'h10 == index2 ? valid1_16 : _GEN_914; // @[icache.scala 81:{33,33}]
  wire  _GEN_916 = 7'h11 == index2 ? valid1_17 : _GEN_915; // @[icache.scala 81:{33,33}]
  wire  _GEN_917 = 7'h12 == index2 ? valid1_18 : _GEN_916; // @[icache.scala 81:{33,33}]
  wire  _GEN_918 = 7'h13 == index2 ? valid1_19 : _GEN_917; // @[icache.scala 81:{33,33}]
  wire  _GEN_919 = 7'h14 == index2 ? valid1_20 : _GEN_918; // @[icache.scala 81:{33,33}]
  wire  _GEN_920 = 7'h15 == index2 ? valid1_21 : _GEN_919; // @[icache.scala 81:{33,33}]
  wire  _GEN_921 = 7'h16 == index2 ? valid1_22 : _GEN_920; // @[icache.scala 81:{33,33}]
  wire  _GEN_922 = 7'h17 == index2 ? valid1_23 : _GEN_921; // @[icache.scala 81:{33,33}]
  wire  _GEN_923 = 7'h18 == index2 ? valid1_24 : _GEN_922; // @[icache.scala 81:{33,33}]
  wire  _GEN_924 = 7'h19 == index2 ? valid1_25 : _GEN_923; // @[icache.scala 81:{33,33}]
  wire  _GEN_925 = 7'h1a == index2 ? valid1_26 : _GEN_924; // @[icache.scala 81:{33,33}]
  wire  _GEN_926 = 7'h1b == index2 ? valid1_27 : _GEN_925; // @[icache.scala 81:{33,33}]
  wire  _GEN_927 = 7'h1c == index2 ? valid1_28 : _GEN_926; // @[icache.scala 81:{33,33}]
  wire  _GEN_928 = 7'h1d == index2 ? valid1_29 : _GEN_927; // @[icache.scala 81:{33,33}]
  wire  _GEN_929 = 7'h1e == index2 ? valid1_30 : _GEN_928; // @[icache.scala 81:{33,33}]
  wire  _GEN_930 = 7'h1f == index2 ? valid1_31 : _GEN_929; // @[icache.scala 81:{33,33}]
  wire  _GEN_931 = 7'h20 == index2 ? valid1_32 : _GEN_930; // @[icache.scala 81:{33,33}]
  wire  _GEN_932 = 7'h21 == index2 ? valid1_33 : _GEN_931; // @[icache.scala 81:{33,33}]
  wire  _GEN_933 = 7'h22 == index2 ? valid1_34 : _GEN_932; // @[icache.scala 81:{33,33}]
  wire  _GEN_934 = 7'h23 == index2 ? valid1_35 : _GEN_933; // @[icache.scala 81:{33,33}]
  wire  _GEN_935 = 7'h24 == index2 ? valid1_36 : _GEN_934; // @[icache.scala 81:{33,33}]
  wire  _GEN_936 = 7'h25 == index2 ? valid1_37 : _GEN_935; // @[icache.scala 81:{33,33}]
  wire  _GEN_937 = 7'h26 == index2 ? valid1_38 : _GEN_936; // @[icache.scala 81:{33,33}]
  wire  _GEN_938 = 7'h27 == index2 ? valid1_39 : _GEN_937; // @[icache.scala 81:{33,33}]
  wire  _GEN_939 = 7'h28 == index2 ? valid1_40 : _GEN_938; // @[icache.scala 81:{33,33}]
  wire  _GEN_940 = 7'h29 == index2 ? valid1_41 : _GEN_939; // @[icache.scala 81:{33,33}]
  wire  _GEN_941 = 7'h2a == index2 ? valid1_42 : _GEN_940; // @[icache.scala 81:{33,33}]
  wire  _GEN_942 = 7'h2b == index2 ? valid1_43 : _GEN_941; // @[icache.scala 81:{33,33}]
  wire  _GEN_943 = 7'h2c == index2 ? valid1_44 : _GEN_942; // @[icache.scala 81:{33,33}]
  wire  _GEN_944 = 7'h2d == index2 ? valid1_45 : _GEN_943; // @[icache.scala 81:{33,33}]
  wire  _GEN_945 = 7'h2e == index2 ? valid1_46 : _GEN_944; // @[icache.scala 81:{33,33}]
  wire  _GEN_946 = 7'h2f == index2 ? valid1_47 : _GEN_945; // @[icache.scala 81:{33,33}]
  wire  _GEN_947 = 7'h30 == index2 ? valid1_48 : _GEN_946; // @[icache.scala 81:{33,33}]
  wire  _GEN_948 = 7'h31 == index2 ? valid1_49 : _GEN_947; // @[icache.scala 81:{33,33}]
  wire  _GEN_949 = 7'h32 == index2 ? valid1_50 : _GEN_948; // @[icache.scala 81:{33,33}]
  wire  _GEN_950 = 7'h33 == index2 ? valid1_51 : _GEN_949; // @[icache.scala 81:{33,33}]
  wire  _GEN_951 = 7'h34 == index2 ? valid1_52 : _GEN_950; // @[icache.scala 81:{33,33}]
  wire  _GEN_952 = 7'h35 == index2 ? valid1_53 : _GEN_951; // @[icache.scala 81:{33,33}]
  wire  _GEN_953 = 7'h36 == index2 ? valid1_54 : _GEN_952; // @[icache.scala 81:{33,33}]
  wire  _GEN_954 = 7'h37 == index2 ? valid1_55 : _GEN_953; // @[icache.scala 81:{33,33}]
  wire  _GEN_955 = 7'h38 == index2 ? valid1_56 : _GEN_954; // @[icache.scala 81:{33,33}]
  wire  _GEN_956 = 7'h39 == index2 ? valid1_57 : _GEN_955; // @[icache.scala 81:{33,33}]
  wire  _GEN_957 = 7'h3a == index2 ? valid1_58 : _GEN_956; // @[icache.scala 81:{33,33}]
  wire  _GEN_958 = 7'h3b == index2 ? valid1_59 : _GEN_957; // @[icache.scala 81:{33,33}]
  wire  _GEN_959 = 7'h3c == index2 ? valid1_60 : _GEN_958; // @[icache.scala 81:{33,33}]
  wire  _GEN_960 = 7'h3d == index2 ? valid1_61 : _GEN_959; // @[icache.scala 81:{33,33}]
  wire  _GEN_961 = 7'h3e == index2 ? valid1_62 : _GEN_960; // @[icache.scala 81:{33,33}]
  wire  _GEN_962 = 7'h3f == index2 ? valid1_63 : _GEN_961; // @[icache.scala 81:{33,33}]
  wire  _GEN_963 = 7'h40 == index2 ? valid1_64 : _GEN_962; // @[icache.scala 81:{33,33}]
  wire  _GEN_964 = 7'h41 == index2 ? valid1_65 : _GEN_963; // @[icache.scala 81:{33,33}]
  wire  _GEN_965 = 7'h42 == index2 ? valid1_66 : _GEN_964; // @[icache.scala 81:{33,33}]
  wire  _GEN_966 = 7'h43 == index2 ? valid1_67 : _GEN_965; // @[icache.scala 81:{33,33}]
  wire  _GEN_967 = 7'h44 == index2 ? valid1_68 : _GEN_966; // @[icache.scala 81:{33,33}]
  wire  _GEN_968 = 7'h45 == index2 ? valid1_69 : _GEN_967; // @[icache.scala 81:{33,33}]
  wire  _GEN_969 = 7'h46 == index2 ? valid1_70 : _GEN_968; // @[icache.scala 81:{33,33}]
  wire  _GEN_970 = 7'h47 == index2 ? valid1_71 : _GEN_969; // @[icache.scala 81:{33,33}]
  wire  _GEN_971 = 7'h48 == index2 ? valid1_72 : _GEN_970; // @[icache.scala 81:{33,33}]
  wire  _GEN_972 = 7'h49 == index2 ? valid1_73 : _GEN_971; // @[icache.scala 81:{33,33}]
  wire  _GEN_973 = 7'h4a == index2 ? valid1_74 : _GEN_972; // @[icache.scala 81:{33,33}]
  wire  _GEN_974 = 7'h4b == index2 ? valid1_75 : _GEN_973; // @[icache.scala 81:{33,33}]
  wire  _GEN_975 = 7'h4c == index2 ? valid1_76 : _GEN_974; // @[icache.scala 81:{33,33}]
  wire  _GEN_976 = 7'h4d == index2 ? valid1_77 : _GEN_975; // @[icache.scala 81:{33,33}]
  wire  _GEN_977 = 7'h4e == index2 ? valid1_78 : _GEN_976; // @[icache.scala 81:{33,33}]
  wire  _GEN_978 = 7'h4f == index2 ? valid1_79 : _GEN_977; // @[icache.scala 81:{33,33}]
  wire  _GEN_979 = 7'h50 == index2 ? valid1_80 : _GEN_978; // @[icache.scala 81:{33,33}]
  wire  _GEN_980 = 7'h51 == index2 ? valid1_81 : _GEN_979; // @[icache.scala 81:{33,33}]
  wire  _GEN_981 = 7'h52 == index2 ? valid1_82 : _GEN_980; // @[icache.scala 81:{33,33}]
  wire  _GEN_982 = 7'h53 == index2 ? valid1_83 : _GEN_981; // @[icache.scala 81:{33,33}]
  wire  _GEN_983 = 7'h54 == index2 ? valid1_84 : _GEN_982; // @[icache.scala 81:{33,33}]
  wire  _GEN_984 = 7'h55 == index2 ? valid1_85 : _GEN_983; // @[icache.scala 81:{33,33}]
  wire  _GEN_985 = 7'h56 == index2 ? valid1_86 : _GEN_984; // @[icache.scala 81:{33,33}]
  wire  _GEN_986 = 7'h57 == index2 ? valid1_87 : _GEN_985; // @[icache.scala 81:{33,33}]
  wire  _GEN_987 = 7'h58 == index2 ? valid1_88 : _GEN_986; // @[icache.scala 81:{33,33}]
  wire  _GEN_988 = 7'h59 == index2 ? valid1_89 : _GEN_987; // @[icache.scala 81:{33,33}]
  wire  _GEN_989 = 7'h5a == index2 ? valid1_90 : _GEN_988; // @[icache.scala 81:{33,33}]
  wire  _GEN_990 = 7'h5b == index2 ? valid1_91 : _GEN_989; // @[icache.scala 81:{33,33}]
  wire  _GEN_991 = 7'h5c == index2 ? valid1_92 : _GEN_990; // @[icache.scala 81:{33,33}]
  wire  _GEN_992 = 7'h5d == index2 ? valid1_93 : _GEN_991; // @[icache.scala 81:{33,33}]
  wire  _GEN_993 = 7'h5e == index2 ? valid1_94 : _GEN_992; // @[icache.scala 81:{33,33}]
  wire  _GEN_994 = 7'h5f == index2 ? valid1_95 : _GEN_993; // @[icache.scala 81:{33,33}]
  wire  _GEN_995 = 7'h60 == index2 ? valid1_96 : _GEN_994; // @[icache.scala 81:{33,33}]
  wire  _GEN_996 = 7'h61 == index2 ? valid1_97 : _GEN_995; // @[icache.scala 81:{33,33}]
  wire  _GEN_997 = 7'h62 == index2 ? valid1_98 : _GEN_996; // @[icache.scala 81:{33,33}]
  wire  _GEN_998 = 7'h63 == index2 ? valid1_99 : _GEN_997; // @[icache.scala 81:{33,33}]
  wire  _GEN_999 = 7'h64 == index2 ? valid1_100 : _GEN_998; // @[icache.scala 81:{33,33}]
  wire  _GEN_1000 = 7'h65 == index2 ? valid1_101 : _GEN_999; // @[icache.scala 81:{33,33}]
  wire  _GEN_1001 = 7'h66 == index2 ? valid1_102 : _GEN_1000; // @[icache.scala 81:{33,33}]
  wire  _GEN_1002 = 7'h67 == index2 ? valid1_103 : _GEN_1001; // @[icache.scala 81:{33,33}]
  wire  _GEN_1003 = 7'h68 == index2 ? valid1_104 : _GEN_1002; // @[icache.scala 81:{33,33}]
  wire  _GEN_1004 = 7'h69 == index2 ? valid1_105 : _GEN_1003; // @[icache.scala 81:{33,33}]
  wire  _GEN_1005 = 7'h6a == index2 ? valid1_106 : _GEN_1004; // @[icache.scala 81:{33,33}]
  wire  _GEN_1006 = 7'h6b == index2 ? valid1_107 : _GEN_1005; // @[icache.scala 81:{33,33}]
  wire  _GEN_1007 = 7'h6c == index2 ? valid1_108 : _GEN_1006; // @[icache.scala 81:{33,33}]
  wire  _GEN_1008 = 7'h6d == index2 ? valid1_109 : _GEN_1007; // @[icache.scala 81:{33,33}]
  wire  _GEN_1009 = 7'h6e == index2 ? valid1_110 : _GEN_1008; // @[icache.scala 81:{33,33}]
  wire  _GEN_1010 = 7'h6f == index2 ? valid1_111 : _GEN_1009; // @[icache.scala 81:{33,33}]
  wire  _GEN_1011 = 7'h70 == index2 ? valid1_112 : _GEN_1010; // @[icache.scala 81:{33,33}]
  wire  _GEN_1012 = 7'h71 == index2 ? valid1_113 : _GEN_1011; // @[icache.scala 81:{33,33}]
  wire  _GEN_1013 = 7'h72 == index2 ? valid1_114 : _GEN_1012; // @[icache.scala 81:{33,33}]
  wire  _GEN_1014 = 7'h73 == index2 ? valid1_115 : _GEN_1013; // @[icache.scala 81:{33,33}]
  wire  _GEN_1015 = 7'h74 == index2 ? valid1_116 : _GEN_1014; // @[icache.scala 81:{33,33}]
  wire  _GEN_1016 = 7'h75 == index2 ? valid1_117 : _GEN_1015; // @[icache.scala 81:{33,33}]
  wire  _GEN_1017 = 7'h76 == index2 ? valid1_118 : _GEN_1016; // @[icache.scala 81:{33,33}]
  wire  _GEN_1018 = 7'h77 == index2 ? valid1_119 : _GEN_1017; // @[icache.scala 81:{33,33}]
  wire  _GEN_1019 = 7'h78 == index2 ? valid1_120 : _GEN_1018; // @[icache.scala 81:{33,33}]
  wire  _GEN_1020 = 7'h79 == index2 ? valid1_121 : _GEN_1019; // @[icache.scala 81:{33,33}]
  wire  _GEN_1021 = 7'h7a == index2 ? valid1_122 : _GEN_1020; // @[icache.scala 81:{33,33}]
  wire  _GEN_1022 = 7'h7b == index2 ? valid1_123 : _GEN_1021; // @[icache.scala 81:{33,33}]
  wire  _GEN_1023 = 7'h7c == index2 ? valid1_124 : _GEN_1022; // @[icache.scala 81:{33,33}]
  wire  _GEN_1024 = 7'h7d == index2 ? valid1_125 : _GEN_1023; // @[icache.scala 81:{33,33}]
  wire  _GEN_1025 = 7'h7e == index2 ? valid1_126 : _GEN_1024; // @[icache.scala 81:{33,33}]
  wire  _GEN_1026 = 7'h7f == index2 ? valid1_127 : _GEN_1025; // @[icache.scala 81:{33,33}]
  wire  hit = hit_bank_0 | hit_bank_1; // @[icache.scala 83:20]
  wire  _victim_T_1 = ~_GEN_770; // @[icache.scala 85:6]
  wire  _victim_T_5 = _GEN_770 & ~_GEN_1026; // @[icache.scala 86:28]
  wire  victim = _victim_T_1 ? 1'h0 : _victim_T_5; // @[Mux.scala 101:16]
  wire  _next_state_T = state == 2'h0; // @[icache.scala 111:12]
  wire  _next_state_T_1 = state == 2'h1; // @[icache.scala 112:12]
  wire  _next_state_T_3 = state == 2'h1 & ~hit; // @[icache.scala 112:23]
  wire  _next_state_T_5 = _out_reg_T & io_mem_master_readData_valid; // @[icache.scala 113:22]
  wire  _next_state_T_7 = _next_state_T_1 & hit; // @[icache.scala 114:23]
  wire [1:0] _next_state_T_8 = _next_state_T_7 ? 2'h1 : state; // @[Mux.scala 101:16]
  wire [1:0] _next_state_T_9 = _next_state_T_5 ? 2'h1 : _next_state_T_8; // @[Mux.scala 101:16]
  wire [1:0] _next_state_T_10 = _next_state_T_3 ? 2'h2 : _next_state_T_9; // @[Mux.scala 101:16]
  wire [1:0] next_state = _next_state_T ? 2'h1 : _next_state_T_10; // @[Mux.scala 101:16]
  wire  _data_array_0_io_i_wen_T_4 = next_state == 2'h1 & _out_reg_T & ~victim; // @[icache.scala 95:76]
  wire  _data_array_1_io_i_wen_T_4 = next_state == 2'h1 & _out_reg_T & victim; // @[icache.scala 95:76]
  wire  _GEN_2051 = 7'h0 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1027 = 7'h0 == index2 | valid0_0; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2052 = 7'h1 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1028 = 7'h1 == index2 | valid0_1; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2053 = 7'h2 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1029 = 7'h2 == index2 | valid0_2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2054 = 7'h3 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1030 = 7'h3 == index2 | valid0_3; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2055 = 7'h4 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1031 = 7'h4 == index2 | valid0_4; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2056 = 7'h5 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1032 = 7'h5 == index2 | valid0_5; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2057 = 7'h6 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1033 = 7'h6 == index2 | valid0_6; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2058 = 7'h7 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1034 = 7'h7 == index2 | valid0_7; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2059 = 7'h8 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1035 = 7'h8 == index2 | valid0_8; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2060 = 7'h9 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1036 = 7'h9 == index2 | valid0_9; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2061 = 7'ha == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1037 = 7'ha == index2 | valid0_10; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2062 = 7'hb == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1038 = 7'hb == index2 | valid0_11; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2063 = 7'hc == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1039 = 7'hc == index2 | valid0_12; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2064 = 7'hd == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1040 = 7'hd == index2 | valid0_13; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2065 = 7'he == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1041 = 7'he == index2 | valid0_14; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2066 = 7'hf == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1042 = 7'hf == index2 | valid0_15; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2067 = 7'h10 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1043 = 7'h10 == index2 | valid0_16; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2068 = 7'h11 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1044 = 7'h11 == index2 | valid0_17; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2069 = 7'h12 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1045 = 7'h12 == index2 | valid0_18; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2070 = 7'h13 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1046 = 7'h13 == index2 | valid0_19; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2071 = 7'h14 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1047 = 7'h14 == index2 | valid0_20; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2072 = 7'h15 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1048 = 7'h15 == index2 | valid0_21; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2073 = 7'h16 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1049 = 7'h16 == index2 | valid0_22; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2074 = 7'h17 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1050 = 7'h17 == index2 | valid0_23; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2075 = 7'h18 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1051 = 7'h18 == index2 | valid0_24; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2076 = 7'h19 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1052 = 7'h19 == index2 | valid0_25; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2077 = 7'h1a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1053 = 7'h1a == index2 | valid0_26; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2078 = 7'h1b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1054 = 7'h1b == index2 | valid0_27; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2079 = 7'h1c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1055 = 7'h1c == index2 | valid0_28; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2080 = 7'h1d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1056 = 7'h1d == index2 | valid0_29; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2081 = 7'h1e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1057 = 7'h1e == index2 | valid0_30; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2082 = 7'h1f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1058 = 7'h1f == index2 | valid0_31; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2083 = 7'h20 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1059 = 7'h20 == index2 | valid0_32; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2084 = 7'h21 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1060 = 7'h21 == index2 | valid0_33; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2085 = 7'h22 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1061 = 7'h22 == index2 | valid0_34; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2086 = 7'h23 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1062 = 7'h23 == index2 | valid0_35; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2087 = 7'h24 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1063 = 7'h24 == index2 | valid0_36; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2088 = 7'h25 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1064 = 7'h25 == index2 | valid0_37; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2089 = 7'h26 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1065 = 7'h26 == index2 | valid0_38; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2090 = 7'h27 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1066 = 7'h27 == index2 | valid0_39; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2091 = 7'h28 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1067 = 7'h28 == index2 | valid0_40; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2092 = 7'h29 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1068 = 7'h29 == index2 | valid0_41; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2093 = 7'h2a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1069 = 7'h2a == index2 | valid0_42; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2094 = 7'h2b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1070 = 7'h2b == index2 | valid0_43; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2095 = 7'h2c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1071 = 7'h2c == index2 | valid0_44; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2096 = 7'h2d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1072 = 7'h2d == index2 | valid0_45; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2097 = 7'h2e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1073 = 7'h2e == index2 | valid0_46; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2098 = 7'h2f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1074 = 7'h2f == index2 | valid0_47; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2099 = 7'h30 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1075 = 7'h30 == index2 | valid0_48; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2100 = 7'h31 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1076 = 7'h31 == index2 | valid0_49; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2101 = 7'h32 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1077 = 7'h32 == index2 | valid0_50; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2102 = 7'h33 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1078 = 7'h33 == index2 | valid0_51; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2103 = 7'h34 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1079 = 7'h34 == index2 | valid0_52; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2104 = 7'h35 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1080 = 7'h35 == index2 | valid0_53; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2105 = 7'h36 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1081 = 7'h36 == index2 | valid0_54; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2106 = 7'h37 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1082 = 7'h37 == index2 | valid0_55; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2107 = 7'h38 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1083 = 7'h38 == index2 | valid0_56; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2108 = 7'h39 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1084 = 7'h39 == index2 | valid0_57; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2109 = 7'h3a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1085 = 7'h3a == index2 | valid0_58; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2110 = 7'h3b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1086 = 7'h3b == index2 | valid0_59; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2111 = 7'h3c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1087 = 7'h3c == index2 | valid0_60; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2112 = 7'h3d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1088 = 7'h3d == index2 | valid0_61; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2113 = 7'h3e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1089 = 7'h3e == index2 | valid0_62; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2114 = 7'h3f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1090 = 7'h3f == index2 | valid0_63; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2115 = 7'h40 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1091 = 7'h40 == index2 | valid0_64; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2116 = 7'h41 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1092 = 7'h41 == index2 | valid0_65; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2117 = 7'h42 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1093 = 7'h42 == index2 | valid0_66; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2118 = 7'h43 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1094 = 7'h43 == index2 | valid0_67; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2119 = 7'h44 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1095 = 7'h44 == index2 | valid0_68; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2120 = 7'h45 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1096 = 7'h45 == index2 | valid0_69; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2121 = 7'h46 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1097 = 7'h46 == index2 | valid0_70; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2122 = 7'h47 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1098 = 7'h47 == index2 | valid0_71; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2123 = 7'h48 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1099 = 7'h48 == index2 | valid0_72; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2124 = 7'h49 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1100 = 7'h49 == index2 | valid0_73; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2125 = 7'h4a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1101 = 7'h4a == index2 | valid0_74; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2126 = 7'h4b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1102 = 7'h4b == index2 | valid0_75; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2127 = 7'h4c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1103 = 7'h4c == index2 | valid0_76; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2128 = 7'h4d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1104 = 7'h4d == index2 | valid0_77; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2129 = 7'h4e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1105 = 7'h4e == index2 | valid0_78; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2130 = 7'h4f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1106 = 7'h4f == index2 | valid0_79; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2131 = 7'h50 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1107 = 7'h50 == index2 | valid0_80; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2132 = 7'h51 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1108 = 7'h51 == index2 | valid0_81; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2133 = 7'h52 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1109 = 7'h52 == index2 | valid0_82; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2134 = 7'h53 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1110 = 7'h53 == index2 | valid0_83; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2135 = 7'h54 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1111 = 7'h54 == index2 | valid0_84; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2136 = 7'h55 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1112 = 7'h55 == index2 | valid0_85; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2137 = 7'h56 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1113 = 7'h56 == index2 | valid0_86; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2138 = 7'h57 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1114 = 7'h57 == index2 | valid0_87; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2139 = 7'h58 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1115 = 7'h58 == index2 | valid0_88; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2140 = 7'h59 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1116 = 7'h59 == index2 | valid0_89; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2141 = 7'h5a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1117 = 7'h5a == index2 | valid0_90; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2142 = 7'h5b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1118 = 7'h5b == index2 | valid0_91; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2143 = 7'h5c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1119 = 7'h5c == index2 | valid0_92; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2144 = 7'h5d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1120 = 7'h5d == index2 | valid0_93; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2145 = 7'h5e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1121 = 7'h5e == index2 | valid0_94; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2146 = 7'h5f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1122 = 7'h5f == index2 | valid0_95; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2147 = 7'h60 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1123 = 7'h60 == index2 | valid0_96; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2148 = 7'h61 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1124 = 7'h61 == index2 | valid0_97; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2149 = 7'h62 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1125 = 7'h62 == index2 | valid0_98; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2150 = 7'h63 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1126 = 7'h63 == index2 | valid0_99; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2151 = 7'h64 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1127 = 7'h64 == index2 | valid0_100; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2152 = 7'h65 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1128 = 7'h65 == index2 | valid0_101; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2153 = 7'h66 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1129 = 7'h66 == index2 | valid0_102; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2154 = 7'h67 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1130 = 7'h67 == index2 | valid0_103; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2155 = 7'h68 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1131 = 7'h68 == index2 | valid0_104; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2156 = 7'h69 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1132 = 7'h69 == index2 | valid0_105; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2157 = 7'h6a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1133 = 7'h6a == index2 | valid0_106; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2158 = 7'h6b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1134 = 7'h6b == index2 | valid0_107; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2159 = 7'h6c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1135 = 7'h6c == index2 | valid0_108; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2160 = 7'h6d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1136 = 7'h6d == index2 | valid0_109; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2161 = 7'h6e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1137 = 7'h6e == index2 | valid0_110; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2162 = 7'h6f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1138 = 7'h6f == index2 | valid0_111; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2163 = 7'h70 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1139 = 7'h70 == index2 | valid0_112; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2164 = 7'h71 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1140 = 7'h71 == index2 | valid0_113; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2165 = 7'h72 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1141 = 7'h72 == index2 | valid0_114; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2166 = 7'h73 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1142 = 7'h73 == index2 | valid0_115; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2167 = 7'h74 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1143 = 7'h74 == index2 | valid0_116; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2168 = 7'h75 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1144 = 7'h75 == index2 | valid0_117; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2169 = 7'h76 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1145 = 7'h76 == index2 | valid0_118; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2170 = 7'h77 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1146 = 7'h77 == index2 | valid0_119; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2171 = 7'h78 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1147 = 7'h78 == index2 | valid0_120; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2172 = 7'h79 == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1148 = 7'h79 == index2 | valid0_121; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2173 = 7'h7a == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1149 = 7'h7a == index2 | valid0_122; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2174 = 7'h7b == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1150 = 7'h7b == index2 | valid0_123; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2175 = 7'h7c == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1151 = 7'h7c == index2 | valid0_124; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2176 = 7'h7d == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1152 = 7'h7d == index2 | valid0_125; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2177 = 7'h7e == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1153 = 7'h7e == index2 | valid0_126; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_2178 = 7'h7f == index2; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1154 = 7'h7f == index2 | valid0_127; // @[icache.scala 101:{20,20} 30:21]
  wire  _GEN_1539 = _GEN_2051 | valid1_0; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1540 = _GEN_2052 | valid1_1; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1541 = _GEN_2053 | valid1_2; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1542 = _GEN_2054 | valid1_3; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1543 = _GEN_2055 | valid1_4; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1544 = _GEN_2056 | valid1_5; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1545 = _GEN_2057 | valid1_6; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1546 = _GEN_2058 | valid1_7; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1547 = _GEN_2059 | valid1_8; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1548 = _GEN_2060 | valid1_9; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1549 = _GEN_2061 | valid1_10; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1550 = _GEN_2062 | valid1_11; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1551 = _GEN_2063 | valid1_12; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1552 = _GEN_2064 | valid1_13; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1553 = _GEN_2065 | valid1_14; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1554 = _GEN_2066 | valid1_15; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1555 = _GEN_2067 | valid1_16; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1556 = _GEN_2068 | valid1_17; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1557 = _GEN_2069 | valid1_18; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1558 = _GEN_2070 | valid1_19; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1559 = _GEN_2071 | valid1_20; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1560 = _GEN_2072 | valid1_21; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1561 = _GEN_2073 | valid1_22; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1562 = _GEN_2074 | valid1_23; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1563 = _GEN_2075 | valid1_24; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1564 = _GEN_2076 | valid1_25; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1565 = _GEN_2077 | valid1_26; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1566 = _GEN_2078 | valid1_27; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1567 = _GEN_2079 | valid1_28; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1568 = _GEN_2080 | valid1_29; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1569 = _GEN_2081 | valid1_30; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1570 = _GEN_2082 | valid1_31; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1571 = _GEN_2083 | valid1_32; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1572 = _GEN_2084 | valid1_33; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1573 = _GEN_2085 | valid1_34; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1574 = _GEN_2086 | valid1_35; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1575 = _GEN_2087 | valid1_36; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1576 = _GEN_2088 | valid1_37; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1577 = _GEN_2089 | valid1_38; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1578 = _GEN_2090 | valid1_39; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1579 = _GEN_2091 | valid1_40; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1580 = _GEN_2092 | valid1_41; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1581 = _GEN_2093 | valid1_42; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1582 = _GEN_2094 | valid1_43; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1583 = _GEN_2095 | valid1_44; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1584 = _GEN_2096 | valid1_45; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1585 = _GEN_2097 | valid1_46; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1586 = _GEN_2098 | valid1_47; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1587 = _GEN_2099 | valid1_48; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1588 = _GEN_2100 | valid1_49; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1589 = _GEN_2101 | valid1_50; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1590 = _GEN_2102 | valid1_51; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1591 = _GEN_2103 | valid1_52; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1592 = _GEN_2104 | valid1_53; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1593 = _GEN_2105 | valid1_54; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1594 = _GEN_2106 | valid1_55; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1595 = _GEN_2107 | valid1_56; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1596 = _GEN_2108 | valid1_57; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1597 = _GEN_2109 | valid1_58; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1598 = _GEN_2110 | valid1_59; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1599 = _GEN_2111 | valid1_60; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1600 = _GEN_2112 | valid1_61; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1601 = _GEN_2113 | valid1_62; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1602 = _GEN_2114 | valid1_63; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1603 = _GEN_2115 | valid1_64; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1604 = _GEN_2116 | valid1_65; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1605 = _GEN_2117 | valid1_66; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1606 = _GEN_2118 | valid1_67; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1607 = _GEN_2119 | valid1_68; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1608 = _GEN_2120 | valid1_69; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1609 = _GEN_2121 | valid1_70; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1610 = _GEN_2122 | valid1_71; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1611 = _GEN_2123 | valid1_72; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1612 = _GEN_2124 | valid1_73; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1613 = _GEN_2125 | valid1_74; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1614 = _GEN_2126 | valid1_75; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1615 = _GEN_2127 | valid1_76; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1616 = _GEN_2128 | valid1_77; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1617 = _GEN_2129 | valid1_78; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1618 = _GEN_2130 | valid1_79; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1619 = _GEN_2131 | valid1_80; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1620 = _GEN_2132 | valid1_81; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1621 = _GEN_2133 | valid1_82; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1622 = _GEN_2134 | valid1_83; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1623 = _GEN_2135 | valid1_84; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1624 = _GEN_2136 | valid1_85; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1625 = _GEN_2137 | valid1_86; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1626 = _GEN_2138 | valid1_87; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1627 = _GEN_2139 | valid1_88; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1628 = _GEN_2140 | valid1_89; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1629 = _GEN_2141 | valid1_90; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1630 = _GEN_2142 | valid1_91; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1631 = _GEN_2143 | valid1_92; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1632 = _GEN_2144 | valid1_93; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1633 = _GEN_2145 | valid1_94; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1634 = _GEN_2146 | valid1_95; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1635 = _GEN_2147 | valid1_96; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1636 = _GEN_2148 | valid1_97; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1637 = _GEN_2149 | valid1_98; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1638 = _GEN_2150 | valid1_99; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1639 = _GEN_2151 | valid1_100; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1640 = _GEN_2152 | valid1_101; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1641 = _GEN_2153 | valid1_102; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1642 = _GEN_2154 | valid1_103; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1643 = _GEN_2155 | valid1_104; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1644 = _GEN_2156 | valid1_105; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1645 = _GEN_2157 | valid1_106; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1646 = _GEN_2158 | valid1_107; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1647 = _GEN_2159 | valid1_108; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1648 = _GEN_2160 | valid1_109; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1649 = _GEN_2161 | valid1_110; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1650 = _GEN_2162 | valid1_111; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1651 = _GEN_2163 | valid1_112; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1652 = _GEN_2164 | valid1_113; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1653 = _GEN_2165 | valid1_114; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1654 = _GEN_2166 | valid1_115; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1655 = _GEN_2167 | valid1_116; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1656 = _GEN_2168 | valid1_117; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1657 = _GEN_2169 | valid1_118; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1658 = _GEN_2170 | valid1_119; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1659 = _GEN_2171 | valid1_120; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1660 = _GEN_2172 | valid1_121; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1661 = _GEN_2173 | valid1_122; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1662 = _GEN_2174 | valid1_123; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1663 = _GEN_2175 | valid1_124; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1664 = _GEN_2176 | valid1_125; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1665 = _GEN_2177 | valid1_126; // @[icache.scala 105:{20,20} 31:21]
  wire  _GEN_1666 = _GEN_2178 | valid1_127; // @[icache.scala 105:{20,20} 31:21]
  Data_Array data_array_0 ( // @[icache.scala 32:36]
    .clock(data_array_0_clock),
    .reset(data_array_0_reset),
    .io_i_wen(data_array_0_io_i_wen),
    .io_i_wstrb(data_array_0_io_i_wstrb),
    .io_i_addr(data_array_0_io_i_addr),
    .io_i_wdata(data_array_0_io_i_wdata),
    .io_o_rdata(data_array_0_io_o_rdata)
  );
  Data_Array data_array_1 ( // @[icache.scala 32:36]
    .clock(data_array_1_clock),
    .reset(data_array_1_reset),
    .io_i_wen(data_array_1_io_i_wen),
    .io_i_wstrb(data_array_1_io_i_wstrb),
    .io_i_addr(data_array_1_io_i_addr),
    .io_i_wdata(data_array_1_io_i_wdata),
    .io_o_rdata(data_array_1_io_o_rdata)
  );
  assign io_cpu_if_i_data = ~cpu_if2_o_addr[3] ? dout2[63:0] : dout2[127:64]; // @[icache.scala 71:24]
  assign io_cpu_if_i_addr_ready = state != 2'h2; // @[icache.scala 73:34]
  assign io_cpu_if_i_data_valid = state != 2'h2; // @[icache.scala 72:34]
  assign io_mem_master_readAddr_valid = state == 2'h2; // @[icache.scala 118:40]
  assign io_mem_master_readAddr_bits_addr = {cpu_if2_o_addr[63:4],4'h0}; // @[Cat.scala 33:92]
  assign io_mem_master_readAddr_bits_prot = 3'h0; // @[icache.scala 132:34]
  assign io_mem_master_readData_ready = state == 2'h2; // @[icache.scala 120:40]
  assign io_mem_master_writeAddr_valid = 1'h0; // @[icache.scala 125:31]
  assign io_mem_master_writeAddr_bits_addr = 64'h0; // @[icache.scala 131:35]
  assign io_mem_master_writeAddr_bits_prot = 3'h0; // @[icache.scala 129:35]
  assign io_mem_master_writeData_valid = 1'h0; // @[icache.scala 127:31]
  assign io_mem_master_writeData_bits_data = 128'h0; // @[icache.scala 128:34]
  assign io_mem_master_writeData_bits_strb = 16'h0; // @[icache.scala 126:35]
  assign io_mem_master_writeResp_ready = 1'h0; // @[icache.scala 130:31]
  assign data_array_0_clock = clock;
  assign data_array_0_reset = reset;
  assign data_array_0_io_i_wen = next_state == 2'h1 & _out_reg_T & ~victim; // @[icache.scala 95:76]
  assign data_array_0_io_i_wstrb = 16'hffff; // @[icache.scala 96:30]
  assign data_array_0_io_i_addr = _out_reg_T ? index2 : index; // @[icache.scala 97:35]
  assign data_array_0_io_i_wdata = io_mem_master_readData_bits_data; // @[icache.scala 98:30]
  assign data_array_1_clock = clock;
  assign data_array_1_reset = reset;
  assign data_array_1_io_i_wen = next_state == 2'h1 & _out_reg_T & victim; // @[icache.scala 95:76]
  assign data_array_1_io_i_wstrb = 16'hffff; // @[icache.scala 96:30]
  assign data_array_1_io_i_addr = _out_reg_T ? index2 : index; // @[icache.scala 97:35]
  assign data_array_1_io_i_wdata = io_mem_master_readData_bits_data; // @[icache.scala 98:30]
  always @(posedge clock) begin
    if (reset) begin // @[icache.scala 24:22]
      cpu_if1_o_addr <= 64'h0; // @[icache.scala 24:22]
    end else if (!(io_cpu_if_o_stall1)) begin // @[icache.scala 46:25]
      cpu_if1_o_addr <= io_cpu_if_o_addr; // @[icache.scala 49:13]
    end
    if (reset) begin // @[icache.scala 25:22]
      cpu_if2_o_addr <= 64'h0; // @[icache.scala 25:22]
    end else if (~io_cpu_if_o_stall2) begin // @[icache.scala 51:15]
      cpu_if2_o_addr <= cpu_if1_o_addr;
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_0 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h0 == index2) begin // @[icache.scala 102:19]
        tags0_0 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_1 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1 == index2) begin // @[icache.scala 102:19]
        tags0_1 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_2 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2 == index2) begin // @[icache.scala 102:19]
        tags0_2 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_3 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3 == index2) begin // @[icache.scala 102:19]
        tags0_3 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_4 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4 == index2) begin // @[icache.scala 102:19]
        tags0_4 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_5 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5 == index2) begin // @[icache.scala 102:19]
        tags0_5 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_6 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6 == index2) begin // @[icache.scala 102:19]
        tags0_6 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_7 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7 == index2) begin // @[icache.scala 102:19]
        tags0_7 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_8 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h8 == index2) begin // @[icache.scala 102:19]
        tags0_8 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_9 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h9 == index2) begin // @[icache.scala 102:19]
        tags0_9 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_10 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'ha == index2) begin // @[icache.scala 102:19]
        tags0_10 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_11 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'hb == index2) begin // @[icache.scala 102:19]
        tags0_11 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_12 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'hc == index2) begin // @[icache.scala 102:19]
        tags0_12 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_13 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'hd == index2) begin // @[icache.scala 102:19]
        tags0_13 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_14 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'he == index2) begin // @[icache.scala 102:19]
        tags0_14 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_15 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'hf == index2) begin // @[icache.scala 102:19]
        tags0_15 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_16 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h10 == index2) begin // @[icache.scala 102:19]
        tags0_16 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_17 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h11 == index2) begin // @[icache.scala 102:19]
        tags0_17 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_18 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h12 == index2) begin // @[icache.scala 102:19]
        tags0_18 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_19 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h13 == index2) begin // @[icache.scala 102:19]
        tags0_19 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_20 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h14 == index2) begin // @[icache.scala 102:19]
        tags0_20 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_21 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h15 == index2) begin // @[icache.scala 102:19]
        tags0_21 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_22 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h16 == index2) begin // @[icache.scala 102:19]
        tags0_22 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_23 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h17 == index2) begin // @[icache.scala 102:19]
        tags0_23 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_24 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h18 == index2) begin // @[icache.scala 102:19]
        tags0_24 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_25 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h19 == index2) begin // @[icache.scala 102:19]
        tags0_25 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_26 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1a == index2) begin // @[icache.scala 102:19]
        tags0_26 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_27 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1b == index2) begin // @[icache.scala 102:19]
        tags0_27 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_28 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1c == index2) begin // @[icache.scala 102:19]
        tags0_28 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_29 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1d == index2) begin // @[icache.scala 102:19]
        tags0_29 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_30 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1e == index2) begin // @[icache.scala 102:19]
        tags0_30 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_31 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h1f == index2) begin // @[icache.scala 102:19]
        tags0_31 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_32 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h20 == index2) begin // @[icache.scala 102:19]
        tags0_32 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_33 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h21 == index2) begin // @[icache.scala 102:19]
        tags0_33 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_34 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h22 == index2) begin // @[icache.scala 102:19]
        tags0_34 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_35 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h23 == index2) begin // @[icache.scala 102:19]
        tags0_35 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_36 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h24 == index2) begin // @[icache.scala 102:19]
        tags0_36 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_37 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h25 == index2) begin // @[icache.scala 102:19]
        tags0_37 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_38 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h26 == index2) begin // @[icache.scala 102:19]
        tags0_38 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_39 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h27 == index2) begin // @[icache.scala 102:19]
        tags0_39 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_40 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h28 == index2) begin // @[icache.scala 102:19]
        tags0_40 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_41 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h29 == index2) begin // @[icache.scala 102:19]
        tags0_41 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_42 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2a == index2) begin // @[icache.scala 102:19]
        tags0_42 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_43 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2b == index2) begin // @[icache.scala 102:19]
        tags0_43 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_44 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2c == index2) begin // @[icache.scala 102:19]
        tags0_44 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_45 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2d == index2) begin // @[icache.scala 102:19]
        tags0_45 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_46 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2e == index2) begin // @[icache.scala 102:19]
        tags0_46 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_47 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h2f == index2) begin // @[icache.scala 102:19]
        tags0_47 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_48 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h30 == index2) begin // @[icache.scala 102:19]
        tags0_48 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_49 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h31 == index2) begin // @[icache.scala 102:19]
        tags0_49 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_50 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h32 == index2) begin // @[icache.scala 102:19]
        tags0_50 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_51 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h33 == index2) begin // @[icache.scala 102:19]
        tags0_51 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_52 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h34 == index2) begin // @[icache.scala 102:19]
        tags0_52 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_53 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h35 == index2) begin // @[icache.scala 102:19]
        tags0_53 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_54 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h36 == index2) begin // @[icache.scala 102:19]
        tags0_54 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_55 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h37 == index2) begin // @[icache.scala 102:19]
        tags0_55 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_56 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h38 == index2) begin // @[icache.scala 102:19]
        tags0_56 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_57 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h39 == index2) begin // @[icache.scala 102:19]
        tags0_57 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_58 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3a == index2) begin // @[icache.scala 102:19]
        tags0_58 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_59 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3b == index2) begin // @[icache.scala 102:19]
        tags0_59 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_60 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3c == index2) begin // @[icache.scala 102:19]
        tags0_60 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_61 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3d == index2) begin // @[icache.scala 102:19]
        tags0_61 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_62 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3e == index2) begin // @[icache.scala 102:19]
        tags0_62 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_63 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h3f == index2) begin // @[icache.scala 102:19]
        tags0_63 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_64 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h40 == index2) begin // @[icache.scala 102:19]
        tags0_64 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_65 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h41 == index2) begin // @[icache.scala 102:19]
        tags0_65 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_66 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h42 == index2) begin // @[icache.scala 102:19]
        tags0_66 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_67 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h43 == index2) begin // @[icache.scala 102:19]
        tags0_67 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_68 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h44 == index2) begin // @[icache.scala 102:19]
        tags0_68 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_69 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h45 == index2) begin // @[icache.scala 102:19]
        tags0_69 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_70 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h46 == index2) begin // @[icache.scala 102:19]
        tags0_70 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_71 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h47 == index2) begin // @[icache.scala 102:19]
        tags0_71 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_72 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h48 == index2) begin // @[icache.scala 102:19]
        tags0_72 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_73 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h49 == index2) begin // @[icache.scala 102:19]
        tags0_73 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_74 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4a == index2) begin // @[icache.scala 102:19]
        tags0_74 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_75 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4b == index2) begin // @[icache.scala 102:19]
        tags0_75 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_76 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4c == index2) begin // @[icache.scala 102:19]
        tags0_76 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_77 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4d == index2) begin // @[icache.scala 102:19]
        tags0_77 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_78 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4e == index2) begin // @[icache.scala 102:19]
        tags0_78 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_79 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h4f == index2) begin // @[icache.scala 102:19]
        tags0_79 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_80 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h50 == index2) begin // @[icache.scala 102:19]
        tags0_80 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_81 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h51 == index2) begin // @[icache.scala 102:19]
        tags0_81 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_82 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h52 == index2) begin // @[icache.scala 102:19]
        tags0_82 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_83 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h53 == index2) begin // @[icache.scala 102:19]
        tags0_83 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_84 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h54 == index2) begin // @[icache.scala 102:19]
        tags0_84 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_85 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h55 == index2) begin // @[icache.scala 102:19]
        tags0_85 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_86 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h56 == index2) begin // @[icache.scala 102:19]
        tags0_86 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_87 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h57 == index2) begin // @[icache.scala 102:19]
        tags0_87 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_88 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h58 == index2) begin // @[icache.scala 102:19]
        tags0_88 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_89 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h59 == index2) begin // @[icache.scala 102:19]
        tags0_89 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_90 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5a == index2) begin // @[icache.scala 102:19]
        tags0_90 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_91 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5b == index2) begin // @[icache.scala 102:19]
        tags0_91 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_92 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5c == index2) begin // @[icache.scala 102:19]
        tags0_92 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_93 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5d == index2) begin // @[icache.scala 102:19]
        tags0_93 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_94 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5e == index2) begin // @[icache.scala 102:19]
        tags0_94 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_95 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h5f == index2) begin // @[icache.scala 102:19]
        tags0_95 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_96 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h60 == index2) begin // @[icache.scala 102:19]
        tags0_96 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_97 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h61 == index2) begin // @[icache.scala 102:19]
        tags0_97 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_98 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h62 == index2) begin // @[icache.scala 102:19]
        tags0_98 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_99 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h63 == index2) begin // @[icache.scala 102:19]
        tags0_99 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_100 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h64 == index2) begin // @[icache.scala 102:19]
        tags0_100 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_101 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h65 == index2) begin // @[icache.scala 102:19]
        tags0_101 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_102 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h66 == index2) begin // @[icache.scala 102:19]
        tags0_102 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_103 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h67 == index2) begin // @[icache.scala 102:19]
        tags0_103 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_104 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h68 == index2) begin // @[icache.scala 102:19]
        tags0_104 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_105 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h69 == index2) begin // @[icache.scala 102:19]
        tags0_105 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_106 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6a == index2) begin // @[icache.scala 102:19]
        tags0_106 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_107 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6b == index2) begin // @[icache.scala 102:19]
        tags0_107 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_108 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6c == index2) begin // @[icache.scala 102:19]
        tags0_108 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_109 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6d == index2) begin // @[icache.scala 102:19]
        tags0_109 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_110 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6e == index2) begin // @[icache.scala 102:19]
        tags0_110 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_111 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h6f == index2) begin // @[icache.scala 102:19]
        tags0_111 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_112 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h70 == index2) begin // @[icache.scala 102:19]
        tags0_112 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_113 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h71 == index2) begin // @[icache.scala 102:19]
        tags0_113 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_114 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h72 == index2) begin // @[icache.scala 102:19]
        tags0_114 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_115 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h73 == index2) begin // @[icache.scala 102:19]
        tags0_115 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_116 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h74 == index2) begin // @[icache.scala 102:19]
        tags0_116 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_117 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h75 == index2) begin // @[icache.scala 102:19]
        tags0_117 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_118 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h76 == index2) begin // @[icache.scala 102:19]
        tags0_118 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_119 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h77 == index2) begin // @[icache.scala 102:19]
        tags0_119 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_120 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h78 == index2) begin // @[icache.scala 102:19]
        tags0_120 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_121 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h79 == index2) begin // @[icache.scala 102:19]
        tags0_121 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_122 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7a == index2) begin // @[icache.scala 102:19]
        tags0_122 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_123 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7b == index2) begin // @[icache.scala 102:19]
        tags0_123 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_124 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7c == index2) begin // @[icache.scala 102:19]
        tags0_124 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_125 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7d == index2) begin // @[icache.scala 102:19]
        tags0_125 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_126 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7e == index2) begin // @[icache.scala 102:19]
        tags0_126 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 28:20]
      tags0_127 <= 53'h0; // @[icache.scala 28:20]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      if (7'h7f == index2) begin // @[icache.scala 102:19]
        tags0_127 <= cpu_if2_o_addr[63:11]; // @[icache.scala 102:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_0 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h0 == index2) begin // @[icache.scala 106:19]
        tags1_0 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_1 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1 == index2) begin // @[icache.scala 106:19]
        tags1_1 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_2 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2 == index2) begin // @[icache.scala 106:19]
        tags1_2 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_3 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3 == index2) begin // @[icache.scala 106:19]
        tags1_3 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_4 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4 == index2) begin // @[icache.scala 106:19]
        tags1_4 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_5 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5 == index2) begin // @[icache.scala 106:19]
        tags1_5 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_6 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6 == index2) begin // @[icache.scala 106:19]
        tags1_6 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_7 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7 == index2) begin // @[icache.scala 106:19]
        tags1_7 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_8 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h8 == index2) begin // @[icache.scala 106:19]
        tags1_8 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_9 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h9 == index2) begin // @[icache.scala 106:19]
        tags1_9 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_10 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'ha == index2) begin // @[icache.scala 106:19]
        tags1_10 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_11 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'hb == index2) begin // @[icache.scala 106:19]
        tags1_11 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_12 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'hc == index2) begin // @[icache.scala 106:19]
        tags1_12 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_13 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'hd == index2) begin // @[icache.scala 106:19]
        tags1_13 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_14 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'he == index2) begin // @[icache.scala 106:19]
        tags1_14 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_15 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'hf == index2) begin // @[icache.scala 106:19]
        tags1_15 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_16 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h10 == index2) begin // @[icache.scala 106:19]
        tags1_16 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_17 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h11 == index2) begin // @[icache.scala 106:19]
        tags1_17 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_18 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h12 == index2) begin // @[icache.scala 106:19]
        tags1_18 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_19 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h13 == index2) begin // @[icache.scala 106:19]
        tags1_19 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_20 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h14 == index2) begin // @[icache.scala 106:19]
        tags1_20 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_21 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h15 == index2) begin // @[icache.scala 106:19]
        tags1_21 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_22 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h16 == index2) begin // @[icache.scala 106:19]
        tags1_22 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_23 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h17 == index2) begin // @[icache.scala 106:19]
        tags1_23 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_24 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h18 == index2) begin // @[icache.scala 106:19]
        tags1_24 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_25 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h19 == index2) begin // @[icache.scala 106:19]
        tags1_25 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_26 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1a == index2) begin // @[icache.scala 106:19]
        tags1_26 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_27 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1b == index2) begin // @[icache.scala 106:19]
        tags1_27 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_28 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1c == index2) begin // @[icache.scala 106:19]
        tags1_28 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_29 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1d == index2) begin // @[icache.scala 106:19]
        tags1_29 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_30 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1e == index2) begin // @[icache.scala 106:19]
        tags1_30 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_31 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h1f == index2) begin // @[icache.scala 106:19]
        tags1_31 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_32 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h20 == index2) begin // @[icache.scala 106:19]
        tags1_32 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_33 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h21 == index2) begin // @[icache.scala 106:19]
        tags1_33 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_34 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h22 == index2) begin // @[icache.scala 106:19]
        tags1_34 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_35 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h23 == index2) begin // @[icache.scala 106:19]
        tags1_35 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_36 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h24 == index2) begin // @[icache.scala 106:19]
        tags1_36 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_37 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h25 == index2) begin // @[icache.scala 106:19]
        tags1_37 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_38 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h26 == index2) begin // @[icache.scala 106:19]
        tags1_38 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_39 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h27 == index2) begin // @[icache.scala 106:19]
        tags1_39 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_40 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h28 == index2) begin // @[icache.scala 106:19]
        tags1_40 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_41 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h29 == index2) begin // @[icache.scala 106:19]
        tags1_41 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_42 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2a == index2) begin // @[icache.scala 106:19]
        tags1_42 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_43 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2b == index2) begin // @[icache.scala 106:19]
        tags1_43 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_44 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2c == index2) begin // @[icache.scala 106:19]
        tags1_44 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_45 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2d == index2) begin // @[icache.scala 106:19]
        tags1_45 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_46 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2e == index2) begin // @[icache.scala 106:19]
        tags1_46 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_47 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h2f == index2) begin // @[icache.scala 106:19]
        tags1_47 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_48 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h30 == index2) begin // @[icache.scala 106:19]
        tags1_48 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_49 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h31 == index2) begin // @[icache.scala 106:19]
        tags1_49 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_50 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h32 == index2) begin // @[icache.scala 106:19]
        tags1_50 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_51 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h33 == index2) begin // @[icache.scala 106:19]
        tags1_51 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_52 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h34 == index2) begin // @[icache.scala 106:19]
        tags1_52 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_53 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h35 == index2) begin // @[icache.scala 106:19]
        tags1_53 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_54 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h36 == index2) begin // @[icache.scala 106:19]
        tags1_54 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_55 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h37 == index2) begin // @[icache.scala 106:19]
        tags1_55 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_56 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h38 == index2) begin // @[icache.scala 106:19]
        tags1_56 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_57 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h39 == index2) begin // @[icache.scala 106:19]
        tags1_57 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_58 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3a == index2) begin // @[icache.scala 106:19]
        tags1_58 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_59 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3b == index2) begin // @[icache.scala 106:19]
        tags1_59 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_60 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3c == index2) begin // @[icache.scala 106:19]
        tags1_60 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_61 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3d == index2) begin // @[icache.scala 106:19]
        tags1_61 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_62 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3e == index2) begin // @[icache.scala 106:19]
        tags1_62 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_63 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h3f == index2) begin // @[icache.scala 106:19]
        tags1_63 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_64 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h40 == index2) begin // @[icache.scala 106:19]
        tags1_64 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_65 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h41 == index2) begin // @[icache.scala 106:19]
        tags1_65 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_66 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h42 == index2) begin // @[icache.scala 106:19]
        tags1_66 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_67 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h43 == index2) begin // @[icache.scala 106:19]
        tags1_67 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_68 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h44 == index2) begin // @[icache.scala 106:19]
        tags1_68 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_69 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h45 == index2) begin // @[icache.scala 106:19]
        tags1_69 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_70 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h46 == index2) begin // @[icache.scala 106:19]
        tags1_70 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_71 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h47 == index2) begin // @[icache.scala 106:19]
        tags1_71 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_72 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h48 == index2) begin // @[icache.scala 106:19]
        tags1_72 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_73 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h49 == index2) begin // @[icache.scala 106:19]
        tags1_73 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_74 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4a == index2) begin // @[icache.scala 106:19]
        tags1_74 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_75 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4b == index2) begin // @[icache.scala 106:19]
        tags1_75 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_76 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4c == index2) begin // @[icache.scala 106:19]
        tags1_76 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_77 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4d == index2) begin // @[icache.scala 106:19]
        tags1_77 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_78 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4e == index2) begin // @[icache.scala 106:19]
        tags1_78 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_79 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h4f == index2) begin // @[icache.scala 106:19]
        tags1_79 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_80 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h50 == index2) begin // @[icache.scala 106:19]
        tags1_80 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_81 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h51 == index2) begin // @[icache.scala 106:19]
        tags1_81 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_82 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h52 == index2) begin // @[icache.scala 106:19]
        tags1_82 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_83 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h53 == index2) begin // @[icache.scala 106:19]
        tags1_83 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_84 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h54 == index2) begin // @[icache.scala 106:19]
        tags1_84 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_85 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h55 == index2) begin // @[icache.scala 106:19]
        tags1_85 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_86 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h56 == index2) begin // @[icache.scala 106:19]
        tags1_86 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_87 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h57 == index2) begin // @[icache.scala 106:19]
        tags1_87 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_88 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h58 == index2) begin // @[icache.scala 106:19]
        tags1_88 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_89 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h59 == index2) begin // @[icache.scala 106:19]
        tags1_89 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_90 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5a == index2) begin // @[icache.scala 106:19]
        tags1_90 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_91 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5b == index2) begin // @[icache.scala 106:19]
        tags1_91 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_92 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5c == index2) begin // @[icache.scala 106:19]
        tags1_92 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_93 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5d == index2) begin // @[icache.scala 106:19]
        tags1_93 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_94 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5e == index2) begin // @[icache.scala 106:19]
        tags1_94 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_95 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h5f == index2) begin // @[icache.scala 106:19]
        tags1_95 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_96 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h60 == index2) begin // @[icache.scala 106:19]
        tags1_96 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_97 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h61 == index2) begin // @[icache.scala 106:19]
        tags1_97 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_98 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h62 == index2) begin // @[icache.scala 106:19]
        tags1_98 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_99 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h63 == index2) begin // @[icache.scala 106:19]
        tags1_99 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_100 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h64 == index2) begin // @[icache.scala 106:19]
        tags1_100 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_101 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h65 == index2) begin // @[icache.scala 106:19]
        tags1_101 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_102 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h66 == index2) begin // @[icache.scala 106:19]
        tags1_102 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_103 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h67 == index2) begin // @[icache.scala 106:19]
        tags1_103 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_104 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h68 == index2) begin // @[icache.scala 106:19]
        tags1_104 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_105 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h69 == index2) begin // @[icache.scala 106:19]
        tags1_105 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_106 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6a == index2) begin // @[icache.scala 106:19]
        tags1_106 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_107 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6b == index2) begin // @[icache.scala 106:19]
        tags1_107 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_108 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6c == index2) begin // @[icache.scala 106:19]
        tags1_108 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_109 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6d == index2) begin // @[icache.scala 106:19]
        tags1_109 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_110 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6e == index2) begin // @[icache.scala 106:19]
        tags1_110 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_111 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h6f == index2) begin // @[icache.scala 106:19]
        tags1_111 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_112 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h70 == index2) begin // @[icache.scala 106:19]
        tags1_112 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_113 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h71 == index2) begin // @[icache.scala 106:19]
        tags1_113 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_114 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h72 == index2) begin // @[icache.scala 106:19]
        tags1_114 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_115 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h73 == index2) begin // @[icache.scala 106:19]
        tags1_115 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_116 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h74 == index2) begin // @[icache.scala 106:19]
        tags1_116 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_117 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h75 == index2) begin // @[icache.scala 106:19]
        tags1_117 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_118 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h76 == index2) begin // @[icache.scala 106:19]
        tags1_118 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_119 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h77 == index2) begin // @[icache.scala 106:19]
        tags1_119 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_120 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h78 == index2) begin // @[icache.scala 106:19]
        tags1_120 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_121 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h79 == index2) begin // @[icache.scala 106:19]
        tags1_121 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_122 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7a == index2) begin // @[icache.scala 106:19]
        tags1_122 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_123 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7b == index2) begin // @[icache.scala 106:19]
        tags1_123 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_124 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7c == index2) begin // @[icache.scala 106:19]
        tags1_124 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_125 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7d == index2) begin // @[icache.scala 106:19]
        tags1_125 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_126 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7e == index2) begin // @[icache.scala 106:19]
        tags1_126 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 29:20]
      tags1_127 <= 53'h0; // @[icache.scala 29:20]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      if (7'h7f == index2) begin // @[icache.scala 106:19]
        tags1_127 <= cpu_if2_o_addr[63:11]; // @[icache.scala 106:19]
      end
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_0 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_0 <= _GEN_1027;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_1 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_1 <= _GEN_1028;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_2 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_2 <= _GEN_1029;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_3 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_3 <= _GEN_1030;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_4 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_4 <= _GEN_1031;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_5 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_5 <= _GEN_1032;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_6 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_6 <= _GEN_1033;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_7 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_7 <= _GEN_1034;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_8 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_8 <= _GEN_1035;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_9 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_9 <= _GEN_1036;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_10 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_10 <= _GEN_1037;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_11 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_11 <= _GEN_1038;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_12 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_12 <= _GEN_1039;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_13 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_13 <= _GEN_1040;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_14 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_14 <= _GEN_1041;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_15 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_15 <= _GEN_1042;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_16 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_16 <= _GEN_1043;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_17 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_17 <= _GEN_1044;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_18 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_18 <= _GEN_1045;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_19 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_19 <= _GEN_1046;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_20 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_20 <= _GEN_1047;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_21 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_21 <= _GEN_1048;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_22 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_22 <= _GEN_1049;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_23 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_23 <= _GEN_1050;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_24 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_24 <= _GEN_1051;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_25 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_25 <= _GEN_1052;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_26 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_26 <= _GEN_1053;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_27 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_27 <= _GEN_1054;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_28 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_28 <= _GEN_1055;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_29 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_29 <= _GEN_1056;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_30 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_30 <= _GEN_1057;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_31 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_31 <= _GEN_1058;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_32 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_32 <= _GEN_1059;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_33 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_33 <= _GEN_1060;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_34 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_34 <= _GEN_1061;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_35 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_35 <= _GEN_1062;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_36 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_36 <= _GEN_1063;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_37 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_37 <= _GEN_1064;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_38 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_38 <= _GEN_1065;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_39 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_39 <= _GEN_1066;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_40 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_40 <= _GEN_1067;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_41 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_41 <= _GEN_1068;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_42 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_42 <= _GEN_1069;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_43 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_43 <= _GEN_1070;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_44 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_44 <= _GEN_1071;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_45 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_45 <= _GEN_1072;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_46 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_46 <= _GEN_1073;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_47 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_47 <= _GEN_1074;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_48 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_48 <= _GEN_1075;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_49 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_49 <= _GEN_1076;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_50 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_50 <= _GEN_1077;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_51 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_51 <= _GEN_1078;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_52 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_52 <= _GEN_1079;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_53 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_53 <= _GEN_1080;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_54 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_54 <= _GEN_1081;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_55 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_55 <= _GEN_1082;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_56 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_56 <= _GEN_1083;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_57 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_57 <= _GEN_1084;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_58 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_58 <= _GEN_1085;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_59 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_59 <= _GEN_1086;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_60 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_60 <= _GEN_1087;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_61 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_61 <= _GEN_1088;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_62 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_62 <= _GEN_1089;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_63 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_63 <= _GEN_1090;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_64 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_64 <= _GEN_1091;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_65 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_65 <= _GEN_1092;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_66 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_66 <= _GEN_1093;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_67 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_67 <= _GEN_1094;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_68 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_68 <= _GEN_1095;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_69 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_69 <= _GEN_1096;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_70 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_70 <= _GEN_1097;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_71 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_71 <= _GEN_1098;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_72 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_72 <= _GEN_1099;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_73 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_73 <= _GEN_1100;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_74 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_74 <= _GEN_1101;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_75 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_75 <= _GEN_1102;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_76 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_76 <= _GEN_1103;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_77 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_77 <= _GEN_1104;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_78 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_78 <= _GEN_1105;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_79 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_79 <= _GEN_1106;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_80 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_80 <= _GEN_1107;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_81 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_81 <= _GEN_1108;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_82 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_82 <= _GEN_1109;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_83 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_83 <= _GEN_1110;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_84 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_84 <= _GEN_1111;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_85 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_85 <= _GEN_1112;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_86 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_86 <= _GEN_1113;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_87 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_87 <= _GEN_1114;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_88 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_88 <= _GEN_1115;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_89 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_89 <= _GEN_1116;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_90 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_90 <= _GEN_1117;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_91 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_91 <= _GEN_1118;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_92 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_92 <= _GEN_1119;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_93 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_93 <= _GEN_1120;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_94 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_94 <= _GEN_1121;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_95 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_95 <= _GEN_1122;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_96 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_96 <= _GEN_1123;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_97 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_97 <= _GEN_1124;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_98 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_98 <= _GEN_1125;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_99 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_99 <= _GEN_1126;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_100 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_100 <= _GEN_1127;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_101 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_101 <= _GEN_1128;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_102 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_102 <= _GEN_1129;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_103 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_103 <= _GEN_1130;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_104 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_104 <= _GEN_1131;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_105 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_105 <= _GEN_1132;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_106 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_106 <= _GEN_1133;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_107 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_107 <= _GEN_1134;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_108 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_108 <= _GEN_1135;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_109 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_109 <= _GEN_1136;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_110 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_110 <= _GEN_1137;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_111 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_111 <= _GEN_1138;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_112 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_112 <= _GEN_1139;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_113 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_113 <= _GEN_1140;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_114 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_114 <= _GEN_1141;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_115 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_115 <= _GEN_1142;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_116 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_116 <= _GEN_1143;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_117 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_117 <= _GEN_1144;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_118 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_118 <= _GEN_1145;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_119 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_119 <= _GEN_1146;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_120 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_120 <= _GEN_1147;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_121 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_121 <= _GEN_1148;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_122 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_122 <= _GEN_1149;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_123 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_123 <= _GEN_1150;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_124 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_124 <= _GEN_1151;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_125 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_125 <= _GEN_1152;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_126 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_126 <= _GEN_1153;
    end
    if (reset) begin // @[icache.scala 30:21]
      valid0_127 <= 1'h0; // @[icache.scala 30:21]
    end else if (_data_array_0_io_i_wen_T_4) begin // @[icache.scala 100:71]
      valid0_127 <= _GEN_1154;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_0 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_0 <= _GEN_1539;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_1 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_1 <= _GEN_1540;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_2 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_2 <= _GEN_1541;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_3 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_3 <= _GEN_1542;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_4 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_4 <= _GEN_1543;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_5 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_5 <= _GEN_1544;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_6 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_6 <= _GEN_1545;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_7 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_7 <= _GEN_1546;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_8 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_8 <= _GEN_1547;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_9 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_9 <= _GEN_1548;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_10 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_10 <= _GEN_1549;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_11 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_11 <= _GEN_1550;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_12 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_12 <= _GEN_1551;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_13 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_13 <= _GEN_1552;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_14 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_14 <= _GEN_1553;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_15 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_15 <= _GEN_1554;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_16 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_16 <= _GEN_1555;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_17 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_17 <= _GEN_1556;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_18 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_18 <= _GEN_1557;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_19 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_19 <= _GEN_1558;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_20 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_20 <= _GEN_1559;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_21 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_21 <= _GEN_1560;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_22 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_22 <= _GEN_1561;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_23 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_23 <= _GEN_1562;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_24 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_24 <= _GEN_1563;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_25 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_25 <= _GEN_1564;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_26 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_26 <= _GEN_1565;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_27 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_27 <= _GEN_1566;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_28 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_28 <= _GEN_1567;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_29 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_29 <= _GEN_1568;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_30 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_30 <= _GEN_1569;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_31 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_31 <= _GEN_1570;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_32 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_32 <= _GEN_1571;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_33 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_33 <= _GEN_1572;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_34 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_34 <= _GEN_1573;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_35 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_35 <= _GEN_1574;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_36 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_36 <= _GEN_1575;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_37 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_37 <= _GEN_1576;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_38 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_38 <= _GEN_1577;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_39 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_39 <= _GEN_1578;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_40 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_40 <= _GEN_1579;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_41 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_41 <= _GEN_1580;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_42 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_42 <= _GEN_1581;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_43 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_43 <= _GEN_1582;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_44 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_44 <= _GEN_1583;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_45 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_45 <= _GEN_1584;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_46 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_46 <= _GEN_1585;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_47 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_47 <= _GEN_1586;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_48 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_48 <= _GEN_1587;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_49 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_49 <= _GEN_1588;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_50 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_50 <= _GEN_1589;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_51 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_51 <= _GEN_1590;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_52 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_52 <= _GEN_1591;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_53 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_53 <= _GEN_1592;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_54 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_54 <= _GEN_1593;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_55 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_55 <= _GEN_1594;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_56 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_56 <= _GEN_1595;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_57 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_57 <= _GEN_1596;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_58 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_58 <= _GEN_1597;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_59 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_59 <= _GEN_1598;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_60 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_60 <= _GEN_1599;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_61 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_61 <= _GEN_1600;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_62 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_62 <= _GEN_1601;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_63 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_63 <= _GEN_1602;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_64 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_64 <= _GEN_1603;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_65 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_65 <= _GEN_1604;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_66 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_66 <= _GEN_1605;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_67 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_67 <= _GEN_1606;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_68 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_68 <= _GEN_1607;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_69 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_69 <= _GEN_1608;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_70 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_70 <= _GEN_1609;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_71 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_71 <= _GEN_1610;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_72 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_72 <= _GEN_1611;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_73 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_73 <= _GEN_1612;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_74 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_74 <= _GEN_1613;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_75 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_75 <= _GEN_1614;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_76 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_76 <= _GEN_1615;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_77 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_77 <= _GEN_1616;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_78 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_78 <= _GEN_1617;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_79 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_79 <= _GEN_1618;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_80 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_80 <= _GEN_1619;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_81 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_81 <= _GEN_1620;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_82 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_82 <= _GEN_1621;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_83 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_83 <= _GEN_1622;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_84 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_84 <= _GEN_1623;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_85 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_85 <= _GEN_1624;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_86 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_86 <= _GEN_1625;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_87 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_87 <= _GEN_1626;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_88 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_88 <= _GEN_1627;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_89 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_89 <= _GEN_1628;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_90 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_90 <= _GEN_1629;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_91 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_91 <= _GEN_1630;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_92 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_92 <= _GEN_1631;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_93 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_93 <= _GEN_1632;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_94 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_94 <= _GEN_1633;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_95 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_95 <= _GEN_1634;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_96 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_96 <= _GEN_1635;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_97 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_97 <= _GEN_1636;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_98 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_98 <= _GEN_1637;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_99 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_99 <= _GEN_1638;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_100 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_100 <= _GEN_1639;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_101 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_101 <= _GEN_1640;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_102 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_102 <= _GEN_1641;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_103 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_103 <= _GEN_1642;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_104 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_104 <= _GEN_1643;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_105 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_105 <= _GEN_1644;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_106 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_106 <= _GEN_1645;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_107 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_107 <= _GEN_1646;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_108 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_108 <= _GEN_1647;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_109 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_109 <= _GEN_1648;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_110 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_110 <= _GEN_1649;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_111 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_111 <= _GEN_1650;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_112 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_112 <= _GEN_1651;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_113 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_113 <= _GEN_1652;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_114 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_114 <= _GEN_1653;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_115 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_115 <= _GEN_1654;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_116 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_116 <= _GEN_1655;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_117 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_117 <= _GEN_1656;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_118 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_118 <= _GEN_1657;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_119 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_119 <= _GEN_1658;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_120 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_120 <= _GEN_1659;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_121 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_121 <= _GEN_1660;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_122 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_122 <= _GEN_1661;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_123 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_123 <= _GEN_1662;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_124 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_124 <= _GEN_1663;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_125 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_125 <= _GEN_1664;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_126 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_126 <= _GEN_1665;
    end
    if (reset) begin // @[icache.scala 31:21]
      valid1_127 <= 1'h0; // @[icache.scala 31:21]
    end else if (_data_array_1_io_i_wen_T_4) begin // @[icache.scala 104:71]
      valid1_127 <= _GEN_1666;
    end
    if (reset) begin // @[icache.scala 43:20]
      state <= 2'h0; // @[icache.scala 43:20]
    end else if (_next_state_T) begin // @[Mux.scala 101:16]
      state <= 2'h1;
    end else if (_next_state_T_3) begin // @[Mux.scala 101:16]
      state <= 2'h2;
    end else if (_next_state_T_5) begin // @[Mux.scala 101:16]
      state <= 2'h1;
    end else begin
      state <= _next_state_T_8;
    end
    if (reset) begin // @[icache.scala 64:25]
      last_stall <= 1'h0; // @[icache.scala 64:25]
    end else begin
      last_stall <= io_cpu_if_o_stall2; // @[icache.scala 69:12]
    end
    if (reset) begin // @[icache.scala 65:22]
      out_reg <= 128'h0; // @[icache.scala 65:22]
    end else if (state == 2'h2) begin // @[icache.scala 70:15]
      out_reg <= io_mem_master_readData_bits_data;
    end else if (!(last_stall)) begin // @[icache.scala 67:16]
      if (hit_bank2_0) begin // @[icache.scala 66:15]
        out_reg <= data_array_0_io_o_rdata;
      end else begin
        out_reg <= data_array_1_io_o_rdata;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  cpu_if1_o_addr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  cpu_if2_o_addr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  tags0_0 = _RAND_2[52:0];
  _RAND_3 = {2{`RANDOM}};
  tags0_1 = _RAND_3[52:0];
  _RAND_4 = {2{`RANDOM}};
  tags0_2 = _RAND_4[52:0];
  _RAND_5 = {2{`RANDOM}};
  tags0_3 = _RAND_5[52:0];
  _RAND_6 = {2{`RANDOM}};
  tags0_4 = _RAND_6[52:0];
  _RAND_7 = {2{`RANDOM}};
  tags0_5 = _RAND_7[52:0];
  _RAND_8 = {2{`RANDOM}};
  tags0_6 = _RAND_8[52:0];
  _RAND_9 = {2{`RANDOM}};
  tags0_7 = _RAND_9[52:0];
  _RAND_10 = {2{`RANDOM}};
  tags0_8 = _RAND_10[52:0];
  _RAND_11 = {2{`RANDOM}};
  tags0_9 = _RAND_11[52:0];
  _RAND_12 = {2{`RANDOM}};
  tags0_10 = _RAND_12[52:0];
  _RAND_13 = {2{`RANDOM}};
  tags0_11 = _RAND_13[52:0];
  _RAND_14 = {2{`RANDOM}};
  tags0_12 = _RAND_14[52:0];
  _RAND_15 = {2{`RANDOM}};
  tags0_13 = _RAND_15[52:0];
  _RAND_16 = {2{`RANDOM}};
  tags0_14 = _RAND_16[52:0];
  _RAND_17 = {2{`RANDOM}};
  tags0_15 = _RAND_17[52:0];
  _RAND_18 = {2{`RANDOM}};
  tags0_16 = _RAND_18[52:0];
  _RAND_19 = {2{`RANDOM}};
  tags0_17 = _RAND_19[52:0];
  _RAND_20 = {2{`RANDOM}};
  tags0_18 = _RAND_20[52:0];
  _RAND_21 = {2{`RANDOM}};
  tags0_19 = _RAND_21[52:0];
  _RAND_22 = {2{`RANDOM}};
  tags0_20 = _RAND_22[52:0];
  _RAND_23 = {2{`RANDOM}};
  tags0_21 = _RAND_23[52:0];
  _RAND_24 = {2{`RANDOM}};
  tags0_22 = _RAND_24[52:0];
  _RAND_25 = {2{`RANDOM}};
  tags0_23 = _RAND_25[52:0];
  _RAND_26 = {2{`RANDOM}};
  tags0_24 = _RAND_26[52:0];
  _RAND_27 = {2{`RANDOM}};
  tags0_25 = _RAND_27[52:0];
  _RAND_28 = {2{`RANDOM}};
  tags0_26 = _RAND_28[52:0];
  _RAND_29 = {2{`RANDOM}};
  tags0_27 = _RAND_29[52:0];
  _RAND_30 = {2{`RANDOM}};
  tags0_28 = _RAND_30[52:0];
  _RAND_31 = {2{`RANDOM}};
  tags0_29 = _RAND_31[52:0];
  _RAND_32 = {2{`RANDOM}};
  tags0_30 = _RAND_32[52:0];
  _RAND_33 = {2{`RANDOM}};
  tags0_31 = _RAND_33[52:0];
  _RAND_34 = {2{`RANDOM}};
  tags0_32 = _RAND_34[52:0];
  _RAND_35 = {2{`RANDOM}};
  tags0_33 = _RAND_35[52:0];
  _RAND_36 = {2{`RANDOM}};
  tags0_34 = _RAND_36[52:0];
  _RAND_37 = {2{`RANDOM}};
  tags0_35 = _RAND_37[52:0];
  _RAND_38 = {2{`RANDOM}};
  tags0_36 = _RAND_38[52:0];
  _RAND_39 = {2{`RANDOM}};
  tags0_37 = _RAND_39[52:0];
  _RAND_40 = {2{`RANDOM}};
  tags0_38 = _RAND_40[52:0];
  _RAND_41 = {2{`RANDOM}};
  tags0_39 = _RAND_41[52:0];
  _RAND_42 = {2{`RANDOM}};
  tags0_40 = _RAND_42[52:0];
  _RAND_43 = {2{`RANDOM}};
  tags0_41 = _RAND_43[52:0];
  _RAND_44 = {2{`RANDOM}};
  tags0_42 = _RAND_44[52:0];
  _RAND_45 = {2{`RANDOM}};
  tags0_43 = _RAND_45[52:0];
  _RAND_46 = {2{`RANDOM}};
  tags0_44 = _RAND_46[52:0];
  _RAND_47 = {2{`RANDOM}};
  tags0_45 = _RAND_47[52:0];
  _RAND_48 = {2{`RANDOM}};
  tags0_46 = _RAND_48[52:0];
  _RAND_49 = {2{`RANDOM}};
  tags0_47 = _RAND_49[52:0];
  _RAND_50 = {2{`RANDOM}};
  tags0_48 = _RAND_50[52:0];
  _RAND_51 = {2{`RANDOM}};
  tags0_49 = _RAND_51[52:0];
  _RAND_52 = {2{`RANDOM}};
  tags0_50 = _RAND_52[52:0];
  _RAND_53 = {2{`RANDOM}};
  tags0_51 = _RAND_53[52:0];
  _RAND_54 = {2{`RANDOM}};
  tags0_52 = _RAND_54[52:0];
  _RAND_55 = {2{`RANDOM}};
  tags0_53 = _RAND_55[52:0];
  _RAND_56 = {2{`RANDOM}};
  tags0_54 = _RAND_56[52:0];
  _RAND_57 = {2{`RANDOM}};
  tags0_55 = _RAND_57[52:0];
  _RAND_58 = {2{`RANDOM}};
  tags0_56 = _RAND_58[52:0];
  _RAND_59 = {2{`RANDOM}};
  tags0_57 = _RAND_59[52:0];
  _RAND_60 = {2{`RANDOM}};
  tags0_58 = _RAND_60[52:0];
  _RAND_61 = {2{`RANDOM}};
  tags0_59 = _RAND_61[52:0];
  _RAND_62 = {2{`RANDOM}};
  tags0_60 = _RAND_62[52:0];
  _RAND_63 = {2{`RANDOM}};
  tags0_61 = _RAND_63[52:0];
  _RAND_64 = {2{`RANDOM}};
  tags0_62 = _RAND_64[52:0];
  _RAND_65 = {2{`RANDOM}};
  tags0_63 = _RAND_65[52:0];
  _RAND_66 = {2{`RANDOM}};
  tags0_64 = _RAND_66[52:0];
  _RAND_67 = {2{`RANDOM}};
  tags0_65 = _RAND_67[52:0];
  _RAND_68 = {2{`RANDOM}};
  tags0_66 = _RAND_68[52:0];
  _RAND_69 = {2{`RANDOM}};
  tags0_67 = _RAND_69[52:0];
  _RAND_70 = {2{`RANDOM}};
  tags0_68 = _RAND_70[52:0];
  _RAND_71 = {2{`RANDOM}};
  tags0_69 = _RAND_71[52:0];
  _RAND_72 = {2{`RANDOM}};
  tags0_70 = _RAND_72[52:0];
  _RAND_73 = {2{`RANDOM}};
  tags0_71 = _RAND_73[52:0];
  _RAND_74 = {2{`RANDOM}};
  tags0_72 = _RAND_74[52:0];
  _RAND_75 = {2{`RANDOM}};
  tags0_73 = _RAND_75[52:0];
  _RAND_76 = {2{`RANDOM}};
  tags0_74 = _RAND_76[52:0];
  _RAND_77 = {2{`RANDOM}};
  tags0_75 = _RAND_77[52:0];
  _RAND_78 = {2{`RANDOM}};
  tags0_76 = _RAND_78[52:0];
  _RAND_79 = {2{`RANDOM}};
  tags0_77 = _RAND_79[52:0];
  _RAND_80 = {2{`RANDOM}};
  tags0_78 = _RAND_80[52:0];
  _RAND_81 = {2{`RANDOM}};
  tags0_79 = _RAND_81[52:0];
  _RAND_82 = {2{`RANDOM}};
  tags0_80 = _RAND_82[52:0];
  _RAND_83 = {2{`RANDOM}};
  tags0_81 = _RAND_83[52:0];
  _RAND_84 = {2{`RANDOM}};
  tags0_82 = _RAND_84[52:0];
  _RAND_85 = {2{`RANDOM}};
  tags0_83 = _RAND_85[52:0];
  _RAND_86 = {2{`RANDOM}};
  tags0_84 = _RAND_86[52:0];
  _RAND_87 = {2{`RANDOM}};
  tags0_85 = _RAND_87[52:0];
  _RAND_88 = {2{`RANDOM}};
  tags0_86 = _RAND_88[52:0];
  _RAND_89 = {2{`RANDOM}};
  tags0_87 = _RAND_89[52:0];
  _RAND_90 = {2{`RANDOM}};
  tags0_88 = _RAND_90[52:0];
  _RAND_91 = {2{`RANDOM}};
  tags0_89 = _RAND_91[52:0];
  _RAND_92 = {2{`RANDOM}};
  tags0_90 = _RAND_92[52:0];
  _RAND_93 = {2{`RANDOM}};
  tags0_91 = _RAND_93[52:0];
  _RAND_94 = {2{`RANDOM}};
  tags0_92 = _RAND_94[52:0];
  _RAND_95 = {2{`RANDOM}};
  tags0_93 = _RAND_95[52:0];
  _RAND_96 = {2{`RANDOM}};
  tags0_94 = _RAND_96[52:0];
  _RAND_97 = {2{`RANDOM}};
  tags0_95 = _RAND_97[52:0];
  _RAND_98 = {2{`RANDOM}};
  tags0_96 = _RAND_98[52:0];
  _RAND_99 = {2{`RANDOM}};
  tags0_97 = _RAND_99[52:0];
  _RAND_100 = {2{`RANDOM}};
  tags0_98 = _RAND_100[52:0];
  _RAND_101 = {2{`RANDOM}};
  tags0_99 = _RAND_101[52:0];
  _RAND_102 = {2{`RANDOM}};
  tags0_100 = _RAND_102[52:0];
  _RAND_103 = {2{`RANDOM}};
  tags0_101 = _RAND_103[52:0];
  _RAND_104 = {2{`RANDOM}};
  tags0_102 = _RAND_104[52:0];
  _RAND_105 = {2{`RANDOM}};
  tags0_103 = _RAND_105[52:0];
  _RAND_106 = {2{`RANDOM}};
  tags0_104 = _RAND_106[52:0];
  _RAND_107 = {2{`RANDOM}};
  tags0_105 = _RAND_107[52:0];
  _RAND_108 = {2{`RANDOM}};
  tags0_106 = _RAND_108[52:0];
  _RAND_109 = {2{`RANDOM}};
  tags0_107 = _RAND_109[52:0];
  _RAND_110 = {2{`RANDOM}};
  tags0_108 = _RAND_110[52:0];
  _RAND_111 = {2{`RANDOM}};
  tags0_109 = _RAND_111[52:0];
  _RAND_112 = {2{`RANDOM}};
  tags0_110 = _RAND_112[52:0];
  _RAND_113 = {2{`RANDOM}};
  tags0_111 = _RAND_113[52:0];
  _RAND_114 = {2{`RANDOM}};
  tags0_112 = _RAND_114[52:0];
  _RAND_115 = {2{`RANDOM}};
  tags0_113 = _RAND_115[52:0];
  _RAND_116 = {2{`RANDOM}};
  tags0_114 = _RAND_116[52:0];
  _RAND_117 = {2{`RANDOM}};
  tags0_115 = _RAND_117[52:0];
  _RAND_118 = {2{`RANDOM}};
  tags0_116 = _RAND_118[52:0];
  _RAND_119 = {2{`RANDOM}};
  tags0_117 = _RAND_119[52:0];
  _RAND_120 = {2{`RANDOM}};
  tags0_118 = _RAND_120[52:0];
  _RAND_121 = {2{`RANDOM}};
  tags0_119 = _RAND_121[52:0];
  _RAND_122 = {2{`RANDOM}};
  tags0_120 = _RAND_122[52:0];
  _RAND_123 = {2{`RANDOM}};
  tags0_121 = _RAND_123[52:0];
  _RAND_124 = {2{`RANDOM}};
  tags0_122 = _RAND_124[52:0];
  _RAND_125 = {2{`RANDOM}};
  tags0_123 = _RAND_125[52:0];
  _RAND_126 = {2{`RANDOM}};
  tags0_124 = _RAND_126[52:0];
  _RAND_127 = {2{`RANDOM}};
  tags0_125 = _RAND_127[52:0];
  _RAND_128 = {2{`RANDOM}};
  tags0_126 = _RAND_128[52:0];
  _RAND_129 = {2{`RANDOM}};
  tags0_127 = _RAND_129[52:0];
  _RAND_130 = {2{`RANDOM}};
  tags1_0 = _RAND_130[52:0];
  _RAND_131 = {2{`RANDOM}};
  tags1_1 = _RAND_131[52:0];
  _RAND_132 = {2{`RANDOM}};
  tags1_2 = _RAND_132[52:0];
  _RAND_133 = {2{`RANDOM}};
  tags1_3 = _RAND_133[52:0];
  _RAND_134 = {2{`RANDOM}};
  tags1_4 = _RAND_134[52:0];
  _RAND_135 = {2{`RANDOM}};
  tags1_5 = _RAND_135[52:0];
  _RAND_136 = {2{`RANDOM}};
  tags1_6 = _RAND_136[52:0];
  _RAND_137 = {2{`RANDOM}};
  tags1_7 = _RAND_137[52:0];
  _RAND_138 = {2{`RANDOM}};
  tags1_8 = _RAND_138[52:0];
  _RAND_139 = {2{`RANDOM}};
  tags1_9 = _RAND_139[52:0];
  _RAND_140 = {2{`RANDOM}};
  tags1_10 = _RAND_140[52:0];
  _RAND_141 = {2{`RANDOM}};
  tags1_11 = _RAND_141[52:0];
  _RAND_142 = {2{`RANDOM}};
  tags1_12 = _RAND_142[52:0];
  _RAND_143 = {2{`RANDOM}};
  tags1_13 = _RAND_143[52:0];
  _RAND_144 = {2{`RANDOM}};
  tags1_14 = _RAND_144[52:0];
  _RAND_145 = {2{`RANDOM}};
  tags1_15 = _RAND_145[52:0];
  _RAND_146 = {2{`RANDOM}};
  tags1_16 = _RAND_146[52:0];
  _RAND_147 = {2{`RANDOM}};
  tags1_17 = _RAND_147[52:0];
  _RAND_148 = {2{`RANDOM}};
  tags1_18 = _RAND_148[52:0];
  _RAND_149 = {2{`RANDOM}};
  tags1_19 = _RAND_149[52:0];
  _RAND_150 = {2{`RANDOM}};
  tags1_20 = _RAND_150[52:0];
  _RAND_151 = {2{`RANDOM}};
  tags1_21 = _RAND_151[52:0];
  _RAND_152 = {2{`RANDOM}};
  tags1_22 = _RAND_152[52:0];
  _RAND_153 = {2{`RANDOM}};
  tags1_23 = _RAND_153[52:0];
  _RAND_154 = {2{`RANDOM}};
  tags1_24 = _RAND_154[52:0];
  _RAND_155 = {2{`RANDOM}};
  tags1_25 = _RAND_155[52:0];
  _RAND_156 = {2{`RANDOM}};
  tags1_26 = _RAND_156[52:0];
  _RAND_157 = {2{`RANDOM}};
  tags1_27 = _RAND_157[52:0];
  _RAND_158 = {2{`RANDOM}};
  tags1_28 = _RAND_158[52:0];
  _RAND_159 = {2{`RANDOM}};
  tags1_29 = _RAND_159[52:0];
  _RAND_160 = {2{`RANDOM}};
  tags1_30 = _RAND_160[52:0];
  _RAND_161 = {2{`RANDOM}};
  tags1_31 = _RAND_161[52:0];
  _RAND_162 = {2{`RANDOM}};
  tags1_32 = _RAND_162[52:0];
  _RAND_163 = {2{`RANDOM}};
  tags1_33 = _RAND_163[52:0];
  _RAND_164 = {2{`RANDOM}};
  tags1_34 = _RAND_164[52:0];
  _RAND_165 = {2{`RANDOM}};
  tags1_35 = _RAND_165[52:0];
  _RAND_166 = {2{`RANDOM}};
  tags1_36 = _RAND_166[52:0];
  _RAND_167 = {2{`RANDOM}};
  tags1_37 = _RAND_167[52:0];
  _RAND_168 = {2{`RANDOM}};
  tags1_38 = _RAND_168[52:0];
  _RAND_169 = {2{`RANDOM}};
  tags1_39 = _RAND_169[52:0];
  _RAND_170 = {2{`RANDOM}};
  tags1_40 = _RAND_170[52:0];
  _RAND_171 = {2{`RANDOM}};
  tags1_41 = _RAND_171[52:0];
  _RAND_172 = {2{`RANDOM}};
  tags1_42 = _RAND_172[52:0];
  _RAND_173 = {2{`RANDOM}};
  tags1_43 = _RAND_173[52:0];
  _RAND_174 = {2{`RANDOM}};
  tags1_44 = _RAND_174[52:0];
  _RAND_175 = {2{`RANDOM}};
  tags1_45 = _RAND_175[52:0];
  _RAND_176 = {2{`RANDOM}};
  tags1_46 = _RAND_176[52:0];
  _RAND_177 = {2{`RANDOM}};
  tags1_47 = _RAND_177[52:0];
  _RAND_178 = {2{`RANDOM}};
  tags1_48 = _RAND_178[52:0];
  _RAND_179 = {2{`RANDOM}};
  tags1_49 = _RAND_179[52:0];
  _RAND_180 = {2{`RANDOM}};
  tags1_50 = _RAND_180[52:0];
  _RAND_181 = {2{`RANDOM}};
  tags1_51 = _RAND_181[52:0];
  _RAND_182 = {2{`RANDOM}};
  tags1_52 = _RAND_182[52:0];
  _RAND_183 = {2{`RANDOM}};
  tags1_53 = _RAND_183[52:0];
  _RAND_184 = {2{`RANDOM}};
  tags1_54 = _RAND_184[52:0];
  _RAND_185 = {2{`RANDOM}};
  tags1_55 = _RAND_185[52:0];
  _RAND_186 = {2{`RANDOM}};
  tags1_56 = _RAND_186[52:0];
  _RAND_187 = {2{`RANDOM}};
  tags1_57 = _RAND_187[52:0];
  _RAND_188 = {2{`RANDOM}};
  tags1_58 = _RAND_188[52:0];
  _RAND_189 = {2{`RANDOM}};
  tags1_59 = _RAND_189[52:0];
  _RAND_190 = {2{`RANDOM}};
  tags1_60 = _RAND_190[52:0];
  _RAND_191 = {2{`RANDOM}};
  tags1_61 = _RAND_191[52:0];
  _RAND_192 = {2{`RANDOM}};
  tags1_62 = _RAND_192[52:0];
  _RAND_193 = {2{`RANDOM}};
  tags1_63 = _RAND_193[52:0];
  _RAND_194 = {2{`RANDOM}};
  tags1_64 = _RAND_194[52:0];
  _RAND_195 = {2{`RANDOM}};
  tags1_65 = _RAND_195[52:0];
  _RAND_196 = {2{`RANDOM}};
  tags1_66 = _RAND_196[52:0];
  _RAND_197 = {2{`RANDOM}};
  tags1_67 = _RAND_197[52:0];
  _RAND_198 = {2{`RANDOM}};
  tags1_68 = _RAND_198[52:0];
  _RAND_199 = {2{`RANDOM}};
  tags1_69 = _RAND_199[52:0];
  _RAND_200 = {2{`RANDOM}};
  tags1_70 = _RAND_200[52:0];
  _RAND_201 = {2{`RANDOM}};
  tags1_71 = _RAND_201[52:0];
  _RAND_202 = {2{`RANDOM}};
  tags1_72 = _RAND_202[52:0];
  _RAND_203 = {2{`RANDOM}};
  tags1_73 = _RAND_203[52:0];
  _RAND_204 = {2{`RANDOM}};
  tags1_74 = _RAND_204[52:0];
  _RAND_205 = {2{`RANDOM}};
  tags1_75 = _RAND_205[52:0];
  _RAND_206 = {2{`RANDOM}};
  tags1_76 = _RAND_206[52:0];
  _RAND_207 = {2{`RANDOM}};
  tags1_77 = _RAND_207[52:0];
  _RAND_208 = {2{`RANDOM}};
  tags1_78 = _RAND_208[52:0];
  _RAND_209 = {2{`RANDOM}};
  tags1_79 = _RAND_209[52:0];
  _RAND_210 = {2{`RANDOM}};
  tags1_80 = _RAND_210[52:0];
  _RAND_211 = {2{`RANDOM}};
  tags1_81 = _RAND_211[52:0];
  _RAND_212 = {2{`RANDOM}};
  tags1_82 = _RAND_212[52:0];
  _RAND_213 = {2{`RANDOM}};
  tags1_83 = _RAND_213[52:0];
  _RAND_214 = {2{`RANDOM}};
  tags1_84 = _RAND_214[52:0];
  _RAND_215 = {2{`RANDOM}};
  tags1_85 = _RAND_215[52:0];
  _RAND_216 = {2{`RANDOM}};
  tags1_86 = _RAND_216[52:0];
  _RAND_217 = {2{`RANDOM}};
  tags1_87 = _RAND_217[52:0];
  _RAND_218 = {2{`RANDOM}};
  tags1_88 = _RAND_218[52:0];
  _RAND_219 = {2{`RANDOM}};
  tags1_89 = _RAND_219[52:0];
  _RAND_220 = {2{`RANDOM}};
  tags1_90 = _RAND_220[52:0];
  _RAND_221 = {2{`RANDOM}};
  tags1_91 = _RAND_221[52:0];
  _RAND_222 = {2{`RANDOM}};
  tags1_92 = _RAND_222[52:0];
  _RAND_223 = {2{`RANDOM}};
  tags1_93 = _RAND_223[52:0];
  _RAND_224 = {2{`RANDOM}};
  tags1_94 = _RAND_224[52:0];
  _RAND_225 = {2{`RANDOM}};
  tags1_95 = _RAND_225[52:0];
  _RAND_226 = {2{`RANDOM}};
  tags1_96 = _RAND_226[52:0];
  _RAND_227 = {2{`RANDOM}};
  tags1_97 = _RAND_227[52:0];
  _RAND_228 = {2{`RANDOM}};
  tags1_98 = _RAND_228[52:0];
  _RAND_229 = {2{`RANDOM}};
  tags1_99 = _RAND_229[52:0];
  _RAND_230 = {2{`RANDOM}};
  tags1_100 = _RAND_230[52:0];
  _RAND_231 = {2{`RANDOM}};
  tags1_101 = _RAND_231[52:0];
  _RAND_232 = {2{`RANDOM}};
  tags1_102 = _RAND_232[52:0];
  _RAND_233 = {2{`RANDOM}};
  tags1_103 = _RAND_233[52:0];
  _RAND_234 = {2{`RANDOM}};
  tags1_104 = _RAND_234[52:0];
  _RAND_235 = {2{`RANDOM}};
  tags1_105 = _RAND_235[52:0];
  _RAND_236 = {2{`RANDOM}};
  tags1_106 = _RAND_236[52:0];
  _RAND_237 = {2{`RANDOM}};
  tags1_107 = _RAND_237[52:0];
  _RAND_238 = {2{`RANDOM}};
  tags1_108 = _RAND_238[52:0];
  _RAND_239 = {2{`RANDOM}};
  tags1_109 = _RAND_239[52:0];
  _RAND_240 = {2{`RANDOM}};
  tags1_110 = _RAND_240[52:0];
  _RAND_241 = {2{`RANDOM}};
  tags1_111 = _RAND_241[52:0];
  _RAND_242 = {2{`RANDOM}};
  tags1_112 = _RAND_242[52:0];
  _RAND_243 = {2{`RANDOM}};
  tags1_113 = _RAND_243[52:0];
  _RAND_244 = {2{`RANDOM}};
  tags1_114 = _RAND_244[52:0];
  _RAND_245 = {2{`RANDOM}};
  tags1_115 = _RAND_245[52:0];
  _RAND_246 = {2{`RANDOM}};
  tags1_116 = _RAND_246[52:0];
  _RAND_247 = {2{`RANDOM}};
  tags1_117 = _RAND_247[52:0];
  _RAND_248 = {2{`RANDOM}};
  tags1_118 = _RAND_248[52:0];
  _RAND_249 = {2{`RANDOM}};
  tags1_119 = _RAND_249[52:0];
  _RAND_250 = {2{`RANDOM}};
  tags1_120 = _RAND_250[52:0];
  _RAND_251 = {2{`RANDOM}};
  tags1_121 = _RAND_251[52:0];
  _RAND_252 = {2{`RANDOM}};
  tags1_122 = _RAND_252[52:0];
  _RAND_253 = {2{`RANDOM}};
  tags1_123 = _RAND_253[52:0];
  _RAND_254 = {2{`RANDOM}};
  tags1_124 = _RAND_254[52:0];
  _RAND_255 = {2{`RANDOM}};
  tags1_125 = _RAND_255[52:0];
  _RAND_256 = {2{`RANDOM}};
  tags1_126 = _RAND_256[52:0];
  _RAND_257 = {2{`RANDOM}};
  tags1_127 = _RAND_257[52:0];
  _RAND_258 = {1{`RANDOM}};
  valid0_0 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  valid0_1 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  valid0_2 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  valid0_3 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  valid0_4 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  valid0_5 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  valid0_6 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  valid0_7 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  valid0_8 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  valid0_9 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  valid0_10 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  valid0_11 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  valid0_12 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  valid0_13 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  valid0_14 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  valid0_15 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  valid0_16 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  valid0_17 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  valid0_18 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  valid0_19 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  valid0_20 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  valid0_21 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  valid0_22 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  valid0_23 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  valid0_24 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  valid0_25 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  valid0_26 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  valid0_27 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  valid0_28 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  valid0_29 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  valid0_30 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  valid0_31 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  valid0_32 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  valid0_33 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  valid0_34 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  valid0_35 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  valid0_36 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  valid0_37 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  valid0_38 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  valid0_39 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  valid0_40 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  valid0_41 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  valid0_42 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  valid0_43 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  valid0_44 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  valid0_45 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  valid0_46 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  valid0_47 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  valid0_48 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  valid0_49 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  valid0_50 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  valid0_51 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  valid0_52 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  valid0_53 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  valid0_54 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  valid0_55 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  valid0_56 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  valid0_57 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  valid0_58 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  valid0_59 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  valid0_60 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  valid0_61 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  valid0_62 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  valid0_63 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  valid0_64 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  valid0_65 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  valid0_66 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  valid0_67 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  valid0_68 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  valid0_69 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  valid0_70 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  valid0_71 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  valid0_72 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  valid0_73 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  valid0_74 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  valid0_75 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  valid0_76 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  valid0_77 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  valid0_78 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  valid0_79 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  valid0_80 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  valid0_81 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  valid0_82 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  valid0_83 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  valid0_84 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  valid0_85 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  valid0_86 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  valid0_87 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  valid0_88 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  valid0_89 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  valid0_90 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  valid0_91 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  valid0_92 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  valid0_93 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  valid0_94 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  valid0_95 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  valid0_96 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  valid0_97 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  valid0_98 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  valid0_99 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  valid0_100 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  valid0_101 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  valid0_102 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  valid0_103 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  valid0_104 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  valid0_105 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  valid0_106 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  valid0_107 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  valid0_108 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  valid0_109 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  valid0_110 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  valid0_111 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  valid0_112 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  valid0_113 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  valid0_114 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  valid0_115 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  valid0_116 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  valid0_117 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  valid0_118 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  valid0_119 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  valid0_120 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  valid0_121 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  valid0_122 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  valid0_123 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  valid0_124 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  valid0_125 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  valid0_126 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  valid0_127 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  valid1_0 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  valid1_1 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  valid1_2 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  valid1_3 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  valid1_4 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  valid1_5 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  valid1_6 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  valid1_7 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  valid1_8 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  valid1_9 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  valid1_10 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  valid1_11 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  valid1_12 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  valid1_13 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  valid1_14 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  valid1_15 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  valid1_16 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  valid1_17 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  valid1_18 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  valid1_19 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  valid1_20 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  valid1_21 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  valid1_22 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  valid1_23 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  valid1_24 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  valid1_25 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  valid1_26 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  valid1_27 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  valid1_28 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  valid1_29 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  valid1_30 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  valid1_31 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  valid1_32 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  valid1_33 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  valid1_34 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  valid1_35 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  valid1_36 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  valid1_37 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  valid1_38 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  valid1_39 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  valid1_40 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  valid1_41 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  valid1_42 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  valid1_43 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  valid1_44 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  valid1_45 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  valid1_46 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  valid1_47 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  valid1_48 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  valid1_49 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  valid1_50 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  valid1_51 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  valid1_52 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  valid1_53 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  valid1_54 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  valid1_55 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  valid1_56 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  valid1_57 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  valid1_58 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  valid1_59 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  valid1_60 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  valid1_61 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  valid1_62 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  valid1_63 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  valid1_64 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  valid1_65 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  valid1_66 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  valid1_67 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  valid1_68 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  valid1_69 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  valid1_70 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  valid1_71 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  valid1_72 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  valid1_73 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  valid1_74 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  valid1_75 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  valid1_76 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  valid1_77 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  valid1_78 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  valid1_79 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  valid1_80 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  valid1_81 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  valid1_82 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  valid1_83 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  valid1_84 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  valid1_85 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  valid1_86 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  valid1_87 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  valid1_88 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  valid1_89 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  valid1_90 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  valid1_91 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  valid1_92 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  valid1_93 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  valid1_94 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  valid1_95 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  valid1_96 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  valid1_97 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  valid1_98 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  valid1_99 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  valid1_100 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  valid1_101 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  valid1_102 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  valid1_103 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  valid1_104 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  valid1_105 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  valid1_106 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  valid1_107 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  valid1_108 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  valid1_109 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  valid1_110 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  valid1_111 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  valid1_112 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  valid1_113 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  valid1_114 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  valid1_115 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  valid1_116 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  valid1_117 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  valid1_118 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  valid1_119 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  valid1_120 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  valid1_121 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  valid1_122 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  valid1_123 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  valid1_124 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  valid1_125 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  valid1_126 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  valid1_127 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  state = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  last_stall = _RAND_515[0:0];
  _RAND_516 = {4{`RANDOM}};
  out_reg = _RAND_516[127:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

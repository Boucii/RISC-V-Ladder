module Reservation_Station(
  input          clock,
  input          reset,
  input          io_i_dispatch_packs_0_valid,
  input  [31:0]  io_i_dispatch_packs_0_pc,
  input  [31:0]  io_i_dispatch_packs_0_inst,
  input  [6:0]   io_i_dispatch_packs_0_func_code,
  input          io_i_dispatch_packs_0_branch_predict_pack_valid,
  input  [63:0]  io_i_dispatch_packs_0_branch_predict_pack_target,
  input  [3:0]   io_i_dispatch_packs_0_branch_predict_pack_branch_type,
  input          io_i_dispatch_packs_0_branch_predict_pack_select,
  input          io_i_dispatch_packs_0_branch_predict_pack_taken,
  input  [6:0]   io_i_dispatch_packs_0_phy_dst,
  input  [6:0]   io_i_dispatch_packs_0_stale_dst,
  input  [4:0]   io_i_dispatch_packs_0_arch_dst,
  input  [2:0]   io_i_dispatch_packs_0_inst_type,
  input          io_i_dispatch_packs_0_regWen,
  input          io_i_dispatch_packs_0_src1_valid,
  input  [6:0]   io_i_dispatch_packs_0_phy_rs1,
  input  [4:0]   io_i_dispatch_packs_0_arch_rs1,
  input          io_i_dispatch_packs_0_src2_valid,
  input  [6:0]   io_i_dispatch_packs_0_phy_rs2,
  input  [4:0]   io_i_dispatch_packs_0_arch_rs2,
  input  [6:0]   io_i_dispatch_packs_0_rob_idx,
  input  [63:0]  io_i_dispatch_packs_0_imm,
  input  [63:0]  io_i_dispatch_packs_0_src1_value,
  input  [63:0]  io_i_dispatch_packs_0_src2_value,
  input  [2:0]   io_i_dispatch_packs_0_op1_sel,
  input  [2:0]   io_i_dispatch_packs_0_op2_sel,
  input  [4:0]   io_i_dispatch_packs_0_alu_sel,
  input  [3:0]   io_i_dispatch_packs_0_branch_type,
  input  [1:0]   io_i_dispatch_packs_0_mem_type,
  input          io_i_dispatch_packs_1_valid,
  input  [31:0]  io_i_dispatch_packs_1_pc,
  input  [31:0]  io_i_dispatch_packs_1_inst,
  input  [6:0]   io_i_dispatch_packs_1_func_code,
  input          io_i_dispatch_packs_1_branch_predict_pack_valid,
  input  [63:0]  io_i_dispatch_packs_1_branch_predict_pack_target,
  input  [3:0]   io_i_dispatch_packs_1_branch_predict_pack_branch_type,
  input          io_i_dispatch_packs_1_branch_predict_pack_select,
  input          io_i_dispatch_packs_1_branch_predict_pack_taken,
  input  [6:0]   io_i_dispatch_packs_1_phy_dst,
  input  [6:0]   io_i_dispatch_packs_1_stale_dst,
  input  [4:0]   io_i_dispatch_packs_1_arch_dst,
  input  [2:0]   io_i_dispatch_packs_1_inst_type,
  input          io_i_dispatch_packs_1_regWen,
  input          io_i_dispatch_packs_1_src1_valid,
  input  [6:0]   io_i_dispatch_packs_1_phy_rs1,
  input  [4:0]   io_i_dispatch_packs_1_arch_rs1,
  input          io_i_dispatch_packs_1_src2_valid,
  input  [6:0]   io_i_dispatch_packs_1_phy_rs2,
  input  [4:0]   io_i_dispatch_packs_1_arch_rs2,
  input  [6:0]   io_i_dispatch_packs_1_rob_idx,
  input  [63:0]  io_i_dispatch_packs_1_imm,
  input  [63:0]  io_i_dispatch_packs_1_src1_value,
  input  [63:0]  io_i_dispatch_packs_1_src2_value,
  input  [2:0]   io_i_dispatch_packs_1_op1_sel,
  input  [2:0]   io_i_dispatch_packs_1_op2_sel,
  input  [4:0]   io_i_dispatch_packs_1_alu_sel,
  input  [3:0]   io_i_dispatch_packs_1_branch_type,
  input  [1:0]   io_i_dispatch_packs_1_mem_type,
  output         io_o_issue_packs_0_valid,
  output [31:0]  io_o_issue_packs_0_pc,
  output [31:0]  io_o_issue_packs_0_inst,
  output [6:0]   io_o_issue_packs_0_func_code,
  output         io_o_issue_packs_0_branch_predict_pack_valid,
  output [63:0]  io_o_issue_packs_0_branch_predict_pack_target,
  output [3:0]   io_o_issue_packs_0_branch_predict_pack_branch_type,
  output         io_o_issue_packs_0_branch_predict_pack_select,
  output         io_o_issue_packs_0_branch_predict_pack_taken,
  output [6:0]   io_o_issue_packs_0_phy_dst,
  output [6:0]   io_o_issue_packs_0_stale_dst,
  output [4:0]   io_o_issue_packs_0_arch_dst,
  output [2:0]   io_o_issue_packs_0_inst_type,
  output         io_o_issue_packs_0_regWen,
  output         io_o_issue_packs_0_src1_valid,
  output [6:0]   io_o_issue_packs_0_phy_rs1,
  output [4:0]   io_o_issue_packs_0_arch_rs1,
  output         io_o_issue_packs_0_src2_valid,
  output [6:0]   io_o_issue_packs_0_phy_rs2,
  output [4:0]   io_o_issue_packs_0_arch_rs2,
  output [6:0]   io_o_issue_packs_0_rob_idx,
  output [63:0]  io_o_issue_packs_0_imm,
  output [63:0]  io_o_issue_packs_0_src1_value,
  output [63:0]  io_o_issue_packs_0_src2_value,
  output [2:0]   io_o_issue_packs_0_op1_sel,
  output [2:0]   io_o_issue_packs_0_op2_sel,
  output [4:0]   io_o_issue_packs_0_alu_sel,
  output [3:0]   io_o_issue_packs_0_branch_type,
  output [1:0]   io_o_issue_packs_0_mem_type,
  output         io_o_issue_packs_1_valid,
  output [31:0]  io_o_issue_packs_1_pc,
  output [31:0]  io_o_issue_packs_1_inst,
  output [6:0]   io_o_issue_packs_1_func_code,
  output         io_o_issue_packs_1_branch_predict_pack_valid,
  output [63:0]  io_o_issue_packs_1_branch_predict_pack_target,
  output [3:0]   io_o_issue_packs_1_branch_predict_pack_branch_type,
  output         io_o_issue_packs_1_branch_predict_pack_select,
  output         io_o_issue_packs_1_branch_predict_pack_taken,
  output [6:0]   io_o_issue_packs_1_phy_dst,
  output [6:0]   io_o_issue_packs_1_stale_dst,
  output [4:0]   io_o_issue_packs_1_arch_dst,
  output [2:0]   io_o_issue_packs_1_inst_type,
  output         io_o_issue_packs_1_regWen,
  output         io_o_issue_packs_1_src1_valid,
  output [6:0]   io_o_issue_packs_1_phy_rs1,
  output [4:0]   io_o_issue_packs_1_arch_rs1,
  output         io_o_issue_packs_1_src2_valid,
  output [6:0]   io_o_issue_packs_1_phy_rs2,
  output [4:0]   io_o_issue_packs_1_arch_rs2,
  output [6:0]   io_o_issue_packs_1_rob_idx,
  output [63:0]  io_o_issue_packs_1_imm,
  output [63:0]  io_o_issue_packs_1_src1_value,
  output [63:0]  io_o_issue_packs_1_src2_value,
  output [2:0]   io_o_issue_packs_1_op1_sel,
  output [2:0]   io_o_issue_packs_1_op2_sel,
  output [4:0]   io_o_issue_packs_1_alu_sel,
  output [3:0]   io_o_issue_packs_1_branch_type,
  output [1:0]   io_o_issue_packs_1_mem_type,
  input  [127:0] io_i_wakeup_port,
  input          io_i_ex_res_packs_0_valid,
  input  [6:0]   io_i_ex_res_packs_0_uop_func_code,
  input  [6:0]   io_i_ex_res_packs_0_uop_phy_dst,
  input  [63:0]  io_i_ex_res_packs_0_uop_dst_value,
  input          io_i_ex_res_packs_1_valid,
  input  [6:0]   io_i_ex_res_packs_1_uop_func_code,
  input  [6:0]   io_i_ex_res_packs_1_uop_phy_dst,
  input  [63:0]  io_i_ex_res_packs_1_uop_dst_value,
  input          io_i_branch_resolve_pack_valid,
  input          io_i_branch_resolve_pack_mispred,
  input  [6:0]   io_i_branch_resolve_pack_rob_idx,
  output         io_o_full,
  input          io_i_exception,
  input          io_i_rollback_valid,
  input  [1:0]   io_i_available_funcs_0,
  input  [1:0]   io_i_available_funcs_1,
  input  [1:0]   io_i_available_funcs_2,
  input  [1:0]   io_i_available_funcs_3,
  input  [1:0]   io_i_available_funcs_4,
  input  [1:0]   io_i_available_funcs_5,
  input  [6:0]   io_i_ROB_first_entry
);
  wire  reservation_station_0_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_0_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_0_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_0_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_0_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_0_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_0_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_0_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_0_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_0_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_0_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_1_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_1_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_1_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_1_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_1_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_1_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_1_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_1_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_1_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_1_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_2_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_2_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_2_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_2_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_2_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_2_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_2_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_2_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_2_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_2_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_3_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_3_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_3_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_3_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_3_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_3_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_3_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_3_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_3_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_3_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_4_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_4_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_4_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_4_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_4_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_4_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_4_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_4_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_4_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_4_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_5_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_5_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_5_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_5_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_5_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_5_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_5_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_5_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_5_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_5_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_6_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_6_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_6_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_6_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_6_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_6_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_6_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_6_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_6_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_6_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_7_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_7_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_7_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_7_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_7_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_7_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_7_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_7_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_7_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_7_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_8_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_8_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_8_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_8_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_8_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_8_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_8_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_8_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_8_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_8_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_9_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_9_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_9_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_9_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_9_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_9_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_9_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_9_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_9_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_9_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_10_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_10_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_10_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_10_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_10_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_10_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_10_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_10_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_10_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_10_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_11_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_11_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_11_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_11_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_11_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_11_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_11_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_11_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_11_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_11_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_12_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_12_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_12_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_12_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_12_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_12_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_12_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_12_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_12_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_12_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_13_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_13_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_13_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_13_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_13_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_13_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_13_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_13_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_13_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_13_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_14_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_14_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_14_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_14_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_14_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_14_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_14_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_14_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_14_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_14_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_15_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_15_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_15_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_15_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_15_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_15_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_15_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_15_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_15_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_15_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_16_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_16_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_16_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_16_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_16_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_16_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_16_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_16_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_16_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_16_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_17_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_17_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_17_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_17_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_17_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_17_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_17_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_17_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_17_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_17_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_18_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_18_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_18_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_18_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_18_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_18_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_18_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_18_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_18_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_18_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_19_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_19_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_19_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_19_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_19_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_19_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_19_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_19_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_19_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_19_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_20_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_20_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_20_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_20_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_20_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_20_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_20_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_20_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_20_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_20_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_21_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_21_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_21_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_21_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_21_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_21_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_21_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_21_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_21_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_21_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_22_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_22_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_22_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_22_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_22_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_22_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_22_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_22_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_22_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_22_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_23_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_23_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_23_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_23_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_23_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_23_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_23_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_23_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_23_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_23_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_24_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_24_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_24_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_24_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_24_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_24_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_24_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_24_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_24_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_24_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_25_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_25_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_25_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_25_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_25_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_25_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_25_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_25_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_25_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_25_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_26_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_26_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_26_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_26_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_26_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_26_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_26_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_26_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_26_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_26_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_27_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_27_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_27_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_27_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_27_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_27_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_27_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_27_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_27_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_27_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_28_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_28_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_28_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_28_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_28_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_28_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_28_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_28_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_28_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_28_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_29_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_29_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_29_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_29_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_29_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_29_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_29_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_29_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_29_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_29_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_30_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_30_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_30_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_30_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_30_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_30_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_30_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_30_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_30_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_30_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_31_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_31_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_31_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_31_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_31_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_31_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_31_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_31_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_31_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_31_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_32_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_32_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_32_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_32_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_32_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_32_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_32_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_32_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_32_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_32_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_33_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_33_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_33_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_33_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_33_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_33_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_33_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_33_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_33_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_33_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_34_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_34_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_34_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_34_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_34_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_34_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_34_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_34_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_34_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_34_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_35_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_35_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_35_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_35_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_35_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_35_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_35_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_35_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_35_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_35_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_36_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_36_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_36_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_36_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_36_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_36_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_36_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_36_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_36_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_36_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_37_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_37_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_37_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_37_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_37_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_37_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_37_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_37_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_37_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_37_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_38_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_38_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_38_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_38_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_38_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_38_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_38_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_38_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_38_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_38_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_39_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_39_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_39_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_39_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_39_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_39_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_39_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_39_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_39_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_39_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_40_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_40_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_40_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_40_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_40_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_40_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_40_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_40_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_40_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_40_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_41_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_41_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_41_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_41_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_41_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_41_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_41_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_41_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_41_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_41_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_42_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_42_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_42_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_42_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_42_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_42_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_42_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_42_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_42_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_42_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_43_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_43_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_43_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_43_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_43_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_43_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_43_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_43_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_43_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_43_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_44_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_44_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_44_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_44_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_44_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_44_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_44_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_44_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_44_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_44_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_45_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_45_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_45_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_45_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_45_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_45_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_45_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_45_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_45_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_45_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_46_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_46_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_46_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_46_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_46_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_46_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_46_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_46_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_46_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_46_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_47_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_47_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_47_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_47_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_47_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_47_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_47_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_47_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_47_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_47_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_48_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_48_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_48_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_48_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_48_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_48_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_48_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_48_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_48_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_48_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_49_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_49_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_49_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_49_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_49_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_49_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_49_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_49_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_49_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_49_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_50_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_50_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_50_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_50_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_50_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_50_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_50_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_50_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_50_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_50_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_51_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_51_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_51_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_51_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_51_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_51_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_51_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_51_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_51_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_51_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_52_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_52_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_52_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_52_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_52_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_52_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_52_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_52_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_52_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_52_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_53_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_53_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_53_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_53_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_53_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_53_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_53_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_53_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_53_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_53_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_54_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_54_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_54_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_54_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_54_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_54_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_54_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_54_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_54_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_54_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_55_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_55_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_55_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_55_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_55_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_55_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_55_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_55_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_55_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_55_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_56_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_56_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_56_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_56_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_56_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_56_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_56_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_56_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_56_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_56_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_57_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_57_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_57_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_57_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_57_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_57_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_57_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_57_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_57_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_57_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_58_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_58_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_58_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_58_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_58_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_58_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_58_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_58_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_58_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_58_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_59_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_59_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_59_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_59_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_59_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_59_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_59_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_59_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_59_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_59_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_60_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_60_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_60_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_60_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_60_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_60_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_60_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_60_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_60_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_60_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_61_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_61_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_61_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_61_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_61_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_61_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_61_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_61_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_61_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_61_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_62_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_62_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_62_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_62_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_62_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_62_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_62_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_62_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_62_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_62_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_clock; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_reset; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_ready_to_issue; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_issue_granted; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_branch_resolve_pack_valid; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_exception; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_write_slot; // @[reservation_station.scala 38:51]
  wire [127:0] reservation_station_63_io_i_wakeup_port; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_valid; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_i_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_i_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_i_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_i_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_i_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_i_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_i_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_i_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_i_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_63_io_i_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_o_uop_pc; // @[reservation_station.scala 38:51]
  wire [31:0] reservation_station_63_io_o_uop_inst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_func_code; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_branch_predict_pack_valid; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_branch_predict_pack_target; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_o_uop_branch_predict_pack_branch_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_branch_predict_pack_select; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_branch_predict_pack_taken; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_phy_dst; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_stale_dst; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_arch_dst; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_o_uop_inst_type; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_regWen; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_src1_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_phy_rs1; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_arch_rs1; // @[reservation_station.scala 38:51]
  wire  reservation_station_63_io_o_uop_src2_valid; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_phy_rs2; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_arch_rs2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_o_uop_rob_idx; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_imm; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_src1_value; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_o_uop_src2_value; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_o_uop_op1_sel; // @[reservation_station.scala 38:51]
  wire [2:0] reservation_station_63_io_o_uop_op2_sel; // @[reservation_station.scala 38:51]
  wire [4:0] reservation_station_63_io_o_uop_alu_sel; // @[reservation_station.scala 38:51]
  wire [3:0] reservation_station_63_io_o_uop_branch_type; // @[reservation_station.scala 38:51]
  wire [1:0] reservation_station_63_io_o_uop_mem_type; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_exe_dst1; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_exe_dst2; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_exe_value1; // @[reservation_station.scala 38:51]
  wire [63:0] reservation_station_63_io_i_exe_value2; // @[reservation_station.scala 38:51]
  wire [6:0] reservation_station_63_io_i_ROB_first_entry; // @[reservation_station.scala 38:51]
  wire  temp_1 = reservation_station_1_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_0 = reservation_station_0_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_3 = reservation_station_3_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_2 = reservation_station_2_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_5 = reservation_station_5_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_4 = reservation_station_4_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_7 = reservation_station_7_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_6 = reservation_station_6_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_lo_lo_lo = {temp_7,temp_6,temp_5,temp_4,temp_3,temp_2,temp_1,temp_0}; // @[reservation_station.scala 48:46]
  wire  temp_9 = reservation_station_9_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_8 = reservation_station_8_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_11 = reservation_station_11_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_10 = reservation_station_10_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_13 = reservation_station_13_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_12 = reservation_station_12_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_15 = reservation_station_15_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_14 = reservation_station_14_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [15:0] reservation_station_valid_lo_lo = {temp_15,temp_14,temp_13,temp_12,temp_11,temp_10,temp_9,temp_8,
    reservation_station_valid_lo_lo_lo}; // @[reservation_station.scala 48:46]
  wire  temp_17 = reservation_station_17_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_16 = reservation_station_16_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_19 = reservation_station_19_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_18 = reservation_station_18_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_21 = reservation_station_21_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_20 = reservation_station_20_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_23 = reservation_station_23_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_22 = reservation_station_22_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_lo_hi_lo = {temp_23,temp_22,temp_21,temp_20,temp_19,temp_18,temp_17,temp_16}; // @[reservation_station.scala 48:46]
  wire  temp_25 = reservation_station_25_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_24 = reservation_station_24_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_27 = reservation_station_27_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_26 = reservation_station_26_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_29 = reservation_station_29_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_28 = reservation_station_28_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_31 = reservation_station_31_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_30 = reservation_station_30_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [31:0] reservation_station_valid_lo = {temp_31,temp_30,temp_29,temp_28,temp_27,temp_26,temp_25,temp_24,
    reservation_station_valid_lo_hi_lo,reservation_station_valid_lo_lo}; // @[reservation_station.scala 48:46]
  wire  temp_33 = reservation_station_33_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_32 = reservation_station_32_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_35 = reservation_station_35_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_34 = reservation_station_34_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_37 = reservation_station_37_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_36 = reservation_station_36_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_39 = reservation_station_39_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_38 = reservation_station_38_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_hi_lo_lo = {temp_39,temp_38,temp_37,temp_36,temp_35,temp_34,temp_33,temp_32}; // @[reservation_station.scala 48:46]
  wire  temp_41 = reservation_station_41_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_40 = reservation_station_40_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_43 = reservation_station_43_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_42 = reservation_station_42_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_45 = reservation_station_45_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_44 = reservation_station_44_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_47 = reservation_station_47_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_46 = reservation_station_46_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [15:0] reservation_station_valid_hi_lo = {temp_47,temp_46,temp_45,temp_44,temp_43,temp_42,temp_41,temp_40,
    reservation_station_valid_hi_lo_lo}; // @[reservation_station.scala 48:46]
  wire  temp_49 = reservation_station_49_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_48 = reservation_station_48_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_51 = reservation_station_51_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_50 = reservation_station_50_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_53 = reservation_station_53_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_52 = reservation_station_52_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_55 = reservation_station_55_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_54 = reservation_station_54_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [7:0] reservation_station_valid_hi_hi_lo = {temp_55,temp_54,temp_53,temp_52,temp_51,temp_50,temp_49,temp_48}; // @[reservation_station.scala 48:46]
  wire  temp_57 = reservation_station_57_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_56 = reservation_station_56_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_59 = reservation_station_59_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_58 = reservation_station_58_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_61 = reservation_station_61_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_60 = reservation_station_60_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_63 = reservation_station_63_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire  temp_62 = reservation_station_62_io_o_valid; // @[reservation_station.scala 41:21 43:16]
  wire [31:0] reservation_station_valid_hi = {temp_63,temp_62,temp_61,temp_60,temp_59,temp_58,temp_57,temp_56,
    reservation_station_valid_hi_hi_lo,reservation_station_valid_hi_lo}; // @[reservation_station.scala 48:46]
  wire [63:0] reservation_station_valid = {reservation_station_valid_hi,reservation_station_valid_lo}; // @[reservation_station.scala 48:46]
  wire [63:0] _write_idx1_T = ~reservation_station_valid; // @[reservation_station.scala 49:34]
  wire [5:0] _write_idx1_T_65 = _write_idx1_T[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_66 = _write_idx1_T[61] ? 6'h3d : _write_idx1_T_65; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_67 = _write_idx1_T[60] ? 6'h3c : _write_idx1_T_66; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_68 = _write_idx1_T[59] ? 6'h3b : _write_idx1_T_67; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_69 = _write_idx1_T[58] ? 6'h3a : _write_idx1_T_68; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_70 = _write_idx1_T[57] ? 6'h39 : _write_idx1_T_69; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_71 = _write_idx1_T[56] ? 6'h38 : _write_idx1_T_70; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_72 = _write_idx1_T[55] ? 6'h37 : _write_idx1_T_71; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_73 = _write_idx1_T[54] ? 6'h36 : _write_idx1_T_72; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_74 = _write_idx1_T[53] ? 6'h35 : _write_idx1_T_73; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_75 = _write_idx1_T[52] ? 6'h34 : _write_idx1_T_74; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_76 = _write_idx1_T[51] ? 6'h33 : _write_idx1_T_75; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_77 = _write_idx1_T[50] ? 6'h32 : _write_idx1_T_76; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_78 = _write_idx1_T[49] ? 6'h31 : _write_idx1_T_77; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_79 = _write_idx1_T[48] ? 6'h30 : _write_idx1_T_78; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_80 = _write_idx1_T[47] ? 6'h2f : _write_idx1_T_79; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_81 = _write_idx1_T[46] ? 6'h2e : _write_idx1_T_80; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_82 = _write_idx1_T[45] ? 6'h2d : _write_idx1_T_81; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_83 = _write_idx1_T[44] ? 6'h2c : _write_idx1_T_82; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_84 = _write_idx1_T[43] ? 6'h2b : _write_idx1_T_83; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_85 = _write_idx1_T[42] ? 6'h2a : _write_idx1_T_84; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_86 = _write_idx1_T[41] ? 6'h29 : _write_idx1_T_85; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_87 = _write_idx1_T[40] ? 6'h28 : _write_idx1_T_86; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_88 = _write_idx1_T[39] ? 6'h27 : _write_idx1_T_87; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_89 = _write_idx1_T[38] ? 6'h26 : _write_idx1_T_88; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_90 = _write_idx1_T[37] ? 6'h25 : _write_idx1_T_89; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_91 = _write_idx1_T[36] ? 6'h24 : _write_idx1_T_90; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_92 = _write_idx1_T[35] ? 6'h23 : _write_idx1_T_91; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_93 = _write_idx1_T[34] ? 6'h22 : _write_idx1_T_92; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_94 = _write_idx1_T[33] ? 6'h21 : _write_idx1_T_93; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_95 = _write_idx1_T[32] ? 6'h20 : _write_idx1_T_94; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_96 = _write_idx1_T[31] ? 6'h1f : _write_idx1_T_95; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_97 = _write_idx1_T[30] ? 6'h1e : _write_idx1_T_96; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_98 = _write_idx1_T[29] ? 6'h1d : _write_idx1_T_97; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_99 = _write_idx1_T[28] ? 6'h1c : _write_idx1_T_98; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_100 = _write_idx1_T[27] ? 6'h1b : _write_idx1_T_99; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_101 = _write_idx1_T[26] ? 6'h1a : _write_idx1_T_100; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_102 = _write_idx1_T[25] ? 6'h19 : _write_idx1_T_101; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_103 = _write_idx1_T[24] ? 6'h18 : _write_idx1_T_102; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_104 = _write_idx1_T[23] ? 6'h17 : _write_idx1_T_103; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_105 = _write_idx1_T[22] ? 6'h16 : _write_idx1_T_104; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_106 = _write_idx1_T[21] ? 6'h15 : _write_idx1_T_105; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_107 = _write_idx1_T[20] ? 6'h14 : _write_idx1_T_106; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_108 = _write_idx1_T[19] ? 6'h13 : _write_idx1_T_107; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_109 = _write_idx1_T[18] ? 6'h12 : _write_idx1_T_108; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_110 = _write_idx1_T[17] ? 6'h11 : _write_idx1_T_109; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_111 = _write_idx1_T[16] ? 6'h10 : _write_idx1_T_110; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_112 = _write_idx1_T[15] ? 6'hf : _write_idx1_T_111; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_113 = _write_idx1_T[14] ? 6'he : _write_idx1_T_112; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_114 = _write_idx1_T[13] ? 6'hd : _write_idx1_T_113; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_115 = _write_idx1_T[12] ? 6'hc : _write_idx1_T_114; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_116 = _write_idx1_T[11] ? 6'hb : _write_idx1_T_115; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_117 = _write_idx1_T[10] ? 6'ha : _write_idx1_T_116; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_118 = _write_idx1_T[9] ? 6'h9 : _write_idx1_T_117; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_119 = _write_idx1_T[8] ? 6'h8 : _write_idx1_T_118; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_120 = _write_idx1_T[7] ? 6'h7 : _write_idx1_T_119; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_121 = _write_idx1_T[6] ? 6'h6 : _write_idx1_T_120; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_122 = _write_idx1_T[5] ? 6'h5 : _write_idx1_T_121; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_123 = _write_idx1_T[4] ? 6'h4 : _write_idx1_T_122; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_124 = _write_idx1_T[3] ? 6'h3 : _write_idx1_T_123; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_125 = _write_idx1_T[2] ? 6'h2 : _write_idx1_T_124; // @[Mux.scala 47:70]
  wire [5:0] _write_idx1_T_126 = _write_idx1_T[1] ? 6'h1 : _write_idx1_T_125; // @[Mux.scala 47:70]
  wire [5:0] write_idx1 = _write_idx1_T[0] ? 6'h0 : _write_idx1_T_126; // @[Mux.scala 47:70]
  wire [63:0] _reservation_station_valid_withmask_T = 64'h1 << write_idx1; // @[OneHot.scala 57:35]
  wire [63:0] reservation_station_valid_withmask = reservation_station_valid | _reservation_station_valid_withmask_T; // @[reservation_station.scala 50:69]
  wire [63:0] _write_idx2_T = ~reservation_station_valid_withmask; // @[reservation_station.scala 51:34]
  wire [5:0] _write_idx2_T_65 = _write_idx2_T[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_66 = _write_idx2_T[61] ? 6'h3d : _write_idx2_T_65; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_67 = _write_idx2_T[60] ? 6'h3c : _write_idx2_T_66; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_68 = _write_idx2_T[59] ? 6'h3b : _write_idx2_T_67; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_69 = _write_idx2_T[58] ? 6'h3a : _write_idx2_T_68; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_70 = _write_idx2_T[57] ? 6'h39 : _write_idx2_T_69; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_71 = _write_idx2_T[56] ? 6'h38 : _write_idx2_T_70; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_72 = _write_idx2_T[55] ? 6'h37 : _write_idx2_T_71; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_73 = _write_idx2_T[54] ? 6'h36 : _write_idx2_T_72; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_74 = _write_idx2_T[53] ? 6'h35 : _write_idx2_T_73; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_75 = _write_idx2_T[52] ? 6'h34 : _write_idx2_T_74; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_76 = _write_idx2_T[51] ? 6'h33 : _write_idx2_T_75; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_77 = _write_idx2_T[50] ? 6'h32 : _write_idx2_T_76; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_78 = _write_idx2_T[49] ? 6'h31 : _write_idx2_T_77; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_79 = _write_idx2_T[48] ? 6'h30 : _write_idx2_T_78; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_80 = _write_idx2_T[47] ? 6'h2f : _write_idx2_T_79; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_81 = _write_idx2_T[46] ? 6'h2e : _write_idx2_T_80; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_82 = _write_idx2_T[45] ? 6'h2d : _write_idx2_T_81; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_83 = _write_idx2_T[44] ? 6'h2c : _write_idx2_T_82; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_84 = _write_idx2_T[43] ? 6'h2b : _write_idx2_T_83; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_85 = _write_idx2_T[42] ? 6'h2a : _write_idx2_T_84; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_86 = _write_idx2_T[41] ? 6'h29 : _write_idx2_T_85; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_87 = _write_idx2_T[40] ? 6'h28 : _write_idx2_T_86; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_88 = _write_idx2_T[39] ? 6'h27 : _write_idx2_T_87; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_89 = _write_idx2_T[38] ? 6'h26 : _write_idx2_T_88; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_90 = _write_idx2_T[37] ? 6'h25 : _write_idx2_T_89; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_91 = _write_idx2_T[36] ? 6'h24 : _write_idx2_T_90; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_92 = _write_idx2_T[35] ? 6'h23 : _write_idx2_T_91; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_93 = _write_idx2_T[34] ? 6'h22 : _write_idx2_T_92; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_94 = _write_idx2_T[33] ? 6'h21 : _write_idx2_T_93; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_95 = _write_idx2_T[32] ? 6'h20 : _write_idx2_T_94; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_96 = _write_idx2_T[31] ? 6'h1f : _write_idx2_T_95; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_97 = _write_idx2_T[30] ? 6'h1e : _write_idx2_T_96; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_98 = _write_idx2_T[29] ? 6'h1d : _write_idx2_T_97; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_99 = _write_idx2_T[28] ? 6'h1c : _write_idx2_T_98; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_100 = _write_idx2_T[27] ? 6'h1b : _write_idx2_T_99; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_101 = _write_idx2_T[26] ? 6'h1a : _write_idx2_T_100; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_102 = _write_idx2_T[25] ? 6'h19 : _write_idx2_T_101; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_103 = _write_idx2_T[24] ? 6'h18 : _write_idx2_T_102; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_104 = _write_idx2_T[23] ? 6'h17 : _write_idx2_T_103; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_105 = _write_idx2_T[22] ? 6'h16 : _write_idx2_T_104; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_106 = _write_idx2_T[21] ? 6'h15 : _write_idx2_T_105; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_107 = _write_idx2_T[20] ? 6'h14 : _write_idx2_T_106; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_108 = _write_idx2_T[19] ? 6'h13 : _write_idx2_T_107; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_109 = _write_idx2_T[18] ? 6'h12 : _write_idx2_T_108; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_110 = _write_idx2_T[17] ? 6'h11 : _write_idx2_T_109; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_111 = _write_idx2_T[16] ? 6'h10 : _write_idx2_T_110; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_112 = _write_idx2_T[15] ? 6'hf : _write_idx2_T_111; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_113 = _write_idx2_T[14] ? 6'he : _write_idx2_T_112; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_114 = _write_idx2_T[13] ? 6'hd : _write_idx2_T_113; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_115 = _write_idx2_T[12] ? 6'hc : _write_idx2_T_114; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_116 = _write_idx2_T[11] ? 6'hb : _write_idx2_T_115; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_117 = _write_idx2_T[10] ? 6'ha : _write_idx2_T_116; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_118 = _write_idx2_T[9] ? 6'h9 : _write_idx2_T_117; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_119 = _write_idx2_T[8] ? 6'h8 : _write_idx2_T_118; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_120 = _write_idx2_T[7] ? 6'h7 : _write_idx2_T_119; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_121 = _write_idx2_T[6] ? 6'h6 : _write_idx2_T_120; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_122 = _write_idx2_T[5] ? 6'h5 : _write_idx2_T_121; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_123 = _write_idx2_T[4] ? 6'h4 : _write_idx2_T_122; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_124 = _write_idx2_T[3] ? 6'h3 : _write_idx2_T_123; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_125 = _write_idx2_T[2] ? 6'h2 : _write_idx2_T_124; // @[Mux.scala 47:70]
  wire [5:0] _write_idx2_T_126 = _write_idx2_T[1] ? 6'h1 : _write_idx2_T_125; // @[Mux.scala 47:70]
  wire [5:0] write_idx2 = _write_idx2_T[0] ? 6'h0 : _write_idx2_T_126; // @[Mux.scala 47:70]
  wire  temp2_0 = |io_i_available_funcs_0; // @[reservation_station.scala 59:44]
  wire  temp2_1 = |io_i_available_funcs_1; // @[reservation_station.scala 59:44]
  wire  temp2_2 = |io_i_available_funcs_2; // @[reservation_station.scala 59:44]
  wire  temp2_3 = |io_i_available_funcs_3; // @[reservation_station.scala 59:44]
  wire  temp2_4 = |io_i_available_funcs_4; // @[reservation_station.scala 59:44]
  wire  temp2_5 = |io_i_available_funcs_5; // @[reservation_station.scala 59:44]
  wire [6:0] available_funcs = {1'h0,temp2_5,temp2_4,temp2_3,temp2_2,temp2_1,temp2_0}; // @[reservation_station.scala 61:37]
  wire [6:0] _slots_can_issue_T = reservation_station_0_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_0 = reservation_station_0_io_o_ready_to_issue & |_slots_can_issue_T; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_4 = reservation_station_1_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_1 = reservation_station_1_io_o_ready_to_issue & |_slots_can_issue_T_4; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_8 = reservation_station_2_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_2 = reservation_station_2_io_o_ready_to_issue & |_slots_can_issue_T_8; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_12 = reservation_station_3_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_3 = reservation_station_3_io_o_ready_to_issue & |_slots_can_issue_T_12; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_16 = reservation_station_4_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_4 = reservation_station_4_io_o_ready_to_issue & |_slots_can_issue_T_16; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_20 = reservation_station_5_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_5 = reservation_station_5_io_o_ready_to_issue & |_slots_can_issue_T_20; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_24 = reservation_station_6_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_6 = reservation_station_6_io_o_ready_to_issue & |_slots_can_issue_T_24; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_28 = reservation_station_7_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_7 = reservation_station_7_io_o_ready_to_issue & |_slots_can_issue_T_28; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_32 = reservation_station_8_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_8 = reservation_station_8_io_o_ready_to_issue & |_slots_can_issue_T_32; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_36 = reservation_station_9_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_9 = reservation_station_9_io_o_ready_to_issue & |_slots_can_issue_T_36; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_40 = reservation_station_10_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_10 = reservation_station_10_io_o_ready_to_issue & |_slots_can_issue_T_40; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_44 = reservation_station_11_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_11 = reservation_station_11_io_o_ready_to_issue & |_slots_can_issue_T_44; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_48 = reservation_station_12_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_12 = reservation_station_12_io_o_ready_to_issue & |_slots_can_issue_T_48; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_52 = reservation_station_13_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_13 = reservation_station_13_io_o_ready_to_issue & |_slots_can_issue_T_52; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_56 = reservation_station_14_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_14 = reservation_station_14_io_o_ready_to_issue & |_slots_can_issue_T_56; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_60 = reservation_station_15_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_15 = reservation_station_15_io_o_ready_to_issue & |_slots_can_issue_T_60; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_64 = reservation_station_16_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_16 = reservation_station_16_io_o_ready_to_issue & |_slots_can_issue_T_64; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_68 = reservation_station_17_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_17 = reservation_station_17_io_o_ready_to_issue & |_slots_can_issue_T_68; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_72 = reservation_station_18_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_18 = reservation_station_18_io_o_ready_to_issue & |_slots_can_issue_T_72; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_76 = reservation_station_19_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_19 = reservation_station_19_io_o_ready_to_issue & |_slots_can_issue_T_76; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_80 = reservation_station_20_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_20 = reservation_station_20_io_o_ready_to_issue & |_slots_can_issue_T_80; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_84 = reservation_station_21_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_21 = reservation_station_21_io_o_ready_to_issue & |_slots_can_issue_T_84; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_88 = reservation_station_22_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_22 = reservation_station_22_io_o_ready_to_issue & |_slots_can_issue_T_88; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_92 = reservation_station_23_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_23 = reservation_station_23_io_o_ready_to_issue & |_slots_can_issue_T_92; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_96 = reservation_station_24_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_24 = reservation_station_24_io_o_ready_to_issue & |_slots_can_issue_T_96; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_100 = reservation_station_25_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_25 = reservation_station_25_io_o_ready_to_issue & |_slots_can_issue_T_100; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_104 = reservation_station_26_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_26 = reservation_station_26_io_o_ready_to_issue & |_slots_can_issue_T_104; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_108 = reservation_station_27_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_27 = reservation_station_27_io_o_ready_to_issue & |_slots_can_issue_T_108; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_112 = reservation_station_28_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_28 = reservation_station_28_io_o_ready_to_issue & |_slots_can_issue_T_112; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_116 = reservation_station_29_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_29 = reservation_station_29_io_o_ready_to_issue & |_slots_can_issue_T_116; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_120 = reservation_station_30_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_30 = reservation_station_30_io_o_ready_to_issue & |_slots_can_issue_T_120; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_124 = reservation_station_31_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_31 = reservation_station_31_io_o_ready_to_issue & |_slots_can_issue_T_124; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_128 = reservation_station_32_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_32 = reservation_station_32_io_o_ready_to_issue & |_slots_can_issue_T_128; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_132 = reservation_station_33_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_33 = reservation_station_33_io_o_ready_to_issue & |_slots_can_issue_T_132; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_136 = reservation_station_34_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_34 = reservation_station_34_io_o_ready_to_issue & |_slots_can_issue_T_136; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_140 = reservation_station_35_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_35 = reservation_station_35_io_o_ready_to_issue & |_slots_can_issue_T_140; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_144 = reservation_station_36_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_36 = reservation_station_36_io_o_ready_to_issue & |_slots_can_issue_T_144; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_148 = reservation_station_37_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_37 = reservation_station_37_io_o_ready_to_issue & |_slots_can_issue_T_148; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_152 = reservation_station_38_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_38 = reservation_station_38_io_o_ready_to_issue & |_slots_can_issue_T_152; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_156 = reservation_station_39_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_39 = reservation_station_39_io_o_ready_to_issue & |_slots_can_issue_T_156; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_160 = reservation_station_40_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_40 = reservation_station_40_io_o_ready_to_issue & |_slots_can_issue_T_160; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_164 = reservation_station_41_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_41 = reservation_station_41_io_o_ready_to_issue & |_slots_can_issue_T_164; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_168 = reservation_station_42_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_42 = reservation_station_42_io_o_ready_to_issue & |_slots_can_issue_T_168; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_172 = reservation_station_43_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_43 = reservation_station_43_io_o_ready_to_issue & |_slots_can_issue_T_172; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_176 = reservation_station_44_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_44 = reservation_station_44_io_o_ready_to_issue & |_slots_can_issue_T_176; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_180 = reservation_station_45_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_45 = reservation_station_45_io_o_ready_to_issue & |_slots_can_issue_T_180; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_184 = reservation_station_46_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_46 = reservation_station_46_io_o_ready_to_issue & |_slots_can_issue_T_184; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_188 = reservation_station_47_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_47 = reservation_station_47_io_o_ready_to_issue & |_slots_can_issue_T_188; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_192 = reservation_station_48_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_48 = reservation_station_48_io_o_ready_to_issue & |_slots_can_issue_T_192; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_196 = reservation_station_49_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_49 = reservation_station_49_io_o_ready_to_issue & |_slots_can_issue_T_196; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_200 = reservation_station_50_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_50 = reservation_station_50_io_o_ready_to_issue & |_slots_can_issue_T_200; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_204 = reservation_station_51_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_51 = reservation_station_51_io_o_ready_to_issue & |_slots_can_issue_T_204; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_208 = reservation_station_52_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_52 = reservation_station_52_io_o_ready_to_issue & |_slots_can_issue_T_208; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_212 = reservation_station_53_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_53 = reservation_station_53_io_o_ready_to_issue & |_slots_can_issue_T_212; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_216 = reservation_station_54_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_54 = reservation_station_54_io_o_ready_to_issue & |_slots_can_issue_T_216; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_220 = reservation_station_55_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_55 = reservation_station_55_io_o_ready_to_issue & |_slots_can_issue_T_220; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_224 = reservation_station_56_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_56 = reservation_station_56_io_o_ready_to_issue & |_slots_can_issue_T_224; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_228 = reservation_station_57_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_57 = reservation_station_57_io_o_ready_to_issue & |_slots_can_issue_T_228; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_232 = reservation_station_58_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_58 = reservation_station_58_io_o_ready_to_issue & |_slots_can_issue_T_232; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_236 = reservation_station_59_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_59 = reservation_station_59_io_o_ready_to_issue & |_slots_can_issue_T_236; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_240 = reservation_station_60_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_60 = reservation_station_60_io_o_ready_to_issue & |_slots_can_issue_T_240; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_244 = reservation_station_61_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_61 = reservation_station_61_io_o_ready_to_issue & |_slots_can_issue_T_244; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_248 = reservation_station_62_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_62 = reservation_station_62_io_o_ready_to_issue & |_slots_can_issue_T_248; // @[reservation_station.scala 63:98]
  wire [6:0] _slots_can_issue_T_252 = reservation_station_63_io_o_uop_func_code & available_funcs; // @[reservation_station.scala 63:145]
  wire  slots_can_issue_63 = reservation_station_63_io_o_ready_to_issue & |_slots_can_issue_T_252; // @[reservation_station.scala 63:98]
  wire [7:0] issue1_idx_lo_lo_lo = {slots_can_issue_7,slots_can_issue_6,slots_can_issue_5,slots_can_issue_4,
    slots_can_issue_3,slots_can_issue_2,slots_can_issue_1,slots_can_issue_0}; // @[reservation_station.scala 65:58]
  wire [15:0] issue1_idx_lo_lo = {slots_can_issue_15,slots_can_issue_14,slots_can_issue_13,slots_can_issue_12,
    slots_can_issue_11,slots_can_issue_10,slots_can_issue_9,slots_can_issue_8,issue1_idx_lo_lo_lo}; // @[reservation_station.scala 65:58]
  wire [7:0] issue1_idx_lo_hi_lo = {slots_can_issue_23,slots_can_issue_22,slots_can_issue_21,slots_can_issue_20,
    slots_can_issue_19,slots_can_issue_18,slots_can_issue_17,slots_can_issue_16}; // @[reservation_station.scala 65:58]
  wire [31:0] issue1_idx_lo = {slots_can_issue_31,slots_can_issue_30,slots_can_issue_29,slots_can_issue_28,
    slots_can_issue_27,slots_can_issue_26,slots_can_issue_25,slots_can_issue_24,issue1_idx_lo_hi_lo,issue1_idx_lo_lo}; // @[reservation_station.scala 65:58]
  wire [7:0] issue1_idx_hi_lo_lo = {slots_can_issue_39,slots_can_issue_38,slots_can_issue_37,slots_can_issue_36,
    slots_can_issue_35,slots_can_issue_34,slots_can_issue_33,slots_can_issue_32}; // @[reservation_station.scala 65:58]
  wire [15:0] issue1_idx_hi_lo = {slots_can_issue_47,slots_can_issue_46,slots_can_issue_45,slots_can_issue_44,
    slots_can_issue_43,slots_can_issue_42,slots_can_issue_41,slots_can_issue_40,issue1_idx_hi_lo_lo}; // @[reservation_station.scala 65:58]
  wire [7:0] issue1_idx_hi_hi_lo = {slots_can_issue_55,slots_can_issue_54,slots_can_issue_53,slots_can_issue_52,
    slots_can_issue_51,slots_can_issue_50,slots_can_issue_49,slots_can_issue_48}; // @[reservation_station.scala 65:58]
  wire [31:0] issue1_idx_hi = {slots_can_issue_63,slots_can_issue_62,slots_can_issue_61,slots_can_issue_60,
    slots_can_issue_59,slots_can_issue_58,slots_can_issue_57,slots_can_issue_56,issue1_idx_hi_hi_lo,issue1_idx_hi_lo}; // @[reservation_station.scala 65:58]
  wire [63:0] _issue1_idx_T = {issue1_idx_hi,issue1_idx_lo}; // @[reservation_station.scala 65:58]
  wire [5:0] _issue1_idx_T_65 = _issue1_idx_T[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_66 = _issue1_idx_T[61] ? 6'h3d : _issue1_idx_T_65; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_67 = _issue1_idx_T[60] ? 6'h3c : _issue1_idx_T_66; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_68 = _issue1_idx_T[59] ? 6'h3b : _issue1_idx_T_67; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_69 = _issue1_idx_T[58] ? 6'h3a : _issue1_idx_T_68; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_70 = _issue1_idx_T[57] ? 6'h39 : _issue1_idx_T_69; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_71 = _issue1_idx_T[56] ? 6'h38 : _issue1_idx_T_70; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_72 = _issue1_idx_T[55] ? 6'h37 : _issue1_idx_T_71; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_73 = _issue1_idx_T[54] ? 6'h36 : _issue1_idx_T_72; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_74 = _issue1_idx_T[53] ? 6'h35 : _issue1_idx_T_73; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_75 = _issue1_idx_T[52] ? 6'h34 : _issue1_idx_T_74; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_76 = _issue1_idx_T[51] ? 6'h33 : _issue1_idx_T_75; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_77 = _issue1_idx_T[50] ? 6'h32 : _issue1_idx_T_76; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_78 = _issue1_idx_T[49] ? 6'h31 : _issue1_idx_T_77; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_79 = _issue1_idx_T[48] ? 6'h30 : _issue1_idx_T_78; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_80 = _issue1_idx_T[47] ? 6'h2f : _issue1_idx_T_79; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_81 = _issue1_idx_T[46] ? 6'h2e : _issue1_idx_T_80; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_82 = _issue1_idx_T[45] ? 6'h2d : _issue1_idx_T_81; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_83 = _issue1_idx_T[44] ? 6'h2c : _issue1_idx_T_82; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_84 = _issue1_idx_T[43] ? 6'h2b : _issue1_idx_T_83; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_85 = _issue1_idx_T[42] ? 6'h2a : _issue1_idx_T_84; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_86 = _issue1_idx_T[41] ? 6'h29 : _issue1_idx_T_85; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_87 = _issue1_idx_T[40] ? 6'h28 : _issue1_idx_T_86; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_88 = _issue1_idx_T[39] ? 6'h27 : _issue1_idx_T_87; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_89 = _issue1_idx_T[38] ? 6'h26 : _issue1_idx_T_88; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_90 = _issue1_idx_T[37] ? 6'h25 : _issue1_idx_T_89; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_91 = _issue1_idx_T[36] ? 6'h24 : _issue1_idx_T_90; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_92 = _issue1_idx_T[35] ? 6'h23 : _issue1_idx_T_91; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_93 = _issue1_idx_T[34] ? 6'h22 : _issue1_idx_T_92; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_94 = _issue1_idx_T[33] ? 6'h21 : _issue1_idx_T_93; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_95 = _issue1_idx_T[32] ? 6'h20 : _issue1_idx_T_94; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_96 = _issue1_idx_T[31] ? 6'h1f : _issue1_idx_T_95; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_97 = _issue1_idx_T[30] ? 6'h1e : _issue1_idx_T_96; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_98 = _issue1_idx_T[29] ? 6'h1d : _issue1_idx_T_97; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_99 = _issue1_idx_T[28] ? 6'h1c : _issue1_idx_T_98; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_100 = _issue1_idx_T[27] ? 6'h1b : _issue1_idx_T_99; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_101 = _issue1_idx_T[26] ? 6'h1a : _issue1_idx_T_100; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_102 = _issue1_idx_T[25] ? 6'h19 : _issue1_idx_T_101; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_103 = _issue1_idx_T[24] ? 6'h18 : _issue1_idx_T_102; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_104 = _issue1_idx_T[23] ? 6'h17 : _issue1_idx_T_103; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_105 = _issue1_idx_T[22] ? 6'h16 : _issue1_idx_T_104; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_106 = _issue1_idx_T[21] ? 6'h15 : _issue1_idx_T_105; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_107 = _issue1_idx_T[20] ? 6'h14 : _issue1_idx_T_106; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_108 = _issue1_idx_T[19] ? 6'h13 : _issue1_idx_T_107; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_109 = _issue1_idx_T[18] ? 6'h12 : _issue1_idx_T_108; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_110 = _issue1_idx_T[17] ? 6'h11 : _issue1_idx_T_109; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_111 = _issue1_idx_T[16] ? 6'h10 : _issue1_idx_T_110; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_112 = _issue1_idx_T[15] ? 6'hf : _issue1_idx_T_111; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_113 = _issue1_idx_T[14] ? 6'he : _issue1_idx_T_112; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_114 = _issue1_idx_T[13] ? 6'hd : _issue1_idx_T_113; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_115 = _issue1_idx_T[12] ? 6'hc : _issue1_idx_T_114; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_116 = _issue1_idx_T[11] ? 6'hb : _issue1_idx_T_115; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_117 = _issue1_idx_T[10] ? 6'ha : _issue1_idx_T_116; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_118 = _issue1_idx_T[9] ? 6'h9 : _issue1_idx_T_117; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_119 = _issue1_idx_T[8] ? 6'h8 : _issue1_idx_T_118; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_120 = _issue1_idx_T[7] ? 6'h7 : _issue1_idx_T_119; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_121 = _issue1_idx_T[6] ? 6'h6 : _issue1_idx_T_120; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_122 = _issue1_idx_T[5] ? 6'h5 : _issue1_idx_T_121; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_123 = _issue1_idx_T[4] ? 6'h4 : _issue1_idx_T_122; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_124 = _issue1_idx_T[3] ? 6'h3 : _issue1_idx_T_123; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_125 = _issue1_idx_T[2] ? 6'h2 : _issue1_idx_T_124; // @[Mux.scala 47:70]
  wire [5:0] _issue1_idx_T_126 = _issue1_idx_T[1] ? 6'h1 : _issue1_idx_T_125; // @[Mux.scala 47:70]
  wire [5:0] issue1_idx = _issue1_idx_T[0] ? 6'h0 : _issue1_idx_T_126; // @[Mux.scala 47:70]
  wire  _issue1_func_code_T = 6'h0 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_1 = 6'h1 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_2 = 6'h2 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_3 = 6'h3 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_4 = 6'h4 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_5 = 6'h5 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_6 = 6'h6 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_7 = 6'h7 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_8 = 6'h8 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_9 = 6'h9 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_10 = 6'ha == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_11 = 6'hb == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_12 = 6'hc == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_13 = 6'hd == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_14 = 6'he == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_15 = 6'hf == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_16 = 6'h10 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_17 = 6'h11 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_18 = 6'h12 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_19 = 6'h13 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_20 = 6'h14 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_21 = 6'h15 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_22 = 6'h16 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_23 = 6'h17 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_24 = 6'h18 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_25 = 6'h19 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_26 = 6'h1a == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_27 = 6'h1b == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_28 = 6'h1c == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_29 = 6'h1d == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_30 = 6'h1e == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_31 = 6'h1f == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_32 = 6'h20 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_33 = 6'h21 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_34 = 6'h22 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_35 = 6'h23 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_36 = 6'h24 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_37 = 6'h25 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_38 = 6'h26 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_39 = 6'h27 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_40 = 6'h28 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_41 = 6'h29 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_42 = 6'h2a == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_43 = 6'h2b == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_44 = 6'h2c == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_45 = 6'h2d == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_46 = 6'h2e == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_47 = 6'h2f == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_48 = 6'h30 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_49 = 6'h31 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_50 = 6'h32 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_51 = 6'h33 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_52 = 6'h34 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_53 = 6'h35 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_54 = 6'h36 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_55 = 6'h37 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_56 = 6'h38 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_57 = 6'h39 == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_58 = 6'h3a == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_59 = 6'h3b == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_60 = 6'h3c == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_61 = 6'h3d == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_62 = 6'h3e == issue1_idx; // @[reservation_station.scala 68:80]
  wire  _issue1_func_code_T_63 = 6'h3f == issue1_idx; // @[reservation_station.scala 68:80]
  wire [6:0] _issue1_func_code_T_64 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_func_code : 7'h40; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_65 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_func_code :
    _issue1_func_code_T_64; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_66 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_func_code :
    _issue1_func_code_T_65; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_67 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_func_code :
    _issue1_func_code_T_66; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_68 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_func_code :
    _issue1_func_code_T_67; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_69 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_func_code :
    _issue1_func_code_T_68; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_70 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_func_code :
    _issue1_func_code_T_69; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_71 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_func_code :
    _issue1_func_code_T_70; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_72 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_func_code :
    _issue1_func_code_T_71; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_73 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_func_code :
    _issue1_func_code_T_72; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_74 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_func_code :
    _issue1_func_code_T_73; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_75 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_func_code :
    _issue1_func_code_T_74; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_76 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_func_code :
    _issue1_func_code_T_75; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_77 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_func_code :
    _issue1_func_code_T_76; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_78 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_func_code :
    _issue1_func_code_T_77; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_79 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_func_code :
    _issue1_func_code_T_78; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_80 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_func_code :
    _issue1_func_code_T_79; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_81 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_func_code :
    _issue1_func_code_T_80; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_82 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_func_code :
    _issue1_func_code_T_81; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_83 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_func_code :
    _issue1_func_code_T_82; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_84 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_func_code :
    _issue1_func_code_T_83; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_85 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_func_code :
    _issue1_func_code_T_84; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_86 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_func_code :
    _issue1_func_code_T_85; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_87 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_func_code :
    _issue1_func_code_T_86; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_88 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_func_code :
    _issue1_func_code_T_87; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_89 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_func_code :
    _issue1_func_code_T_88; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_90 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_func_code :
    _issue1_func_code_T_89; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_91 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_func_code :
    _issue1_func_code_T_90; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_92 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_func_code :
    _issue1_func_code_T_91; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_93 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_func_code :
    _issue1_func_code_T_92; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_94 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_func_code :
    _issue1_func_code_T_93; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_95 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_func_code :
    _issue1_func_code_T_94; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_96 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_func_code :
    _issue1_func_code_T_95; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_97 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_func_code :
    _issue1_func_code_T_96; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_98 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_func_code :
    _issue1_func_code_T_97; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_99 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_func_code :
    _issue1_func_code_T_98; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_100 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_func_code :
    _issue1_func_code_T_99; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_101 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_func_code :
    _issue1_func_code_T_100; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_102 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_func_code :
    _issue1_func_code_T_101; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_103 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_func_code :
    _issue1_func_code_T_102; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_104 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_func_code :
    _issue1_func_code_T_103; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_105 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_func_code :
    _issue1_func_code_T_104; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_106 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_func_code :
    _issue1_func_code_T_105; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_107 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_func_code :
    _issue1_func_code_T_106; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_108 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_func_code :
    _issue1_func_code_T_107; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_109 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_func_code :
    _issue1_func_code_T_108; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_110 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_func_code :
    _issue1_func_code_T_109; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_111 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_func_code :
    _issue1_func_code_T_110; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_112 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_func_code :
    _issue1_func_code_T_111; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_113 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_func_code :
    _issue1_func_code_T_112; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_114 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_func_code :
    _issue1_func_code_T_113; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_115 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_func_code :
    _issue1_func_code_T_114; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_116 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_func_code :
    _issue1_func_code_T_115; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_117 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_func_code :
    _issue1_func_code_T_116; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_118 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_func_code :
    _issue1_func_code_T_117; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_119 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_func_code :
    _issue1_func_code_T_118; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_120 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_func_code :
    _issue1_func_code_T_119; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_121 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_func_code :
    _issue1_func_code_T_120; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_122 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_func_code :
    _issue1_func_code_T_121; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_123 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_func_code :
    _issue1_func_code_T_122; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_124 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_func_code :
    _issue1_func_code_T_123; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_125 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_func_code :
    _issue1_func_code_T_124; // @[Mux.scala 101:16]
  wire [6:0] _issue1_func_code_T_126 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_func_code :
    _issue1_func_code_T_125; // @[Mux.scala 101:16]
  wire [6:0] issue1_func_code = _issue1_func_code_T ? reservation_station_0_io_o_uop_func_code : _issue1_func_code_T_126
    ; // @[Mux.scala 101:16]
  wire [2:0] hi = issue1_func_code[6:4]; // @[OneHot.scala 30:18]
  wire [3:0] lo = issue1_func_code[3:0]; // @[OneHot.scala 31:18]
  wire  _T = |hi; // @[OneHot.scala 32:14]
  wire [3:0] _GEN_14 = {{1'd0}, hi}; // @[OneHot.scala 32:28]
  wire [3:0] _T_1 = _GEN_14 | lo; // @[OneHot.scala 32:28]
  wire [1:0] hi_1 = _T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_1 = _T_1[1:0]; // @[OneHot.scala 31:18]
  wire  _T_2 = |hi_1; // @[OneHot.scala 32:14]
  wire [1:0] _T_3 = hi_1 | lo_1; // @[OneHot.scala 32:28]
  wire [2:0] _T_6 = {_T,_T_2,_T_3[1]}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_1 = 3'h1 == _T_6 ? io_i_available_funcs_1 : io_i_available_funcs_0; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_2 = 3'h2 == _T_6 ? io_i_available_funcs_2 : _GEN_1; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_3 = 3'h3 == _T_6 ? io_i_available_funcs_3 : _GEN_2; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_4 = 3'h4 == _T_6 ? io_i_available_funcs_4 : _GEN_3; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_5 = 3'h5 == _T_6 ? io_i_available_funcs_5 : _GEN_4; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _GEN_6 = 3'h6 == _T_6 ? 2'h0 : _GEN_5; // @[reservation_station.scala 71:{109,109}]
  wire [1:0] _available_funcs_with_mask_T_8 = _GEN_6 - 2'h1; // @[reservation_station.scala 71:109]
  wire [1:0] available_funcs_with_mask_0 = 3'h0 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_0; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_1 = 3'h1 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_1; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_2 = 3'h2 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_2; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_3 = 3'h3 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_3; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_4 = 3'h4 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_4; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_5 = 3'h5 == _T_6 ? _available_funcs_with_mask_T_8 : io_i_available_funcs_5; // @[reservation_station.scala 70:31 71:{59,59}]
  wire [1:0] available_funcs_with_mask_6 = 3'h6 == _T_6 ? _available_funcs_with_mask_T_8 : 2'h0; // @[reservation_station.scala 70:31 71:{59,59}]
  wire  temp3_0 = |available_funcs_with_mask_0; // @[reservation_station.scala 75:49]
  wire  temp3_1 = |available_funcs_with_mask_1; // @[reservation_station.scala 75:49]
  wire  temp3_2 = |available_funcs_with_mask_2; // @[reservation_station.scala 75:49]
  wire  temp3_3 = |available_funcs_with_mask_3; // @[reservation_station.scala 75:49]
  wire  temp3_4 = |available_funcs_with_mask_4; // @[reservation_station.scala 75:49]
  wire  temp3_5 = |available_funcs_with_mask_5; // @[reservation_station.scala 75:49]
  wire  temp3_6 = |available_funcs_with_mask_6; // @[reservation_station.scala 75:49]
  wire [6:0] available_funcs2_bits = {temp3_6,temp3_5,temp3_4,temp3_3,temp3_2,temp3_1,temp3_0}; // @[reservation_station.scala 78:46]
  wire [6:0] _slots_can_issue2_T_2 = reservation_station_0_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_3 = |_slots_can_issue2_T_2; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_0 = slots_can_issue_0 & 6'h0 != issue1_idx & _slots_can_issue2_T_3; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_8 = reservation_station_1_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_9 = |_slots_can_issue2_T_8; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_1 = slots_can_issue_1 & 6'h1 != issue1_idx & _slots_can_issue2_T_9; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_14 = reservation_station_2_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_15 = |_slots_can_issue2_T_14; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_2 = slots_can_issue_2 & 6'h2 != issue1_idx & _slots_can_issue2_T_15; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_20 = reservation_station_3_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_21 = |_slots_can_issue2_T_20; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_3 = slots_can_issue_3 & 6'h3 != issue1_idx & _slots_can_issue2_T_21; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_26 = reservation_station_4_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_27 = |_slots_can_issue2_T_26; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_4 = slots_can_issue_4 & 6'h4 != issue1_idx & _slots_can_issue2_T_27; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_32 = reservation_station_5_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_33 = |_slots_can_issue2_T_32; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_5 = slots_can_issue_5 & 6'h5 != issue1_idx & _slots_can_issue2_T_33; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_38 = reservation_station_6_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_39 = |_slots_can_issue2_T_38; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_6 = slots_can_issue_6 & 6'h6 != issue1_idx & _slots_can_issue2_T_39; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_44 = reservation_station_7_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_45 = |_slots_can_issue2_T_44; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_7 = slots_can_issue_7 & 6'h7 != issue1_idx & _slots_can_issue2_T_45; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_50 = reservation_station_8_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_51 = |_slots_can_issue2_T_50; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_8 = slots_can_issue_8 & 6'h8 != issue1_idx & _slots_can_issue2_T_51; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_56 = reservation_station_9_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_57 = |_slots_can_issue2_T_56; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_9 = slots_can_issue_9 & 6'h9 != issue1_idx & _slots_can_issue2_T_57; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_62 = reservation_station_10_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_63 = |_slots_can_issue2_T_62; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_10 = slots_can_issue_10 & 6'ha != issue1_idx & _slots_can_issue2_T_63; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_68 = reservation_station_11_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_69 = |_slots_can_issue2_T_68; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_11 = slots_can_issue_11 & 6'hb != issue1_idx & _slots_can_issue2_T_69; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_74 = reservation_station_12_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_75 = |_slots_can_issue2_T_74; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_12 = slots_can_issue_12 & 6'hc != issue1_idx & _slots_can_issue2_T_75; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_80 = reservation_station_13_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_81 = |_slots_can_issue2_T_80; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_13 = slots_can_issue_13 & 6'hd != issue1_idx & _slots_can_issue2_T_81; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_86 = reservation_station_14_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_87 = |_slots_can_issue2_T_86; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_14 = slots_can_issue_14 & 6'he != issue1_idx & _slots_can_issue2_T_87; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_92 = reservation_station_15_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_93 = |_slots_can_issue2_T_92; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_15 = slots_can_issue_15 & 6'hf != issue1_idx & _slots_can_issue2_T_93; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_98 = reservation_station_16_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_99 = |_slots_can_issue2_T_98; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_16 = slots_can_issue_16 & 6'h10 != issue1_idx & _slots_can_issue2_T_99; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_104 = reservation_station_17_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_105 = |_slots_can_issue2_T_104; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_17 = slots_can_issue_17 & 6'h11 != issue1_idx & _slots_can_issue2_T_105; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_110 = reservation_station_18_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_111 = |_slots_can_issue2_T_110; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_18 = slots_can_issue_18 & 6'h12 != issue1_idx & _slots_can_issue2_T_111; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_116 = reservation_station_19_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_117 = |_slots_can_issue2_T_116; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_19 = slots_can_issue_19 & 6'h13 != issue1_idx & _slots_can_issue2_T_117; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_122 = reservation_station_20_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_123 = |_slots_can_issue2_T_122; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_20 = slots_can_issue_20 & 6'h14 != issue1_idx & _slots_can_issue2_T_123; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_128 = reservation_station_21_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_129 = |_slots_can_issue2_T_128; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_21 = slots_can_issue_21 & 6'h15 != issue1_idx & _slots_can_issue2_T_129; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_134 = reservation_station_22_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_135 = |_slots_can_issue2_T_134; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_22 = slots_can_issue_22 & 6'h16 != issue1_idx & _slots_can_issue2_T_135; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_140 = reservation_station_23_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_141 = |_slots_can_issue2_T_140; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_23 = slots_can_issue_23 & 6'h17 != issue1_idx & _slots_can_issue2_T_141; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_146 = reservation_station_24_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_147 = |_slots_can_issue2_T_146; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_24 = slots_can_issue_24 & 6'h18 != issue1_idx & _slots_can_issue2_T_147; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_152 = reservation_station_25_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_153 = |_slots_can_issue2_T_152; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_25 = slots_can_issue_25 & 6'h19 != issue1_idx & _slots_can_issue2_T_153; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_158 = reservation_station_26_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_159 = |_slots_can_issue2_T_158; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_26 = slots_can_issue_26 & 6'h1a != issue1_idx & _slots_can_issue2_T_159; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_164 = reservation_station_27_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_165 = |_slots_can_issue2_T_164; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_27 = slots_can_issue_27 & 6'h1b != issue1_idx & _slots_can_issue2_T_165; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_170 = reservation_station_28_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_171 = |_slots_can_issue2_T_170; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_28 = slots_can_issue_28 & 6'h1c != issue1_idx & _slots_can_issue2_T_171; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_176 = reservation_station_29_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_177 = |_slots_can_issue2_T_176; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_29 = slots_can_issue_29 & 6'h1d != issue1_idx & _slots_can_issue2_T_177; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_182 = reservation_station_30_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_183 = |_slots_can_issue2_T_182; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_30 = slots_can_issue_30 & 6'h1e != issue1_idx & _slots_can_issue2_T_183; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_188 = reservation_station_31_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_189 = |_slots_can_issue2_T_188; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_31 = slots_can_issue_31 & 6'h1f != issue1_idx & _slots_can_issue2_T_189; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_194 = reservation_station_32_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_195 = |_slots_can_issue2_T_194; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_32 = slots_can_issue_32 & 6'h20 != issue1_idx & _slots_can_issue2_T_195; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_200 = reservation_station_33_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_201 = |_slots_can_issue2_T_200; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_33 = slots_can_issue_33 & 6'h21 != issue1_idx & _slots_can_issue2_T_201; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_206 = reservation_station_34_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_207 = |_slots_can_issue2_T_206; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_34 = slots_can_issue_34 & 6'h22 != issue1_idx & _slots_can_issue2_T_207; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_212 = reservation_station_35_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_213 = |_slots_can_issue2_T_212; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_35 = slots_can_issue_35 & 6'h23 != issue1_idx & _slots_can_issue2_T_213; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_218 = reservation_station_36_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_219 = |_slots_can_issue2_T_218; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_36 = slots_can_issue_36 & 6'h24 != issue1_idx & _slots_can_issue2_T_219; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_224 = reservation_station_37_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_225 = |_slots_can_issue2_T_224; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_37 = slots_can_issue_37 & 6'h25 != issue1_idx & _slots_can_issue2_T_225; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_230 = reservation_station_38_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_231 = |_slots_can_issue2_T_230; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_38 = slots_can_issue_38 & 6'h26 != issue1_idx & _slots_can_issue2_T_231; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_236 = reservation_station_39_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_237 = |_slots_can_issue2_T_236; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_39 = slots_can_issue_39 & 6'h27 != issue1_idx & _slots_can_issue2_T_237; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_242 = reservation_station_40_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_243 = |_slots_can_issue2_T_242; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_40 = slots_can_issue_40 & 6'h28 != issue1_idx & _slots_can_issue2_T_243; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_248 = reservation_station_41_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_249 = |_slots_can_issue2_T_248; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_41 = slots_can_issue_41 & 6'h29 != issue1_idx & _slots_can_issue2_T_249; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_254 = reservation_station_42_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_255 = |_slots_can_issue2_T_254; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_42 = slots_can_issue_42 & 6'h2a != issue1_idx & _slots_can_issue2_T_255; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_260 = reservation_station_43_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_261 = |_slots_can_issue2_T_260; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_43 = slots_can_issue_43 & 6'h2b != issue1_idx & _slots_can_issue2_T_261; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_266 = reservation_station_44_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_267 = |_slots_can_issue2_T_266; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_44 = slots_can_issue_44 & 6'h2c != issue1_idx & _slots_can_issue2_T_267; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_272 = reservation_station_45_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_273 = |_slots_can_issue2_T_272; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_45 = slots_can_issue_45 & 6'h2d != issue1_idx & _slots_can_issue2_T_273; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_278 = reservation_station_46_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_279 = |_slots_can_issue2_T_278; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_46 = slots_can_issue_46 & 6'h2e != issue1_idx & _slots_can_issue2_T_279; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_284 = reservation_station_47_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_285 = |_slots_can_issue2_T_284; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_47 = slots_can_issue_47 & 6'h2f != issue1_idx & _slots_can_issue2_T_285; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_290 = reservation_station_48_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_291 = |_slots_can_issue2_T_290; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_48 = slots_can_issue_48 & 6'h30 != issue1_idx & _slots_can_issue2_T_291; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_296 = reservation_station_49_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_297 = |_slots_can_issue2_T_296; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_49 = slots_can_issue_49 & 6'h31 != issue1_idx & _slots_can_issue2_T_297; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_302 = reservation_station_50_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_303 = |_slots_can_issue2_T_302; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_50 = slots_can_issue_50 & 6'h32 != issue1_idx & _slots_can_issue2_T_303; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_308 = reservation_station_51_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_309 = |_slots_can_issue2_T_308; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_51 = slots_can_issue_51 & 6'h33 != issue1_idx & _slots_can_issue2_T_309; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_314 = reservation_station_52_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_315 = |_slots_can_issue2_T_314; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_52 = slots_can_issue_52 & 6'h34 != issue1_idx & _slots_can_issue2_T_315; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_320 = reservation_station_53_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_321 = |_slots_can_issue2_T_320; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_53 = slots_can_issue_53 & 6'h35 != issue1_idx & _slots_can_issue2_T_321; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_326 = reservation_station_54_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_327 = |_slots_can_issue2_T_326; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_54 = slots_can_issue_54 & 6'h36 != issue1_idx & _slots_can_issue2_T_327; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_332 = reservation_station_55_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_333 = |_slots_can_issue2_T_332; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_55 = slots_can_issue_55 & 6'h37 != issue1_idx & _slots_can_issue2_T_333; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_338 = reservation_station_56_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_339 = |_slots_can_issue2_T_338; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_56 = slots_can_issue_56 & 6'h38 != issue1_idx & _slots_can_issue2_T_339; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_344 = reservation_station_57_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_345 = |_slots_can_issue2_T_344; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_57 = slots_can_issue_57 & 6'h39 != issue1_idx & _slots_can_issue2_T_345; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_350 = reservation_station_58_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_351 = |_slots_can_issue2_T_350; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_58 = slots_can_issue_58 & 6'h3a != issue1_idx & _slots_can_issue2_T_351; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_356 = reservation_station_59_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_357 = |_slots_can_issue2_T_356; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_59 = slots_can_issue_59 & 6'h3b != issue1_idx & _slots_can_issue2_T_357; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_362 = reservation_station_60_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_363 = |_slots_can_issue2_T_362; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_60 = slots_can_issue_60 & 6'h3c != issue1_idx & _slots_can_issue2_T_363; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_368 = reservation_station_61_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_369 = |_slots_can_issue2_T_368; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_61 = slots_can_issue_61 & 6'h3d != issue1_idx & _slots_can_issue2_T_369; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_374 = reservation_station_62_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_375 = |_slots_can_issue2_T_374; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_62 = slots_can_issue_62 & 6'h3e != issue1_idx & _slots_can_issue2_T_375; // @[reservation_station.scala 79:99]
  wire [6:0] _slots_can_issue2_T_380 = reservation_station_63_io_o_uop_func_code & available_funcs2_bits; // @[reservation_station.scala 80:55]
  wire  _slots_can_issue2_T_381 = |_slots_can_issue2_T_380; // @[reservation_station.scala 80:80]
  wire  slots_can_issue2_63 = slots_can_issue_63 & 6'h3f != issue1_idx & _slots_can_issue2_T_381; // @[reservation_station.scala 79:99]
  wire [7:0] issue2_idx_lo_lo_lo = {slots_can_issue2_7,slots_can_issue2_6,slots_can_issue2_5,slots_can_issue2_4,
    slots_can_issue2_3,slots_can_issue2_2,slots_can_issue2_1,slots_can_issue2_0}; // @[reservation_station.scala 83:53]
  wire [15:0] issue2_idx_lo_lo = {slots_can_issue2_15,slots_can_issue2_14,slots_can_issue2_13,slots_can_issue2_12,
    slots_can_issue2_11,slots_can_issue2_10,slots_can_issue2_9,slots_can_issue2_8,issue2_idx_lo_lo_lo}; // @[reservation_station.scala 83:53]
  wire [7:0] issue2_idx_lo_hi_lo = {slots_can_issue2_23,slots_can_issue2_22,slots_can_issue2_21,slots_can_issue2_20,
    slots_can_issue2_19,slots_can_issue2_18,slots_can_issue2_17,slots_can_issue2_16}; // @[reservation_station.scala 83:53]
  wire [31:0] issue2_idx_lo = {slots_can_issue2_31,slots_can_issue2_30,slots_can_issue2_29,slots_can_issue2_28,
    slots_can_issue2_27,slots_can_issue2_26,slots_can_issue2_25,slots_can_issue2_24,issue2_idx_lo_hi_lo,issue2_idx_lo_lo
    }; // @[reservation_station.scala 83:53]
  wire [7:0] issue2_idx_hi_lo_lo = {slots_can_issue2_39,slots_can_issue2_38,slots_can_issue2_37,slots_can_issue2_36,
    slots_can_issue2_35,slots_can_issue2_34,slots_can_issue2_33,slots_can_issue2_32}; // @[reservation_station.scala 83:53]
  wire [15:0] issue2_idx_hi_lo = {slots_can_issue2_47,slots_can_issue2_46,slots_can_issue2_45,slots_can_issue2_44,
    slots_can_issue2_43,slots_can_issue2_42,slots_can_issue2_41,slots_can_issue2_40,issue2_idx_hi_lo_lo}; // @[reservation_station.scala 83:53]
  wire [7:0] issue2_idx_hi_hi_lo = {slots_can_issue2_55,slots_can_issue2_54,slots_can_issue2_53,slots_can_issue2_52,
    slots_can_issue2_51,slots_can_issue2_50,slots_can_issue2_49,slots_can_issue2_48}; // @[reservation_station.scala 83:53]
  wire [31:0] issue2_idx_hi = {slots_can_issue2_63,slots_can_issue2_62,slots_can_issue2_61,slots_can_issue2_60,
    slots_can_issue2_59,slots_can_issue2_58,slots_can_issue2_57,slots_can_issue2_56,issue2_idx_hi_hi_lo,issue2_idx_hi_lo
    }; // @[reservation_station.scala 83:53]
  wire [63:0] _issue2_idx_T = {issue2_idx_hi,issue2_idx_lo}; // @[reservation_station.scala 83:53]
  wire [5:0] _issue2_idx_T_65 = _issue2_idx_T[62] ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_66 = _issue2_idx_T[61] ? 6'h3d : _issue2_idx_T_65; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_67 = _issue2_idx_T[60] ? 6'h3c : _issue2_idx_T_66; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_68 = _issue2_idx_T[59] ? 6'h3b : _issue2_idx_T_67; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_69 = _issue2_idx_T[58] ? 6'h3a : _issue2_idx_T_68; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_70 = _issue2_idx_T[57] ? 6'h39 : _issue2_idx_T_69; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_71 = _issue2_idx_T[56] ? 6'h38 : _issue2_idx_T_70; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_72 = _issue2_idx_T[55] ? 6'h37 : _issue2_idx_T_71; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_73 = _issue2_idx_T[54] ? 6'h36 : _issue2_idx_T_72; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_74 = _issue2_idx_T[53] ? 6'h35 : _issue2_idx_T_73; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_75 = _issue2_idx_T[52] ? 6'h34 : _issue2_idx_T_74; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_76 = _issue2_idx_T[51] ? 6'h33 : _issue2_idx_T_75; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_77 = _issue2_idx_T[50] ? 6'h32 : _issue2_idx_T_76; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_78 = _issue2_idx_T[49] ? 6'h31 : _issue2_idx_T_77; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_79 = _issue2_idx_T[48] ? 6'h30 : _issue2_idx_T_78; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_80 = _issue2_idx_T[47] ? 6'h2f : _issue2_idx_T_79; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_81 = _issue2_idx_T[46] ? 6'h2e : _issue2_idx_T_80; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_82 = _issue2_idx_T[45] ? 6'h2d : _issue2_idx_T_81; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_83 = _issue2_idx_T[44] ? 6'h2c : _issue2_idx_T_82; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_84 = _issue2_idx_T[43] ? 6'h2b : _issue2_idx_T_83; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_85 = _issue2_idx_T[42] ? 6'h2a : _issue2_idx_T_84; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_86 = _issue2_idx_T[41] ? 6'h29 : _issue2_idx_T_85; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_87 = _issue2_idx_T[40] ? 6'h28 : _issue2_idx_T_86; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_88 = _issue2_idx_T[39] ? 6'h27 : _issue2_idx_T_87; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_89 = _issue2_idx_T[38] ? 6'h26 : _issue2_idx_T_88; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_90 = _issue2_idx_T[37] ? 6'h25 : _issue2_idx_T_89; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_91 = _issue2_idx_T[36] ? 6'h24 : _issue2_idx_T_90; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_92 = _issue2_idx_T[35] ? 6'h23 : _issue2_idx_T_91; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_93 = _issue2_idx_T[34] ? 6'h22 : _issue2_idx_T_92; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_94 = _issue2_idx_T[33] ? 6'h21 : _issue2_idx_T_93; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_95 = _issue2_idx_T[32] ? 6'h20 : _issue2_idx_T_94; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_96 = _issue2_idx_T[31] ? 6'h1f : _issue2_idx_T_95; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_97 = _issue2_idx_T[30] ? 6'h1e : _issue2_idx_T_96; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_98 = _issue2_idx_T[29] ? 6'h1d : _issue2_idx_T_97; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_99 = _issue2_idx_T[28] ? 6'h1c : _issue2_idx_T_98; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_100 = _issue2_idx_T[27] ? 6'h1b : _issue2_idx_T_99; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_101 = _issue2_idx_T[26] ? 6'h1a : _issue2_idx_T_100; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_102 = _issue2_idx_T[25] ? 6'h19 : _issue2_idx_T_101; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_103 = _issue2_idx_T[24] ? 6'h18 : _issue2_idx_T_102; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_104 = _issue2_idx_T[23] ? 6'h17 : _issue2_idx_T_103; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_105 = _issue2_idx_T[22] ? 6'h16 : _issue2_idx_T_104; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_106 = _issue2_idx_T[21] ? 6'h15 : _issue2_idx_T_105; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_107 = _issue2_idx_T[20] ? 6'h14 : _issue2_idx_T_106; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_108 = _issue2_idx_T[19] ? 6'h13 : _issue2_idx_T_107; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_109 = _issue2_idx_T[18] ? 6'h12 : _issue2_idx_T_108; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_110 = _issue2_idx_T[17] ? 6'h11 : _issue2_idx_T_109; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_111 = _issue2_idx_T[16] ? 6'h10 : _issue2_idx_T_110; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_112 = _issue2_idx_T[15] ? 6'hf : _issue2_idx_T_111; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_113 = _issue2_idx_T[14] ? 6'he : _issue2_idx_T_112; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_114 = _issue2_idx_T[13] ? 6'hd : _issue2_idx_T_113; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_115 = _issue2_idx_T[12] ? 6'hc : _issue2_idx_T_114; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_116 = _issue2_idx_T[11] ? 6'hb : _issue2_idx_T_115; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_117 = _issue2_idx_T[10] ? 6'ha : _issue2_idx_T_116; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_118 = _issue2_idx_T[9] ? 6'h9 : _issue2_idx_T_117; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_119 = _issue2_idx_T[8] ? 6'h8 : _issue2_idx_T_118; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_120 = _issue2_idx_T[7] ? 6'h7 : _issue2_idx_T_119; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_121 = _issue2_idx_T[6] ? 6'h6 : _issue2_idx_T_120; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_122 = _issue2_idx_T[5] ? 6'h5 : _issue2_idx_T_121; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_123 = _issue2_idx_T[4] ? 6'h4 : _issue2_idx_T_122; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_124 = _issue2_idx_T[3] ? 6'h3 : _issue2_idx_T_123; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_125 = _issue2_idx_T[2] ? 6'h2 : _issue2_idx_T_124; // @[Mux.scala 47:70]
  wire [5:0] _issue2_idx_T_126 = _issue2_idx_T[1] ? 6'h1 : _issue2_idx_T_125; // @[Mux.scala 47:70]
  wire [5:0] issue2_idx = _issue2_idx_T[0] ? 6'h0 : _issue2_idx_T_126; // @[Mux.scala 47:70]
  wire  _issue_num_T = issue1_idx == 6'h3f; // @[reservation_station.scala 87:21]
  wire  _issue_num_T_1 = issue2_idx == 6'h3f; // @[reservation_station.scala 87:42]
  wire  _issue_num_T_2 = issue1_idx == 6'h3f & issue2_idx == 6'h3f; // @[reservation_station.scala 87:29]
  wire  _issue_num_T_4 = issue2_idx != 6'h3f; // @[reservation_station.scala 88:43]
  wire  _issue_num_T_6 = issue1_idx != 6'h3f; // @[reservation_station.scala 88:66]
  wire  _issue_num_T_9 = _issue_num_T & issue2_idx != 6'h3f | issue1_idx != 6'h3f & _issue_num_T_1; // @[reservation_station.scala 88:52]
  wire  _issue_num_T_12 = _issue_num_T_6 & _issue_num_T_4; // @[reservation_station.scala 89:29]
  wire [1:0] _issue_num_T_13 = _issue_num_T_12 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _issue_num_T_14 = _issue_num_T_9 ? 2'h1 : _issue_num_T_13; // @[Mux.scala 101:16]
  wire [1:0] issue_num = _issue_num_T_2 ? 2'h0 : _issue_num_T_14; // @[Mux.scala 101:16]
  wire  _write_num_T = write_idx1 == 6'h3f; // @[reservation_station.scala 98:21]
  wire  _write_num_T_1 = write_idx2 == 6'h3f; // @[reservation_station.scala 98:42]
  wire [31:0] _io_o_issue_packs_0_T_64_pc = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_pc :
    reservation_station_0_io_o_uop_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_64_inst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_inst :
    reservation_station_0_io_o_uop_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_func_code = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_func_code :
    reservation_station_0_io_o_uop_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_branch_predict_pack_valid = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_valid : reservation_station_0_io_o_uop_branch_predict_pack_valid
    ; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_branch_predict_pack_target = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_target :
    reservation_station_0_io_o_uop_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_64_branch_predict_pack_branch_type = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_branch_type :
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_branch_predict_pack_select = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_select :
    reservation_station_0_io_o_uop_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_branch_predict_pack_taken = _issue1_func_code_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_taken : reservation_station_0_io_o_uop_branch_predict_pack_taken
    ; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_phy_dst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_phy_dst :
    reservation_station_0_io_o_uop_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_stale_dst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_stale_dst :
    reservation_station_0_io_o_uop_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_arch_dst = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_arch_dst :
    reservation_station_0_io_o_uop_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_64_inst_type = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_inst_type :
    reservation_station_0_io_o_uop_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_regWen = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_regWen :
    reservation_station_0_io_o_uop_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_src1_valid = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src1_valid :
    reservation_station_0_io_o_uop_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_phy_rs1 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_phy_rs1 :
    reservation_station_0_io_o_uop_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_arch_rs1 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_arch_rs1 :
    reservation_station_0_io_o_uop_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_64_src2_valid = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src2_valid :
    reservation_station_0_io_o_uop_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_phy_rs2 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_phy_rs2 :
    reservation_station_0_io_o_uop_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_arch_rs2 = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_arch_rs2 :
    reservation_station_0_io_o_uop_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_64_rob_idx = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_rob_idx :
    reservation_station_0_io_o_uop_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_imm = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_imm :
    reservation_station_0_io_o_uop_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_src1_value = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src1_value
     : reservation_station_0_io_o_uop_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_64_src2_value = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_src2_value
     : reservation_station_0_io_o_uop_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_64_op1_sel = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_op1_sel :
    reservation_station_0_io_o_uop_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_64_op2_sel = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_op2_sel :
    reservation_station_0_io_o_uop_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_64_alu_sel = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_alu_sel :
    reservation_station_0_io_o_uop_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_64_branch_type = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_branch_type
     : reservation_station_0_io_o_uop_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_64_mem_type = _issue1_func_code_T_63 ? reservation_station_63_io_o_uop_mem_type :
    reservation_station_0_io_o_uop_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_65_pc = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_pc :
    _io_o_issue_packs_0_T_64_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_65_inst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_inst :
    _io_o_issue_packs_0_T_64_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_func_code = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_func_code :
    _io_o_issue_packs_0_T_64_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_branch_predict_pack_valid = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_64_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_branch_predict_pack_target = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_64_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_65_branch_predict_pack_branch_type = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_64_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_branch_predict_pack_select = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_64_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_branch_predict_pack_taken = _issue1_func_code_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_64_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_phy_dst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_64_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_stale_dst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_64_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_arch_dst = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_64_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_65_inst_type = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_64_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_regWen = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_regWen :
    _io_o_issue_packs_0_T_64_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_src1_valid = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_64_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_phy_rs1 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_64_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_arch_rs1 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_64_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_65_src2_valid = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_64_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_phy_rs2 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_64_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_arch_rs2 = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_64_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_65_rob_idx = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_64_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_imm = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_imm :
    _io_o_issue_packs_0_T_64_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_src1_value = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_64_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_65_src2_value = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_64_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_65_op1_sel = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_64_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_65_op2_sel = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_64_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_65_alu_sel = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_64_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_65_branch_type = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_64_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_65_mem_type = _issue1_func_code_T_62 ? reservation_station_62_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_64_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_66_pc = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_pc :
    _io_o_issue_packs_0_T_65_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_66_inst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_inst :
    _io_o_issue_packs_0_T_65_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_func_code = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_func_code :
    _io_o_issue_packs_0_T_65_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_branch_predict_pack_valid = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_65_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_branch_predict_pack_target = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_65_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_66_branch_predict_pack_branch_type = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_65_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_branch_predict_pack_select = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_65_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_branch_predict_pack_taken = _issue1_func_code_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_65_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_phy_dst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_65_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_stale_dst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_65_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_arch_dst = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_65_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_66_inst_type = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_65_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_regWen = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_regWen :
    _io_o_issue_packs_0_T_65_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_src1_valid = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_65_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_phy_rs1 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_65_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_arch_rs1 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_65_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_66_src2_valid = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_65_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_phy_rs2 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_65_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_arch_rs2 = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_65_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_66_rob_idx = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_65_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_imm = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_imm :
    _io_o_issue_packs_0_T_65_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_src1_value = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_65_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_66_src2_value = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_65_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_66_op1_sel = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_65_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_66_op2_sel = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_65_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_66_alu_sel = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_65_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_66_branch_type = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_65_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_66_mem_type = _issue1_func_code_T_61 ? reservation_station_61_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_65_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_67_pc = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_pc :
    _io_o_issue_packs_0_T_66_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_67_inst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_inst :
    _io_o_issue_packs_0_T_66_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_func_code = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_func_code :
    _io_o_issue_packs_0_T_66_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_branch_predict_pack_valid = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_66_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_branch_predict_pack_target = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_66_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_67_branch_predict_pack_branch_type = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_66_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_branch_predict_pack_select = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_66_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_branch_predict_pack_taken = _issue1_func_code_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_66_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_phy_dst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_66_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_stale_dst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_66_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_arch_dst = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_66_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_67_inst_type = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_66_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_regWen = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_regWen :
    _io_o_issue_packs_0_T_66_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_src1_valid = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_66_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_phy_rs1 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_66_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_arch_rs1 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_66_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_67_src2_valid = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_66_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_phy_rs2 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_66_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_arch_rs2 = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_66_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_67_rob_idx = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_66_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_imm = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_imm :
    _io_o_issue_packs_0_T_66_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_src1_value = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_66_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_67_src2_value = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_66_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_67_op1_sel = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_66_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_67_op2_sel = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_66_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_67_alu_sel = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_66_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_67_branch_type = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_66_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_67_mem_type = _issue1_func_code_T_60 ? reservation_station_60_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_66_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_68_pc = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_pc :
    _io_o_issue_packs_0_T_67_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_68_inst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_inst :
    _io_o_issue_packs_0_T_67_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_func_code = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_func_code :
    _io_o_issue_packs_0_T_67_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_branch_predict_pack_valid = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_67_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_branch_predict_pack_target = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_67_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_68_branch_predict_pack_branch_type = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_67_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_branch_predict_pack_select = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_67_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_branch_predict_pack_taken = _issue1_func_code_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_67_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_phy_dst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_67_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_stale_dst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_67_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_arch_dst = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_67_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_68_inst_type = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_67_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_regWen = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_regWen :
    _io_o_issue_packs_0_T_67_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_src1_valid = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_67_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_phy_rs1 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_67_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_arch_rs1 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_67_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_68_src2_valid = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_67_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_phy_rs2 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_67_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_arch_rs2 = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_67_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_68_rob_idx = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_67_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_imm = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_imm :
    _io_o_issue_packs_0_T_67_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_src1_value = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_67_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_68_src2_value = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_67_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_68_op1_sel = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_67_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_68_op2_sel = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_67_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_68_alu_sel = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_67_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_68_branch_type = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_67_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_68_mem_type = _issue1_func_code_T_59 ? reservation_station_59_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_67_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_69_pc = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_pc :
    _io_o_issue_packs_0_T_68_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_69_inst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_inst :
    _io_o_issue_packs_0_T_68_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_func_code = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_func_code :
    _io_o_issue_packs_0_T_68_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_branch_predict_pack_valid = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_68_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_branch_predict_pack_target = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_68_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_69_branch_predict_pack_branch_type = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_68_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_branch_predict_pack_select = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_68_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_branch_predict_pack_taken = _issue1_func_code_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_68_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_phy_dst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_68_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_stale_dst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_68_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_arch_dst = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_68_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_69_inst_type = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_68_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_regWen = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_regWen :
    _io_o_issue_packs_0_T_68_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_src1_valid = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_68_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_phy_rs1 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_68_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_arch_rs1 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_68_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_69_src2_valid = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_68_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_phy_rs2 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_68_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_arch_rs2 = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_68_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_69_rob_idx = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_68_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_imm = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_imm :
    _io_o_issue_packs_0_T_68_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_src1_value = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_68_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_69_src2_value = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_68_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_69_op1_sel = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_68_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_69_op2_sel = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_68_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_69_alu_sel = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_68_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_69_branch_type = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_68_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_69_mem_type = _issue1_func_code_T_58 ? reservation_station_58_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_68_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_70_pc = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_pc :
    _io_o_issue_packs_0_T_69_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_70_inst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_inst :
    _io_o_issue_packs_0_T_69_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_func_code = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_func_code :
    _io_o_issue_packs_0_T_69_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_branch_predict_pack_valid = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_69_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_branch_predict_pack_target = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_69_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_70_branch_predict_pack_branch_type = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_69_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_branch_predict_pack_select = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_69_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_branch_predict_pack_taken = _issue1_func_code_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_69_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_phy_dst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_69_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_stale_dst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_69_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_arch_dst = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_69_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_70_inst_type = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_69_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_regWen = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_regWen :
    _io_o_issue_packs_0_T_69_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_src1_valid = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_69_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_phy_rs1 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_69_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_arch_rs1 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_69_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_70_src2_valid = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_69_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_phy_rs2 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_69_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_arch_rs2 = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_69_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_70_rob_idx = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_69_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_imm = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_imm :
    _io_o_issue_packs_0_T_69_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_src1_value = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_69_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_70_src2_value = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_69_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_70_op1_sel = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_69_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_70_op2_sel = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_69_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_70_alu_sel = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_69_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_70_branch_type = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_69_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_70_mem_type = _issue1_func_code_T_57 ? reservation_station_57_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_69_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_71_pc = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_pc :
    _io_o_issue_packs_0_T_70_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_71_inst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_inst :
    _io_o_issue_packs_0_T_70_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_func_code = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_func_code :
    _io_o_issue_packs_0_T_70_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_branch_predict_pack_valid = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_70_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_branch_predict_pack_target = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_70_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_71_branch_predict_pack_branch_type = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_70_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_branch_predict_pack_select = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_70_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_branch_predict_pack_taken = _issue1_func_code_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_70_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_phy_dst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_70_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_stale_dst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_70_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_arch_dst = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_70_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_71_inst_type = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_70_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_regWen = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_regWen :
    _io_o_issue_packs_0_T_70_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_src1_valid = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_70_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_phy_rs1 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_70_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_arch_rs1 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_70_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_71_src2_valid = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_70_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_phy_rs2 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_70_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_arch_rs2 = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_70_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_71_rob_idx = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_70_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_imm = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_imm :
    _io_o_issue_packs_0_T_70_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_src1_value = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_70_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_71_src2_value = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_70_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_71_op1_sel = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_70_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_71_op2_sel = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_70_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_71_alu_sel = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_70_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_71_branch_type = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_70_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_71_mem_type = _issue1_func_code_T_56 ? reservation_station_56_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_70_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_72_pc = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_pc :
    _io_o_issue_packs_0_T_71_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_72_inst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_inst :
    _io_o_issue_packs_0_T_71_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_func_code = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_func_code :
    _io_o_issue_packs_0_T_71_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_branch_predict_pack_valid = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_71_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_branch_predict_pack_target = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_71_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_72_branch_predict_pack_branch_type = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_71_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_branch_predict_pack_select = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_71_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_branch_predict_pack_taken = _issue1_func_code_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_71_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_phy_dst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_71_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_stale_dst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_71_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_arch_dst = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_71_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_72_inst_type = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_71_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_regWen = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_regWen :
    _io_o_issue_packs_0_T_71_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_src1_valid = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_71_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_phy_rs1 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_71_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_arch_rs1 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_71_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_72_src2_valid = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_71_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_phy_rs2 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_71_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_arch_rs2 = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_71_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_72_rob_idx = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_71_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_imm = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_imm :
    _io_o_issue_packs_0_T_71_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_src1_value = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_71_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_72_src2_value = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_71_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_72_op1_sel = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_71_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_72_op2_sel = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_71_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_72_alu_sel = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_71_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_72_branch_type = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_71_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_72_mem_type = _issue1_func_code_T_55 ? reservation_station_55_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_71_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_73_pc = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_pc :
    _io_o_issue_packs_0_T_72_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_73_inst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_inst :
    _io_o_issue_packs_0_T_72_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_func_code = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_func_code :
    _io_o_issue_packs_0_T_72_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_branch_predict_pack_valid = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_72_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_branch_predict_pack_target = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_72_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_73_branch_predict_pack_branch_type = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_72_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_branch_predict_pack_select = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_72_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_branch_predict_pack_taken = _issue1_func_code_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_72_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_phy_dst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_72_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_stale_dst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_72_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_arch_dst = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_72_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_73_inst_type = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_72_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_regWen = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_regWen :
    _io_o_issue_packs_0_T_72_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_src1_valid = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_72_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_phy_rs1 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_72_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_arch_rs1 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_72_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_73_src2_valid = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_72_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_phy_rs2 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_72_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_arch_rs2 = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_72_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_73_rob_idx = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_72_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_imm = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_imm :
    _io_o_issue_packs_0_T_72_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_src1_value = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_72_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_73_src2_value = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_72_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_73_op1_sel = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_72_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_73_op2_sel = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_72_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_73_alu_sel = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_72_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_73_branch_type = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_72_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_73_mem_type = _issue1_func_code_T_54 ? reservation_station_54_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_72_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_74_pc = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_pc :
    _io_o_issue_packs_0_T_73_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_74_inst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_inst :
    _io_o_issue_packs_0_T_73_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_func_code = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_func_code :
    _io_o_issue_packs_0_T_73_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_branch_predict_pack_valid = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_73_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_branch_predict_pack_target = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_73_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_74_branch_predict_pack_branch_type = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_73_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_branch_predict_pack_select = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_73_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_branch_predict_pack_taken = _issue1_func_code_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_73_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_phy_dst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_73_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_stale_dst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_73_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_arch_dst = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_73_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_74_inst_type = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_73_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_regWen = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_regWen :
    _io_o_issue_packs_0_T_73_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_src1_valid = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_73_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_phy_rs1 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_73_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_arch_rs1 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_73_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_74_src2_valid = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_73_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_phy_rs2 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_73_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_arch_rs2 = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_73_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_74_rob_idx = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_73_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_imm = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_imm :
    _io_o_issue_packs_0_T_73_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_src1_value = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_73_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_74_src2_value = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_73_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_74_op1_sel = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_73_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_74_op2_sel = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_73_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_74_alu_sel = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_73_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_74_branch_type = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_73_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_74_mem_type = _issue1_func_code_T_53 ? reservation_station_53_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_73_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_75_pc = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_pc :
    _io_o_issue_packs_0_T_74_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_75_inst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_inst :
    _io_o_issue_packs_0_T_74_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_func_code = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_func_code :
    _io_o_issue_packs_0_T_74_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_branch_predict_pack_valid = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_74_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_branch_predict_pack_target = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_74_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_75_branch_predict_pack_branch_type = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_74_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_branch_predict_pack_select = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_74_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_branch_predict_pack_taken = _issue1_func_code_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_74_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_phy_dst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_74_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_stale_dst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_74_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_arch_dst = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_74_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_75_inst_type = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_74_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_regWen = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_regWen :
    _io_o_issue_packs_0_T_74_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_src1_valid = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_74_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_phy_rs1 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_74_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_arch_rs1 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_74_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_75_src2_valid = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_74_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_phy_rs2 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_74_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_arch_rs2 = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_74_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_75_rob_idx = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_74_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_imm = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_imm :
    _io_o_issue_packs_0_T_74_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_src1_value = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_74_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_75_src2_value = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_74_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_75_op1_sel = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_74_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_75_op2_sel = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_74_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_75_alu_sel = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_74_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_75_branch_type = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_74_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_75_mem_type = _issue1_func_code_T_52 ? reservation_station_52_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_74_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_76_pc = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_pc :
    _io_o_issue_packs_0_T_75_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_76_inst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_inst :
    _io_o_issue_packs_0_T_75_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_func_code = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_func_code :
    _io_o_issue_packs_0_T_75_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_branch_predict_pack_valid = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_75_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_branch_predict_pack_target = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_75_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_76_branch_predict_pack_branch_type = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_75_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_branch_predict_pack_select = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_75_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_branch_predict_pack_taken = _issue1_func_code_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_75_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_phy_dst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_75_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_stale_dst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_75_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_arch_dst = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_75_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_76_inst_type = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_75_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_regWen = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_regWen :
    _io_o_issue_packs_0_T_75_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_src1_valid = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_75_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_phy_rs1 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_75_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_arch_rs1 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_75_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_76_src2_valid = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_75_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_phy_rs2 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_75_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_arch_rs2 = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_75_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_76_rob_idx = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_75_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_imm = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_imm :
    _io_o_issue_packs_0_T_75_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_src1_value = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_75_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_76_src2_value = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_75_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_76_op1_sel = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_75_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_76_op2_sel = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_75_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_76_alu_sel = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_75_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_76_branch_type = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_75_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_76_mem_type = _issue1_func_code_T_51 ? reservation_station_51_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_75_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_77_pc = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_pc :
    _io_o_issue_packs_0_T_76_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_77_inst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_inst :
    _io_o_issue_packs_0_T_76_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_func_code = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_func_code :
    _io_o_issue_packs_0_T_76_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_branch_predict_pack_valid = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_76_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_branch_predict_pack_target = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_76_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_77_branch_predict_pack_branch_type = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_76_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_branch_predict_pack_select = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_76_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_branch_predict_pack_taken = _issue1_func_code_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_76_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_phy_dst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_76_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_stale_dst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_76_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_arch_dst = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_76_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_77_inst_type = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_76_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_regWen = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_regWen :
    _io_o_issue_packs_0_T_76_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_src1_valid = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_76_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_phy_rs1 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_76_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_arch_rs1 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_76_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_77_src2_valid = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_76_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_phy_rs2 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_76_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_arch_rs2 = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_76_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_77_rob_idx = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_76_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_imm = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_imm :
    _io_o_issue_packs_0_T_76_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_src1_value = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_76_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_77_src2_value = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_76_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_77_op1_sel = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_76_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_77_op2_sel = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_76_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_77_alu_sel = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_76_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_77_branch_type = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_76_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_77_mem_type = _issue1_func_code_T_50 ? reservation_station_50_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_76_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_78_pc = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_pc :
    _io_o_issue_packs_0_T_77_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_78_inst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_inst :
    _io_o_issue_packs_0_T_77_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_func_code = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_func_code :
    _io_o_issue_packs_0_T_77_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_branch_predict_pack_valid = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_77_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_branch_predict_pack_target = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_77_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_78_branch_predict_pack_branch_type = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_77_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_branch_predict_pack_select = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_77_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_branch_predict_pack_taken = _issue1_func_code_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_77_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_phy_dst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_77_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_stale_dst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_77_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_arch_dst = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_77_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_78_inst_type = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_77_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_regWen = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_regWen :
    _io_o_issue_packs_0_T_77_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_src1_valid = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_77_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_phy_rs1 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_77_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_arch_rs1 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_77_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_78_src2_valid = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_77_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_phy_rs2 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_77_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_arch_rs2 = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_77_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_78_rob_idx = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_77_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_imm = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_imm :
    _io_o_issue_packs_0_T_77_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_src1_value = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_77_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_78_src2_value = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_77_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_78_op1_sel = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_77_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_78_op2_sel = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_77_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_78_alu_sel = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_77_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_78_branch_type = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_77_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_78_mem_type = _issue1_func_code_T_49 ? reservation_station_49_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_77_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_79_pc = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_pc :
    _io_o_issue_packs_0_T_78_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_79_inst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_inst :
    _io_o_issue_packs_0_T_78_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_func_code = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_func_code :
    _io_o_issue_packs_0_T_78_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_branch_predict_pack_valid = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_78_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_branch_predict_pack_target = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_78_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_79_branch_predict_pack_branch_type = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_78_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_branch_predict_pack_select = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_78_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_branch_predict_pack_taken = _issue1_func_code_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_78_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_phy_dst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_78_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_stale_dst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_78_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_arch_dst = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_78_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_79_inst_type = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_78_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_regWen = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_regWen :
    _io_o_issue_packs_0_T_78_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_src1_valid = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_78_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_phy_rs1 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_78_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_arch_rs1 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_78_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_79_src2_valid = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_78_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_phy_rs2 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_78_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_arch_rs2 = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_78_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_79_rob_idx = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_78_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_imm = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_imm :
    _io_o_issue_packs_0_T_78_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_src1_value = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_78_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_79_src2_value = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_78_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_79_op1_sel = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_78_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_79_op2_sel = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_78_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_79_alu_sel = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_78_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_79_branch_type = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_78_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_79_mem_type = _issue1_func_code_T_48 ? reservation_station_48_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_78_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_80_pc = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_pc :
    _io_o_issue_packs_0_T_79_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_80_inst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_inst :
    _io_o_issue_packs_0_T_79_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_func_code = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_func_code :
    _io_o_issue_packs_0_T_79_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_branch_predict_pack_valid = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_79_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_branch_predict_pack_target = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_79_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_80_branch_predict_pack_branch_type = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_79_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_branch_predict_pack_select = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_79_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_branch_predict_pack_taken = _issue1_func_code_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_79_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_phy_dst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_79_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_stale_dst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_79_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_arch_dst = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_79_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_80_inst_type = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_79_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_regWen = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_regWen :
    _io_o_issue_packs_0_T_79_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_src1_valid = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_79_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_phy_rs1 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_79_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_arch_rs1 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_79_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_80_src2_valid = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_79_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_phy_rs2 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_79_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_arch_rs2 = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_79_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_80_rob_idx = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_79_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_imm = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_imm :
    _io_o_issue_packs_0_T_79_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_src1_value = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_79_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_80_src2_value = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_79_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_80_op1_sel = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_79_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_80_op2_sel = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_79_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_80_alu_sel = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_79_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_80_branch_type = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_79_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_80_mem_type = _issue1_func_code_T_47 ? reservation_station_47_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_79_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_81_pc = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_pc :
    _io_o_issue_packs_0_T_80_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_81_inst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_inst :
    _io_o_issue_packs_0_T_80_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_func_code = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_func_code :
    _io_o_issue_packs_0_T_80_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_branch_predict_pack_valid = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_80_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_branch_predict_pack_target = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_80_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_81_branch_predict_pack_branch_type = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_80_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_branch_predict_pack_select = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_80_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_branch_predict_pack_taken = _issue1_func_code_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_80_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_phy_dst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_80_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_stale_dst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_80_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_arch_dst = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_80_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_81_inst_type = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_80_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_regWen = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_regWen :
    _io_o_issue_packs_0_T_80_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_src1_valid = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_80_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_phy_rs1 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_80_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_arch_rs1 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_80_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_81_src2_valid = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_80_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_phy_rs2 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_80_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_arch_rs2 = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_80_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_81_rob_idx = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_80_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_imm = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_imm :
    _io_o_issue_packs_0_T_80_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_src1_value = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_80_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_81_src2_value = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_80_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_81_op1_sel = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_80_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_81_op2_sel = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_80_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_81_alu_sel = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_80_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_81_branch_type = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_80_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_81_mem_type = _issue1_func_code_T_46 ? reservation_station_46_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_80_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_82_pc = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_pc :
    _io_o_issue_packs_0_T_81_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_82_inst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_inst :
    _io_o_issue_packs_0_T_81_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_func_code = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_func_code :
    _io_o_issue_packs_0_T_81_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_branch_predict_pack_valid = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_81_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_branch_predict_pack_target = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_81_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_82_branch_predict_pack_branch_type = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_81_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_branch_predict_pack_select = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_81_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_branch_predict_pack_taken = _issue1_func_code_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_81_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_phy_dst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_81_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_stale_dst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_81_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_arch_dst = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_81_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_82_inst_type = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_81_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_regWen = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_regWen :
    _io_o_issue_packs_0_T_81_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_src1_valid = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_81_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_phy_rs1 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_81_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_arch_rs1 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_81_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_82_src2_valid = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_81_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_phy_rs2 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_81_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_arch_rs2 = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_81_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_82_rob_idx = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_81_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_imm = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_imm :
    _io_o_issue_packs_0_T_81_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_src1_value = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_81_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_82_src2_value = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_81_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_82_op1_sel = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_81_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_82_op2_sel = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_81_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_82_alu_sel = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_81_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_82_branch_type = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_81_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_82_mem_type = _issue1_func_code_T_45 ? reservation_station_45_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_81_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_83_pc = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_pc :
    _io_o_issue_packs_0_T_82_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_83_inst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_inst :
    _io_o_issue_packs_0_T_82_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_func_code = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_func_code :
    _io_o_issue_packs_0_T_82_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_branch_predict_pack_valid = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_82_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_branch_predict_pack_target = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_82_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_83_branch_predict_pack_branch_type = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_82_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_branch_predict_pack_select = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_82_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_branch_predict_pack_taken = _issue1_func_code_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_82_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_phy_dst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_82_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_stale_dst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_82_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_arch_dst = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_82_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_83_inst_type = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_82_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_regWen = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_regWen :
    _io_o_issue_packs_0_T_82_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_src1_valid = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_82_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_phy_rs1 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_82_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_arch_rs1 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_82_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_83_src2_valid = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_82_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_phy_rs2 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_82_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_arch_rs2 = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_82_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_83_rob_idx = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_82_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_imm = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_imm :
    _io_o_issue_packs_0_T_82_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_src1_value = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_82_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_83_src2_value = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_82_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_83_op1_sel = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_82_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_83_op2_sel = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_82_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_83_alu_sel = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_82_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_83_branch_type = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_82_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_83_mem_type = _issue1_func_code_T_44 ? reservation_station_44_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_82_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_84_pc = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_pc :
    _io_o_issue_packs_0_T_83_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_84_inst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_inst :
    _io_o_issue_packs_0_T_83_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_func_code = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_func_code :
    _io_o_issue_packs_0_T_83_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_branch_predict_pack_valid = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_83_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_branch_predict_pack_target = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_83_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_84_branch_predict_pack_branch_type = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_83_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_branch_predict_pack_select = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_83_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_branch_predict_pack_taken = _issue1_func_code_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_83_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_phy_dst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_83_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_stale_dst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_83_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_arch_dst = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_83_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_84_inst_type = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_83_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_regWen = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_regWen :
    _io_o_issue_packs_0_T_83_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_src1_valid = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_83_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_phy_rs1 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_83_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_arch_rs1 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_83_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_84_src2_valid = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_83_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_phy_rs2 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_83_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_arch_rs2 = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_83_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_84_rob_idx = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_83_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_imm = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_imm :
    _io_o_issue_packs_0_T_83_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_src1_value = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_83_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_84_src2_value = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_83_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_84_op1_sel = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_83_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_84_op2_sel = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_83_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_84_alu_sel = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_83_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_84_branch_type = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_83_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_84_mem_type = _issue1_func_code_T_43 ? reservation_station_43_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_83_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_85_pc = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_pc :
    _io_o_issue_packs_0_T_84_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_85_inst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_inst :
    _io_o_issue_packs_0_T_84_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_func_code = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_func_code :
    _io_o_issue_packs_0_T_84_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_branch_predict_pack_valid = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_84_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_branch_predict_pack_target = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_84_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_85_branch_predict_pack_branch_type = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_84_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_branch_predict_pack_select = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_84_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_branch_predict_pack_taken = _issue1_func_code_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_84_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_phy_dst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_84_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_stale_dst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_84_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_arch_dst = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_84_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_85_inst_type = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_84_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_regWen = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_regWen :
    _io_o_issue_packs_0_T_84_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_src1_valid = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_84_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_phy_rs1 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_84_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_arch_rs1 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_84_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_85_src2_valid = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_84_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_phy_rs2 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_84_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_arch_rs2 = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_84_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_85_rob_idx = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_84_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_imm = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_imm :
    _io_o_issue_packs_0_T_84_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_src1_value = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_84_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_85_src2_value = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_84_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_85_op1_sel = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_84_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_85_op2_sel = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_84_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_85_alu_sel = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_84_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_85_branch_type = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_84_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_85_mem_type = _issue1_func_code_T_42 ? reservation_station_42_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_84_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_86_pc = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_pc :
    _io_o_issue_packs_0_T_85_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_86_inst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_inst :
    _io_o_issue_packs_0_T_85_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_func_code = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_func_code :
    _io_o_issue_packs_0_T_85_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_branch_predict_pack_valid = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_85_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_branch_predict_pack_target = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_85_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_86_branch_predict_pack_branch_type = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_85_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_branch_predict_pack_select = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_85_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_branch_predict_pack_taken = _issue1_func_code_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_85_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_phy_dst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_85_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_stale_dst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_85_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_arch_dst = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_85_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_86_inst_type = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_85_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_regWen = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_regWen :
    _io_o_issue_packs_0_T_85_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_src1_valid = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_85_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_phy_rs1 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_85_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_arch_rs1 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_85_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_86_src2_valid = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_85_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_phy_rs2 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_85_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_arch_rs2 = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_85_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_86_rob_idx = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_85_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_imm = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_imm :
    _io_o_issue_packs_0_T_85_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_src1_value = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_85_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_86_src2_value = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_85_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_86_op1_sel = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_85_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_86_op2_sel = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_85_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_86_alu_sel = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_85_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_86_branch_type = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_85_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_86_mem_type = _issue1_func_code_T_41 ? reservation_station_41_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_85_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_87_pc = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_pc :
    _io_o_issue_packs_0_T_86_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_87_inst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_inst :
    _io_o_issue_packs_0_T_86_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_func_code = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_func_code :
    _io_o_issue_packs_0_T_86_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_branch_predict_pack_valid = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_86_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_branch_predict_pack_target = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_86_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_87_branch_predict_pack_branch_type = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_86_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_branch_predict_pack_select = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_86_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_branch_predict_pack_taken = _issue1_func_code_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_86_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_phy_dst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_86_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_stale_dst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_86_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_arch_dst = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_86_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_87_inst_type = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_86_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_regWen = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_regWen :
    _io_o_issue_packs_0_T_86_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_src1_valid = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_86_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_phy_rs1 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_86_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_arch_rs1 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_86_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_87_src2_valid = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_86_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_phy_rs2 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_86_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_arch_rs2 = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_86_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_87_rob_idx = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_86_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_imm = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_imm :
    _io_o_issue_packs_0_T_86_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_src1_value = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_86_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_87_src2_value = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_86_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_87_op1_sel = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_86_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_87_op2_sel = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_86_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_87_alu_sel = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_86_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_87_branch_type = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_86_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_87_mem_type = _issue1_func_code_T_40 ? reservation_station_40_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_86_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_88_pc = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_pc :
    _io_o_issue_packs_0_T_87_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_88_inst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_inst :
    _io_o_issue_packs_0_T_87_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_func_code = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_func_code :
    _io_o_issue_packs_0_T_87_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_branch_predict_pack_valid = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_87_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_branch_predict_pack_target = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_87_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_88_branch_predict_pack_branch_type = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_87_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_branch_predict_pack_select = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_87_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_branch_predict_pack_taken = _issue1_func_code_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_87_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_phy_dst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_87_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_stale_dst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_87_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_arch_dst = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_87_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_88_inst_type = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_87_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_regWen = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_regWen :
    _io_o_issue_packs_0_T_87_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_src1_valid = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_87_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_phy_rs1 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_87_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_arch_rs1 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_87_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_88_src2_valid = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_87_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_phy_rs2 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_87_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_arch_rs2 = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_87_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_88_rob_idx = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_87_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_imm = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_imm :
    _io_o_issue_packs_0_T_87_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_src1_value = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_87_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_88_src2_value = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_87_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_88_op1_sel = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_87_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_88_op2_sel = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_87_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_88_alu_sel = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_87_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_88_branch_type = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_87_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_88_mem_type = _issue1_func_code_T_39 ? reservation_station_39_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_87_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_89_pc = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_pc :
    _io_o_issue_packs_0_T_88_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_89_inst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_inst :
    _io_o_issue_packs_0_T_88_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_func_code = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_func_code :
    _io_o_issue_packs_0_T_88_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_branch_predict_pack_valid = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_88_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_branch_predict_pack_target = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_88_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_89_branch_predict_pack_branch_type = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_88_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_branch_predict_pack_select = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_88_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_branch_predict_pack_taken = _issue1_func_code_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_88_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_phy_dst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_88_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_stale_dst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_88_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_arch_dst = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_88_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_89_inst_type = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_88_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_regWen = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_regWen :
    _io_o_issue_packs_0_T_88_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_src1_valid = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_88_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_phy_rs1 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_88_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_arch_rs1 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_88_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_89_src2_valid = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_88_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_phy_rs2 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_88_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_arch_rs2 = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_88_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_89_rob_idx = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_88_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_imm = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_imm :
    _io_o_issue_packs_0_T_88_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_src1_value = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_88_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_89_src2_value = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_88_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_89_op1_sel = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_88_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_89_op2_sel = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_88_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_89_alu_sel = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_88_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_89_branch_type = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_88_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_89_mem_type = _issue1_func_code_T_38 ? reservation_station_38_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_88_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_90_pc = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_pc :
    _io_o_issue_packs_0_T_89_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_90_inst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_inst :
    _io_o_issue_packs_0_T_89_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_func_code = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_func_code :
    _io_o_issue_packs_0_T_89_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_branch_predict_pack_valid = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_89_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_branch_predict_pack_target = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_89_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_90_branch_predict_pack_branch_type = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_89_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_branch_predict_pack_select = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_89_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_branch_predict_pack_taken = _issue1_func_code_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_89_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_phy_dst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_89_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_stale_dst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_89_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_arch_dst = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_89_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_90_inst_type = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_89_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_regWen = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_regWen :
    _io_o_issue_packs_0_T_89_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_src1_valid = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_89_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_phy_rs1 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_89_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_arch_rs1 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_89_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_90_src2_valid = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_89_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_phy_rs2 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_89_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_arch_rs2 = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_89_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_90_rob_idx = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_89_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_imm = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_imm :
    _io_o_issue_packs_0_T_89_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_src1_value = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_89_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_90_src2_value = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_89_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_90_op1_sel = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_89_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_90_op2_sel = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_89_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_90_alu_sel = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_89_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_90_branch_type = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_89_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_90_mem_type = _issue1_func_code_T_37 ? reservation_station_37_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_89_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_91_pc = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_pc :
    _io_o_issue_packs_0_T_90_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_91_inst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_inst :
    _io_o_issue_packs_0_T_90_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_func_code = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_func_code :
    _io_o_issue_packs_0_T_90_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_branch_predict_pack_valid = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_90_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_branch_predict_pack_target = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_90_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_91_branch_predict_pack_branch_type = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_90_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_branch_predict_pack_select = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_90_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_branch_predict_pack_taken = _issue1_func_code_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_90_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_phy_dst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_90_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_stale_dst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_90_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_arch_dst = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_90_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_91_inst_type = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_90_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_regWen = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_regWen :
    _io_o_issue_packs_0_T_90_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_src1_valid = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_90_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_phy_rs1 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_90_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_arch_rs1 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_90_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_91_src2_valid = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_90_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_phy_rs2 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_90_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_arch_rs2 = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_90_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_91_rob_idx = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_90_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_imm = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_imm :
    _io_o_issue_packs_0_T_90_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_src1_value = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_90_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_91_src2_value = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_90_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_91_op1_sel = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_90_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_91_op2_sel = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_90_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_91_alu_sel = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_90_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_91_branch_type = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_90_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_91_mem_type = _issue1_func_code_T_36 ? reservation_station_36_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_90_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_92_pc = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_pc :
    _io_o_issue_packs_0_T_91_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_92_inst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_inst :
    _io_o_issue_packs_0_T_91_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_func_code = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_func_code :
    _io_o_issue_packs_0_T_91_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_branch_predict_pack_valid = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_91_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_branch_predict_pack_target = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_91_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_92_branch_predict_pack_branch_type = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_91_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_branch_predict_pack_select = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_91_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_branch_predict_pack_taken = _issue1_func_code_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_91_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_phy_dst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_91_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_stale_dst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_91_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_arch_dst = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_91_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_92_inst_type = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_91_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_regWen = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_regWen :
    _io_o_issue_packs_0_T_91_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_src1_valid = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_91_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_phy_rs1 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_91_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_arch_rs1 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_91_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_92_src2_valid = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_91_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_phy_rs2 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_91_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_arch_rs2 = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_91_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_92_rob_idx = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_91_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_imm = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_imm :
    _io_o_issue_packs_0_T_91_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_src1_value = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_91_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_92_src2_value = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_91_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_92_op1_sel = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_91_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_92_op2_sel = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_91_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_92_alu_sel = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_91_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_92_branch_type = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_91_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_92_mem_type = _issue1_func_code_T_35 ? reservation_station_35_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_91_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_93_pc = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_pc :
    _io_o_issue_packs_0_T_92_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_93_inst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_inst :
    _io_o_issue_packs_0_T_92_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_func_code = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_func_code :
    _io_o_issue_packs_0_T_92_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_branch_predict_pack_valid = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_92_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_branch_predict_pack_target = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_92_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_93_branch_predict_pack_branch_type = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_92_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_branch_predict_pack_select = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_92_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_branch_predict_pack_taken = _issue1_func_code_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_92_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_phy_dst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_92_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_stale_dst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_92_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_arch_dst = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_92_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_93_inst_type = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_92_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_regWen = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_regWen :
    _io_o_issue_packs_0_T_92_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_src1_valid = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_92_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_phy_rs1 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_92_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_arch_rs1 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_92_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_93_src2_valid = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_92_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_phy_rs2 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_92_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_arch_rs2 = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_92_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_93_rob_idx = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_92_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_imm = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_imm :
    _io_o_issue_packs_0_T_92_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_src1_value = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_92_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_93_src2_value = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_92_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_93_op1_sel = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_92_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_93_op2_sel = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_92_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_93_alu_sel = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_92_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_93_branch_type = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_92_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_93_mem_type = _issue1_func_code_T_34 ? reservation_station_34_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_92_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_94_pc = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_pc :
    _io_o_issue_packs_0_T_93_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_94_inst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_inst :
    _io_o_issue_packs_0_T_93_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_func_code = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_func_code :
    _io_o_issue_packs_0_T_93_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_branch_predict_pack_valid = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_93_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_branch_predict_pack_target = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_93_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_94_branch_predict_pack_branch_type = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_93_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_branch_predict_pack_select = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_93_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_branch_predict_pack_taken = _issue1_func_code_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_93_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_phy_dst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_93_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_stale_dst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_93_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_arch_dst = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_93_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_94_inst_type = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_93_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_regWen = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_regWen :
    _io_o_issue_packs_0_T_93_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_src1_valid = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_93_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_phy_rs1 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_93_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_arch_rs1 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_93_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_94_src2_valid = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_93_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_phy_rs2 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_93_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_arch_rs2 = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_93_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_94_rob_idx = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_93_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_imm = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_imm :
    _io_o_issue_packs_0_T_93_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_src1_value = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_93_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_94_src2_value = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_93_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_94_op1_sel = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_93_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_94_op2_sel = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_93_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_94_alu_sel = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_93_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_94_branch_type = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_93_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_94_mem_type = _issue1_func_code_T_33 ? reservation_station_33_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_93_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_95_pc = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_pc :
    _io_o_issue_packs_0_T_94_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_95_inst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_inst :
    _io_o_issue_packs_0_T_94_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_func_code = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_func_code :
    _io_o_issue_packs_0_T_94_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_branch_predict_pack_valid = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_94_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_branch_predict_pack_target = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_94_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_95_branch_predict_pack_branch_type = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_94_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_branch_predict_pack_select = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_94_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_branch_predict_pack_taken = _issue1_func_code_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_94_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_phy_dst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_94_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_stale_dst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_94_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_arch_dst = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_94_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_95_inst_type = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_94_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_regWen = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_regWen :
    _io_o_issue_packs_0_T_94_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_src1_valid = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_94_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_phy_rs1 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_94_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_arch_rs1 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_94_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_95_src2_valid = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_94_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_phy_rs2 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_94_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_arch_rs2 = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_94_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_95_rob_idx = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_94_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_imm = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_imm :
    _io_o_issue_packs_0_T_94_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_src1_value = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_94_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_95_src2_value = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_94_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_95_op1_sel = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_94_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_95_op2_sel = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_94_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_95_alu_sel = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_94_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_95_branch_type = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_94_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_95_mem_type = _issue1_func_code_T_32 ? reservation_station_32_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_94_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_96_pc = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_pc :
    _io_o_issue_packs_0_T_95_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_96_inst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_inst :
    _io_o_issue_packs_0_T_95_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_func_code = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_func_code :
    _io_o_issue_packs_0_T_95_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_branch_predict_pack_valid = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_95_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_branch_predict_pack_target = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_95_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_96_branch_predict_pack_branch_type = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_95_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_branch_predict_pack_select = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_95_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_branch_predict_pack_taken = _issue1_func_code_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_95_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_phy_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_95_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_stale_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_95_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_arch_dst = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_95_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_96_inst_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_95_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_regWen = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_regWen :
    _io_o_issue_packs_0_T_95_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_src1_valid = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_95_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_phy_rs1 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_95_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_arch_rs1 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_95_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_96_src2_valid = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_95_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_phy_rs2 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_95_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_arch_rs2 = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_95_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_96_rob_idx = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_95_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_imm = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_imm :
    _io_o_issue_packs_0_T_95_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_src1_value = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_95_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_96_src2_value = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_95_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_96_op1_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_95_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_96_op2_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_95_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_96_alu_sel = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_95_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_96_branch_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_95_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_96_mem_type = _issue1_func_code_T_31 ? reservation_station_31_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_95_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_97_pc = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_pc :
    _io_o_issue_packs_0_T_96_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_97_inst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_inst :
    _io_o_issue_packs_0_T_96_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_func_code = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_func_code :
    _io_o_issue_packs_0_T_96_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_branch_predict_pack_valid = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_96_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_branch_predict_pack_target = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_96_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_97_branch_predict_pack_branch_type = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_96_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_branch_predict_pack_select = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_96_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_branch_predict_pack_taken = _issue1_func_code_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_96_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_phy_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_96_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_stale_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_96_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_arch_dst = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_96_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_97_inst_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_96_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_regWen = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_regWen :
    _io_o_issue_packs_0_T_96_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_src1_valid = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_96_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_phy_rs1 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_96_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_arch_rs1 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_96_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_97_src2_valid = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_96_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_phy_rs2 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_96_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_arch_rs2 = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_96_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_97_rob_idx = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_96_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_imm = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_imm :
    _io_o_issue_packs_0_T_96_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_src1_value = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_96_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_97_src2_value = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_96_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_97_op1_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_96_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_97_op2_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_96_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_97_alu_sel = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_96_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_97_branch_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_96_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_97_mem_type = _issue1_func_code_T_30 ? reservation_station_30_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_96_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_98_pc = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_pc :
    _io_o_issue_packs_0_T_97_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_98_inst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_inst :
    _io_o_issue_packs_0_T_97_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_func_code = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_func_code :
    _io_o_issue_packs_0_T_97_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_branch_predict_pack_valid = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_97_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_branch_predict_pack_target = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_97_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_98_branch_predict_pack_branch_type = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_97_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_branch_predict_pack_select = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_97_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_branch_predict_pack_taken = _issue1_func_code_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_97_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_phy_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_97_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_stale_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_97_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_arch_dst = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_97_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_98_inst_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_97_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_regWen = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_regWen :
    _io_o_issue_packs_0_T_97_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_src1_valid = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_97_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_phy_rs1 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_97_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_arch_rs1 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_97_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_98_src2_valid = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_97_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_phy_rs2 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_97_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_arch_rs2 = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_97_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_98_rob_idx = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_97_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_imm = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_imm :
    _io_o_issue_packs_0_T_97_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_src1_value = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_97_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_98_src2_value = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_97_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_98_op1_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_97_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_98_op2_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_97_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_98_alu_sel = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_97_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_98_branch_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_97_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_98_mem_type = _issue1_func_code_T_29 ? reservation_station_29_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_97_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_99_pc = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_pc :
    _io_o_issue_packs_0_T_98_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_99_inst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_inst :
    _io_o_issue_packs_0_T_98_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_func_code = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_func_code :
    _io_o_issue_packs_0_T_98_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_branch_predict_pack_valid = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_98_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_branch_predict_pack_target = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_98_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_99_branch_predict_pack_branch_type = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_98_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_branch_predict_pack_select = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_98_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_branch_predict_pack_taken = _issue1_func_code_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_98_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_phy_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_98_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_stale_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_98_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_arch_dst = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_98_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_99_inst_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_98_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_regWen = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_regWen :
    _io_o_issue_packs_0_T_98_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_src1_valid = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_98_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_phy_rs1 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_98_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_arch_rs1 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_98_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_99_src2_valid = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_98_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_phy_rs2 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_98_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_arch_rs2 = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_98_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_99_rob_idx = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_98_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_imm = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_imm :
    _io_o_issue_packs_0_T_98_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_src1_value = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_98_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_99_src2_value = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_98_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_99_op1_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_98_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_99_op2_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_98_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_99_alu_sel = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_98_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_99_branch_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_98_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_99_mem_type = _issue1_func_code_T_28 ? reservation_station_28_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_98_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_100_pc = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_pc :
    _io_o_issue_packs_0_T_99_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_100_inst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_inst :
    _io_o_issue_packs_0_T_99_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_func_code = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_func_code :
    _io_o_issue_packs_0_T_99_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_branch_predict_pack_valid = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_99_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_branch_predict_pack_target = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_99_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_100_branch_predict_pack_branch_type = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_99_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_branch_predict_pack_select = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_99_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_branch_predict_pack_taken = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_99_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_phy_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_99_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_stale_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_99_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_arch_dst = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_99_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_100_inst_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_99_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_regWen = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_regWen :
    _io_o_issue_packs_0_T_99_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_src1_valid = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_99_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_phy_rs1 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_99_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_arch_rs1 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_99_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_100_src2_valid = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_99_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_phy_rs2 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_99_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_arch_rs2 = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_99_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_100_rob_idx = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_99_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_imm = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_imm :
    _io_o_issue_packs_0_T_99_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_src1_value = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_99_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_100_src2_value = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_99_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_100_op1_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_99_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_100_op2_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_99_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_100_alu_sel = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_99_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_100_branch_type = _issue1_func_code_T_27 ?
    reservation_station_27_io_o_uop_branch_type : _io_o_issue_packs_0_T_99_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_100_mem_type = _issue1_func_code_T_27 ? reservation_station_27_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_99_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_101_pc = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_pc :
    _io_o_issue_packs_0_T_100_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_101_inst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_inst :
    _io_o_issue_packs_0_T_100_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_func_code = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_func_code :
    _io_o_issue_packs_0_T_100_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_branch_predict_pack_valid = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_100_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_branch_predict_pack_target = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_100_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_101_branch_predict_pack_branch_type = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_100_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_branch_predict_pack_select = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_100_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_branch_predict_pack_taken = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_100_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_phy_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_100_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_stale_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_100_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_arch_dst = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_100_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_101_inst_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_100_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_regWen = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_regWen :
    _io_o_issue_packs_0_T_100_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_src1_valid = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_100_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_phy_rs1 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_100_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_arch_rs1 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_100_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_101_src2_valid = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_100_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_phy_rs2 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_100_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_arch_rs2 = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_100_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_101_rob_idx = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_100_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_imm = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_imm :
    _io_o_issue_packs_0_T_100_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_src1_value = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_100_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_101_src2_value = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_100_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_101_op1_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_100_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_101_op2_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_100_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_101_alu_sel = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_100_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_101_branch_type = _issue1_func_code_T_26 ?
    reservation_station_26_io_o_uop_branch_type : _io_o_issue_packs_0_T_100_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_101_mem_type = _issue1_func_code_T_26 ? reservation_station_26_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_100_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_102_pc = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_pc :
    _io_o_issue_packs_0_T_101_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_102_inst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_inst :
    _io_o_issue_packs_0_T_101_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_func_code = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_func_code :
    _io_o_issue_packs_0_T_101_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_branch_predict_pack_valid = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_101_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_branch_predict_pack_target = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_101_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_102_branch_predict_pack_branch_type = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_101_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_branch_predict_pack_select = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_101_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_branch_predict_pack_taken = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_101_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_phy_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_101_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_stale_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_101_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_arch_dst = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_101_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_102_inst_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_101_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_regWen = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_regWen :
    _io_o_issue_packs_0_T_101_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_src1_valid = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_101_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_phy_rs1 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_101_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_arch_rs1 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_101_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_102_src2_valid = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_101_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_phy_rs2 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_101_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_arch_rs2 = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_101_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_102_rob_idx = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_101_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_imm = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_imm :
    _io_o_issue_packs_0_T_101_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_src1_value = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_101_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_102_src2_value = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_101_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_102_op1_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_101_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_102_op2_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_101_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_102_alu_sel = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_101_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_102_branch_type = _issue1_func_code_T_25 ?
    reservation_station_25_io_o_uop_branch_type : _io_o_issue_packs_0_T_101_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_102_mem_type = _issue1_func_code_T_25 ? reservation_station_25_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_101_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_103_pc = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_pc :
    _io_o_issue_packs_0_T_102_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_103_inst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_inst :
    _io_o_issue_packs_0_T_102_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_func_code = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_func_code :
    _io_o_issue_packs_0_T_102_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_branch_predict_pack_valid = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_102_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_branch_predict_pack_target = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_102_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_103_branch_predict_pack_branch_type = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_102_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_branch_predict_pack_select = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_102_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_branch_predict_pack_taken = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_102_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_phy_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_102_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_stale_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_102_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_arch_dst = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_102_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_103_inst_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_102_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_regWen = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_regWen :
    _io_o_issue_packs_0_T_102_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_src1_valid = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_102_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_phy_rs1 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_102_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_arch_rs1 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_102_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_103_src2_valid = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_102_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_phy_rs2 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_102_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_arch_rs2 = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_102_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_103_rob_idx = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_102_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_imm = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_imm :
    _io_o_issue_packs_0_T_102_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_src1_value = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_102_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_103_src2_value = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_102_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_103_op1_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_102_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_103_op2_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_102_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_103_alu_sel = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_102_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_103_branch_type = _issue1_func_code_T_24 ?
    reservation_station_24_io_o_uop_branch_type : _io_o_issue_packs_0_T_102_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_103_mem_type = _issue1_func_code_T_24 ? reservation_station_24_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_102_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_104_pc = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_pc :
    _io_o_issue_packs_0_T_103_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_104_inst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_inst :
    _io_o_issue_packs_0_T_103_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_func_code = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_func_code :
    _io_o_issue_packs_0_T_103_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_branch_predict_pack_valid = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_103_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_branch_predict_pack_target = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_103_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_104_branch_predict_pack_branch_type = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_103_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_branch_predict_pack_select = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_103_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_branch_predict_pack_taken = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_103_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_phy_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_103_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_stale_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_103_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_arch_dst = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_103_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_104_inst_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_103_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_regWen = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_regWen :
    _io_o_issue_packs_0_T_103_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_src1_valid = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_103_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_phy_rs1 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_103_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_arch_rs1 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_103_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_104_src2_valid = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_103_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_phy_rs2 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_103_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_arch_rs2 = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_103_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_104_rob_idx = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_103_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_imm = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_imm :
    _io_o_issue_packs_0_T_103_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_src1_value = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_103_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_104_src2_value = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_103_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_104_op1_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_103_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_104_op2_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_103_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_104_alu_sel = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_103_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_104_branch_type = _issue1_func_code_T_23 ?
    reservation_station_23_io_o_uop_branch_type : _io_o_issue_packs_0_T_103_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_104_mem_type = _issue1_func_code_T_23 ? reservation_station_23_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_103_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_105_pc = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_pc :
    _io_o_issue_packs_0_T_104_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_105_inst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_inst :
    _io_o_issue_packs_0_T_104_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_func_code = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_func_code :
    _io_o_issue_packs_0_T_104_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_branch_predict_pack_valid = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_104_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_branch_predict_pack_target = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_104_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_105_branch_predict_pack_branch_type = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_104_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_branch_predict_pack_select = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_104_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_branch_predict_pack_taken = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_104_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_phy_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_104_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_stale_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_104_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_arch_dst = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_104_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_105_inst_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_104_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_regWen = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_regWen :
    _io_o_issue_packs_0_T_104_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_src1_valid = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_104_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_phy_rs1 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_104_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_arch_rs1 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_104_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_105_src2_valid = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_104_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_phy_rs2 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_104_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_arch_rs2 = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_104_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_105_rob_idx = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_104_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_imm = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_imm :
    _io_o_issue_packs_0_T_104_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_src1_value = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_104_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_105_src2_value = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_104_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_105_op1_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_104_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_105_op2_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_104_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_105_alu_sel = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_104_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_105_branch_type = _issue1_func_code_T_22 ?
    reservation_station_22_io_o_uop_branch_type : _io_o_issue_packs_0_T_104_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_105_mem_type = _issue1_func_code_T_22 ? reservation_station_22_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_104_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_106_pc = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_pc :
    _io_o_issue_packs_0_T_105_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_106_inst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_inst :
    _io_o_issue_packs_0_T_105_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_func_code = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_func_code :
    _io_o_issue_packs_0_T_105_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_branch_predict_pack_valid = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_105_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_branch_predict_pack_target = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_105_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_106_branch_predict_pack_branch_type = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_105_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_branch_predict_pack_select = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_105_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_branch_predict_pack_taken = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_105_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_phy_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_105_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_stale_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_105_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_arch_dst = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_105_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_106_inst_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_105_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_regWen = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_regWen :
    _io_o_issue_packs_0_T_105_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_src1_valid = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_105_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_phy_rs1 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_105_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_arch_rs1 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_105_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_106_src2_valid = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_105_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_phy_rs2 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_105_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_arch_rs2 = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_105_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_106_rob_idx = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_105_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_imm = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_imm :
    _io_o_issue_packs_0_T_105_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_src1_value = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_105_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_106_src2_value = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_105_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_106_op1_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_105_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_106_op2_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_105_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_106_alu_sel = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_105_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_106_branch_type = _issue1_func_code_T_21 ?
    reservation_station_21_io_o_uop_branch_type : _io_o_issue_packs_0_T_105_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_106_mem_type = _issue1_func_code_T_21 ? reservation_station_21_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_105_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_107_pc = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_pc :
    _io_o_issue_packs_0_T_106_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_107_inst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_inst :
    _io_o_issue_packs_0_T_106_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_func_code = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_func_code :
    _io_o_issue_packs_0_T_106_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_branch_predict_pack_valid = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_106_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_branch_predict_pack_target = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_106_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_107_branch_predict_pack_branch_type = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_106_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_branch_predict_pack_select = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_106_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_branch_predict_pack_taken = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_106_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_phy_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_106_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_stale_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_106_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_arch_dst = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_106_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_107_inst_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_106_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_regWen = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_regWen :
    _io_o_issue_packs_0_T_106_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_src1_valid = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_106_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_phy_rs1 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_106_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_arch_rs1 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_106_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_107_src2_valid = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_106_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_phy_rs2 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_106_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_arch_rs2 = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_106_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_107_rob_idx = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_106_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_imm = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_imm :
    _io_o_issue_packs_0_T_106_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_src1_value = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_106_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_107_src2_value = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_106_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_107_op1_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_106_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_107_op2_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_106_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_107_alu_sel = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_106_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_107_branch_type = _issue1_func_code_T_20 ?
    reservation_station_20_io_o_uop_branch_type : _io_o_issue_packs_0_T_106_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_107_mem_type = _issue1_func_code_T_20 ? reservation_station_20_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_106_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_108_pc = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_pc :
    _io_o_issue_packs_0_T_107_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_108_inst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_inst :
    _io_o_issue_packs_0_T_107_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_func_code = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_func_code :
    _io_o_issue_packs_0_T_107_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_branch_predict_pack_valid = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_107_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_branch_predict_pack_target = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_107_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_108_branch_predict_pack_branch_type = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_107_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_branch_predict_pack_select = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_107_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_branch_predict_pack_taken = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_107_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_phy_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_107_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_stale_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_107_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_arch_dst = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_107_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_108_inst_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_107_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_regWen = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_regWen :
    _io_o_issue_packs_0_T_107_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_src1_valid = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_107_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_phy_rs1 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_107_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_arch_rs1 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_107_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_108_src2_valid = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_107_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_phy_rs2 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_107_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_arch_rs2 = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_107_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_108_rob_idx = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_107_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_imm = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_imm :
    _io_o_issue_packs_0_T_107_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_src1_value = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_107_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_108_src2_value = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_107_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_108_op1_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_107_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_108_op2_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_107_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_108_alu_sel = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_107_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_108_branch_type = _issue1_func_code_T_19 ?
    reservation_station_19_io_o_uop_branch_type : _io_o_issue_packs_0_T_107_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_108_mem_type = _issue1_func_code_T_19 ? reservation_station_19_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_107_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_109_pc = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_pc :
    _io_o_issue_packs_0_T_108_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_109_inst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_inst :
    _io_o_issue_packs_0_T_108_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_func_code = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_func_code :
    _io_o_issue_packs_0_T_108_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_branch_predict_pack_valid = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_108_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_branch_predict_pack_target = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_108_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_109_branch_predict_pack_branch_type = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_108_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_branch_predict_pack_select = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_108_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_branch_predict_pack_taken = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_108_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_phy_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_108_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_stale_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_108_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_arch_dst = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_108_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_109_inst_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_108_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_regWen = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_regWen :
    _io_o_issue_packs_0_T_108_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_src1_valid = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_108_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_phy_rs1 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_108_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_arch_rs1 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_108_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_109_src2_valid = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_108_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_phy_rs2 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_108_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_arch_rs2 = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_108_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_109_rob_idx = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_108_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_imm = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_imm :
    _io_o_issue_packs_0_T_108_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_src1_value = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_108_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_109_src2_value = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_108_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_109_op1_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_108_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_109_op2_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_108_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_109_alu_sel = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_108_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_109_branch_type = _issue1_func_code_T_18 ?
    reservation_station_18_io_o_uop_branch_type : _io_o_issue_packs_0_T_108_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_109_mem_type = _issue1_func_code_T_18 ? reservation_station_18_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_108_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_110_pc = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_pc :
    _io_o_issue_packs_0_T_109_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_110_inst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_inst :
    _io_o_issue_packs_0_T_109_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_func_code = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_func_code :
    _io_o_issue_packs_0_T_109_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_branch_predict_pack_valid = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_109_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_branch_predict_pack_target = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_109_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_110_branch_predict_pack_branch_type = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_109_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_branch_predict_pack_select = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_109_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_branch_predict_pack_taken = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_109_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_phy_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_109_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_stale_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_109_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_arch_dst = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_109_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_110_inst_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_109_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_regWen = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_regWen :
    _io_o_issue_packs_0_T_109_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_src1_valid = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_109_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_phy_rs1 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_109_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_arch_rs1 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_109_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_110_src2_valid = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_109_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_phy_rs2 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_109_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_arch_rs2 = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_109_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_110_rob_idx = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_109_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_imm = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_imm :
    _io_o_issue_packs_0_T_109_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_src1_value = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_109_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_110_src2_value = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_109_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_110_op1_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_109_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_110_op2_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_109_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_110_alu_sel = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_109_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_110_branch_type = _issue1_func_code_T_17 ?
    reservation_station_17_io_o_uop_branch_type : _io_o_issue_packs_0_T_109_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_110_mem_type = _issue1_func_code_T_17 ? reservation_station_17_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_109_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_111_pc = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_pc :
    _io_o_issue_packs_0_T_110_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_111_inst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_inst :
    _io_o_issue_packs_0_T_110_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_func_code = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_func_code :
    _io_o_issue_packs_0_T_110_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_branch_predict_pack_valid = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_110_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_branch_predict_pack_target = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_110_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_111_branch_predict_pack_branch_type = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_110_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_branch_predict_pack_select = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_110_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_branch_predict_pack_taken = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_110_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_phy_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_110_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_stale_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_110_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_arch_dst = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_110_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_111_inst_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_110_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_regWen = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_regWen :
    _io_o_issue_packs_0_T_110_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_src1_valid = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_110_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_phy_rs1 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_110_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_arch_rs1 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_110_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_111_src2_valid = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_110_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_phy_rs2 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_110_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_arch_rs2 = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_110_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_111_rob_idx = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_110_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_imm = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_imm :
    _io_o_issue_packs_0_T_110_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_src1_value = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_110_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_111_src2_value = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_110_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_111_op1_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_110_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_111_op2_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_110_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_111_alu_sel = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_110_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_111_branch_type = _issue1_func_code_T_16 ?
    reservation_station_16_io_o_uop_branch_type : _io_o_issue_packs_0_T_110_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_111_mem_type = _issue1_func_code_T_16 ? reservation_station_16_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_110_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_112_pc = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_pc :
    _io_o_issue_packs_0_T_111_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_112_inst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_inst :
    _io_o_issue_packs_0_T_111_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_func_code = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_func_code :
    _io_o_issue_packs_0_T_111_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_branch_predict_pack_valid = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_111_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_branch_predict_pack_target = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_111_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_112_branch_predict_pack_branch_type = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_111_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_branch_predict_pack_select = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_111_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_branch_predict_pack_taken = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_111_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_phy_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_111_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_stale_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_111_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_arch_dst = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_111_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_112_inst_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_111_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_regWen = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_regWen :
    _io_o_issue_packs_0_T_111_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_src1_valid = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_111_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_phy_rs1 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_111_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_arch_rs1 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_111_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_112_src2_valid = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_111_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_phy_rs2 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_111_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_arch_rs2 = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_111_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_112_rob_idx = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_111_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_imm = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_imm :
    _io_o_issue_packs_0_T_111_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_src1_value = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_111_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_112_src2_value = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_111_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_112_op1_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_111_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_112_op2_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_111_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_112_alu_sel = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_111_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_112_branch_type = _issue1_func_code_T_15 ?
    reservation_station_15_io_o_uop_branch_type : _io_o_issue_packs_0_T_111_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_112_mem_type = _issue1_func_code_T_15 ? reservation_station_15_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_111_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_113_pc = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_pc :
    _io_o_issue_packs_0_T_112_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_113_inst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_inst :
    _io_o_issue_packs_0_T_112_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_func_code = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_func_code :
    _io_o_issue_packs_0_T_112_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_branch_predict_pack_valid = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_112_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_branch_predict_pack_target = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_112_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_113_branch_predict_pack_branch_type = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_112_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_branch_predict_pack_select = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_112_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_branch_predict_pack_taken = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_112_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_phy_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_112_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_stale_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_112_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_arch_dst = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_112_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_113_inst_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_112_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_regWen = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_regWen :
    _io_o_issue_packs_0_T_112_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_src1_valid = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_112_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_phy_rs1 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_112_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_arch_rs1 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_112_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_113_src2_valid = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_112_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_phy_rs2 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_112_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_arch_rs2 = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_112_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_113_rob_idx = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_112_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_imm = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_imm :
    _io_o_issue_packs_0_T_112_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_src1_value = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_112_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_113_src2_value = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_112_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_113_op1_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_112_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_113_op2_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_112_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_113_alu_sel = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_112_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_113_branch_type = _issue1_func_code_T_14 ?
    reservation_station_14_io_o_uop_branch_type : _io_o_issue_packs_0_T_112_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_113_mem_type = _issue1_func_code_T_14 ? reservation_station_14_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_112_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_114_pc = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_pc :
    _io_o_issue_packs_0_T_113_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_114_inst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_inst :
    _io_o_issue_packs_0_T_113_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_func_code = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_func_code :
    _io_o_issue_packs_0_T_113_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_branch_predict_pack_valid = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_113_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_branch_predict_pack_target = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_113_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_114_branch_predict_pack_branch_type = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_113_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_branch_predict_pack_select = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_113_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_branch_predict_pack_taken = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_113_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_phy_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_113_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_stale_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_113_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_arch_dst = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_113_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_114_inst_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_113_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_regWen = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_regWen :
    _io_o_issue_packs_0_T_113_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_src1_valid = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_113_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_phy_rs1 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_113_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_arch_rs1 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_113_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_114_src2_valid = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_113_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_phy_rs2 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_113_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_arch_rs2 = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_113_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_114_rob_idx = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_113_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_imm = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_imm :
    _io_o_issue_packs_0_T_113_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_src1_value = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_113_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_114_src2_value = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_113_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_114_op1_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_113_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_114_op2_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_113_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_114_alu_sel = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_113_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_114_branch_type = _issue1_func_code_T_13 ?
    reservation_station_13_io_o_uop_branch_type : _io_o_issue_packs_0_T_113_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_114_mem_type = _issue1_func_code_T_13 ? reservation_station_13_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_113_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_115_pc = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_pc :
    _io_o_issue_packs_0_T_114_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_115_inst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_inst :
    _io_o_issue_packs_0_T_114_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_func_code = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_func_code :
    _io_o_issue_packs_0_T_114_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_branch_predict_pack_valid = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_114_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_branch_predict_pack_target = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_114_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_115_branch_predict_pack_branch_type = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_114_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_branch_predict_pack_select = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_114_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_branch_predict_pack_taken = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_114_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_phy_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_114_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_stale_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_114_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_arch_dst = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_114_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_115_inst_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_114_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_regWen = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_regWen :
    _io_o_issue_packs_0_T_114_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_src1_valid = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_114_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_phy_rs1 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_114_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_arch_rs1 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_114_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_115_src2_valid = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_114_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_phy_rs2 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_114_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_arch_rs2 = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_114_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_115_rob_idx = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_114_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_imm = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_imm :
    _io_o_issue_packs_0_T_114_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_src1_value = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_114_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_115_src2_value = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_114_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_115_op1_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_114_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_115_op2_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_114_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_115_alu_sel = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_114_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_115_branch_type = _issue1_func_code_T_12 ?
    reservation_station_12_io_o_uop_branch_type : _io_o_issue_packs_0_T_114_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_115_mem_type = _issue1_func_code_T_12 ? reservation_station_12_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_114_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_116_pc = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_pc :
    _io_o_issue_packs_0_T_115_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_116_inst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_inst :
    _io_o_issue_packs_0_T_115_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_func_code = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_func_code :
    _io_o_issue_packs_0_T_115_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_branch_predict_pack_valid = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_115_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_branch_predict_pack_target = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_115_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_116_branch_predict_pack_branch_type = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_115_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_branch_predict_pack_select = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_115_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_branch_predict_pack_taken = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_115_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_phy_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_115_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_stale_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_115_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_arch_dst = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_115_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_116_inst_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_115_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_regWen = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_regWen :
    _io_o_issue_packs_0_T_115_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_src1_valid = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_115_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_phy_rs1 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_115_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_arch_rs1 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_115_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_116_src2_valid = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_115_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_phy_rs2 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_115_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_arch_rs2 = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_115_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_116_rob_idx = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_115_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_imm = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_imm :
    _io_o_issue_packs_0_T_115_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_src1_value = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_115_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_116_src2_value = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_115_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_116_op1_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_115_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_116_op2_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_115_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_116_alu_sel = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_115_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_116_branch_type = _issue1_func_code_T_11 ?
    reservation_station_11_io_o_uop_branch_type : _io_o_issue_packs_0_T_115_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_116_mem_type = _issue1_func_code_T_11 ? reservation_station_11_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_115_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_117_pc = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_pc :
    _io_o_issue_packs_0_T_116_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_117_inst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_inst :
    _io_o_issue_packs_0_T_116_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_func_code = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_func_code :
    _io_o_issue_packs_0_T_116_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_branch_predict_pack_valid = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_116_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_branch_predict_pack_target = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_116_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_117_branch_predict_pack_branch_type = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_116_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_branch_predict_pack_select = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_116_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_branch_predict_pack_taken = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_116_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_phy_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_116_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_stale_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_116_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_arch_dst = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_116_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_117_inst_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_116_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_regWen = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_regWen :
    _io_o_issue_packs_0_T_116_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_src1_valid = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_116_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_phy_rs1 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_116_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_arch_rs1 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_116_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_117_src2_valid = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_116_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_phy_rs2 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_116_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_arch_rs2 = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_116_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_117_rob_idx = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_116_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_imm = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_imm :
    _io_o_issue_packs_0_T_116_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_src1_value = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_116_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_117_src2_value = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_116_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_117_op1_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_116_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_117_op2_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_116_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_117_alu_sel = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_116_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_117_branch_type = _issue1_func_code_T_10 ?
    reservation_station_10_io_o_uop_branch_type : _io_o_issue_packs_0_T_116_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_117_mem_type = _issue1_func_code_T_10 ? reservation_station_10_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_116_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_118_pc = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_pc :
    _io_o_issue_packs_0_T_117_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_118_inst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_inst :
    _io_o_issue_packs_0_T_117_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_func_code = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_func_code :
    _io_o_issue_packs_0_T_117_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_branch_predict_pack_valid = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_117_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_branch_predict_pack_target = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_117_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_118_branch_predict_pack_branch_type = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_117_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_branch_predict_pack_select = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_117_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_branch_predict_pack_taken = _issue1_func_code_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_117_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_phy_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_117_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_stale_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_117_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_arch_dst = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_117_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_118_inst_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_117_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_regWen = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_regWen :
    _io_o_issue_packs_0_T_117_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_src1_valid = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_117_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_phy_rs1 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_117_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_arch_rs1 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_117_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_118_src2_valid = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_117_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_phy_rs2 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_117_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_arch_rs2 = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_117_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_118_rob_idx = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_117_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_imm = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_imm :
    _io_o_issue_packs_0_T_117_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_src1_value = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_117_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_118_src2_value = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_117_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_118_op1_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_117_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_118_op2_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_117_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_118_alu_sel = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_117_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_118_branch_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_117_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_118_mem_type = _issue1_func_code_T_9 ? reservation_station_9_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_117_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_119_pc = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_pc :
    _io_o_issue_packs_0_T_118_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_119_inst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_inst :
    _io_o_issue_packs_0_T_118_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_func_code = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_func_code :
    _io_o_issue_packs_0_T_118_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_branch_predict_pack_valid = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_118_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_branch_predict_pack_target = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_118_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_119_branch_predict_pack_branch_type = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_118_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_branch_predict_pack_select = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_118_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_branch_predict_pack_taken = _issue1_func_code_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_118_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_phy_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_118_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_stale_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_118_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_arch_dst = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_118_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_119_inst_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_118_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_regWen = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_regWen :
    _io_o_issue_packs_0_T_118_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_src1_valid = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_118_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_phy_rs1 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_118_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_arch_rs1 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_118_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_119_src2_valid = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_118_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_phy_rs2 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_118_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_arch_rs2 = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_118_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_119_rob_idx = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_118_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_imm = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_imm :
    _io_o_issue_packs_0_T_118_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_src1_value = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_118_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_119_src2_value = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_118_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_119_op1_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_118_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_119_op2_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_118_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_119_alu_sel = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_118_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_119_branch_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_118_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_119_mem_type = _issue1_func_code_T_8 ? reservation_station_8_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_118_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_120_pc = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_pc :
    _io_o_issue_packs_0_T_119_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_120_inst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_inst :
    _io_o_issue_packs_0_T_119_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_func_code = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_func_code :
    _io_o_issue_packs_0_T_119_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_branch_predict_pack_valid = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_119_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_branch_predict_pack_target = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_119_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_120_branch_predict_pack_branch_type = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_119_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_branch_predict_pack_select = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_119_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_branch_predict_pack_taken = _issue1_func_code_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_119_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_phy_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_119_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_stale_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_119_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_arch_dst = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_119_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_120_inst_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_119_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_regWen = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_regWen :
    _io_o_issue_packs_0_T_119_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_src1_valid = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_119_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_phy_rs1 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_119_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_arch_rs1 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_119_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_120_src2_valid = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_119_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_phy_rs2 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_119_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_arch_rs2 = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_119_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_120_rob_idx = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_119_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_imm = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_imm :
    _io_o_issue_packs_0_T_119_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_src1_value = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_119_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_120_src2_value = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_119_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_120_op1_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_119_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_120_op2_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_119_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_120_alu_sel = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_119_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_120_branch_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_119_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_120_mem_type = _issue1_func_code_T_7 ? reservation_station_7_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_119_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_121_pc = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_pc :
    _io_o_issue_packs_0_T_120_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_121_inst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_inst :
    _io_o_issue_packs_0_T_120_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_func_code = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_func_code :
    _io_o_issue_packs_0_T_120_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_branch_predict_pack_valid = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_120_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_branch_predict_pack_target = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_120_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_121_branch_predict_pack_branch_type = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_120_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_branch_predict_pack_select = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_120_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_branch_predict_pack_taken = _issue1_func_code_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_120_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_phy_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_120_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_stale_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_120_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_arch_dst = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_120_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_121_inst_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_120_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_regWen = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_regWen :
    _io_o_issue_packs_0_T_120_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_src1_valid = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_120_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_phy_rs1 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_120_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_arch_rs1 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_120_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_121_src2_valid = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_120_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_phy_rs2 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_120_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_arch_rs2 = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_120_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_121_rob_idx = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_120_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_imm = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_imm :
    _io_o_issue_packs_0_T_120_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_src1_value = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_120_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_121_src2_value = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_120_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_121_op1_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_120_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_121_op2_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_120_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_121_alu_sel = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_120_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_121_branch_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_120_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_121_mem_type = _issue1_func_code_T_6 ? reservation_station_6_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_120_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_122_pc = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_pc :
    _io_o_issue_packs_0_T_121_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_122_inst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_inst :
    _io_o_issue_packs_0_T_121_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_func_code = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_func_code :
    _io_o_issue_packs_0_T_121_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_branch_predict_pack_valid = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_121_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_branch_predict_pack_target = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_121_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_122_branch_predict_pack_branch_type = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_121_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_branch_predict_pack_select = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_121_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_branch_predict_pack_taken = _issue1_func_code_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_121_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_phy_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_121_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_stale_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_121_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_arch_dst = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_121_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_122_inst_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_121_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_regWen = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_regWen :
    _io_o_issue_packs_0_T_121_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_src1_valid = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_121_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_phy_rs1 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_121_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_arch_rs1 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_121_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_122_src2_valid = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_121_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_phy_rs2 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_121_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_arch_rs2 = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_121_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_122_rob_idx = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_121_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_imm = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_imm :
    _io_o_issue_packs_0_T_121_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_src1_value = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_121_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_122_src2_value = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_121_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_122_op1_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_121_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_122_op2_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_121_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_122_alu_sel = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_121_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_122_branch_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_121_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_122_mem_type = _issue1_func_code_T_5 ? reservation_station_5_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_121_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_123_pc = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_pc :
    _io_o_issue_packs_0_T_122_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_123_inst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_inst :
    _io_o_issue_packs_0_T_122_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_func_code = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_func_code :
    _io_o_issue_packs_0_T_122_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_branch_predict_pack_valid = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_122_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_branch_predict_pack_target = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_122_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_123_branch_predict_pack_branch_type = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_122_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_branch_predict_pack_select = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_122_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_branch_predict_pack_taken = _issue1_func_code_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_122_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_phy_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_122_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_stale_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_122_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_arch_dst = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_122_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_123_inst_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_122_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_regWen = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_regWen :
    _io_o_issue_packs_0_T_122_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_src1_valid = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_122_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_phy_rs1 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_122_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_arch_rs1 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_122_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_123_src2_valid = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_122_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_phy_rs2 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_122_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_arch_rs2 = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_122_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_123_rob_idx = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_122_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_imm = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_imm :
    _io_o_issue_packs_0_T_122_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_src1_value = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_122_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_123_src2_value = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_122_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_123_op1_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_122_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_123_op2_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_122_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_123_alu_sel = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_122_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_123_branch_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_122_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_123_mem_type = _issue1_func_code_T_4 ? reservation_station_4_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_122_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_124_pc = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_pc :
    _io_o_issue_packs_0_T_123_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_124_inst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_inst :
    _io_o_issue_packs_0_T_123_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_func_code = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_func_code :
    _io_o_issue_packs_0_T_123_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_branch_predict_pack_valid = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_123_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_branch_predict_pack_target = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_123_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_124_branch_predict_pack_branch_type = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_123_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_branch_predict_pack_select = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_123_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_branch_predict_pack_taken = _issue1_func_code_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_123_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_phy_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_123_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_stale_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_123_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_arch_dst = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_123_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_124_inst_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_123_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_regWen = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_regWen :
    _io_o_issue_packs_0_T_123_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_src1_valid = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_123_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_phy_rs1 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_123_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_arch_rs1 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_123_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_124_src2_valid = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_123_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_phy_rs2 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_123_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_arch_rs2 = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_123_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_124_rob_idx = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_123_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_imm = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_imm :
    _io_o_issue_packs_0_T_123_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_src1_value = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_123_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_124_src2_value = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_123_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_124_op1_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_123_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_124_op2_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_123_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_124_alu_sel = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_123_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_124_branch_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_123_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_124_mem_type = _issue1_func_code_T_3 ? reservation_station_3_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_123_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_125_pc = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_pc :
    _io_o_issue_packs_0_T_124_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_125_inst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_inst :
    _io_o_issue_packs_0_T_124_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_func_code = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_func_code :
    _io_o_issue_packs_0_T_124_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_branch_predict_pack_valid = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_124_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_branch_predict_pack_target = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_124_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_125_branch_predict_pack_branch_type = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_124_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_branch_predict_pack_select = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_124_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_branch_predict_pack_taken = _issue1_func_code_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_124_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_phy_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_124_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_stale_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_124_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_arch_dst = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_124_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_125_inst_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_124_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_regWen = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_regWen :
    _io_o_issue_packs_0_T_124_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_src1_valid = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_124_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_phy_rs1 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_124_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_arch_rs1 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_124_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_125_src2_valid = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_124_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_phy_rs2 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_124_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_arch_rs2 = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_124_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_125_rob_idx = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_124_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_imm = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_imm :
    _io_o_issue_packs_0_T_124_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_src1_value = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_124_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_125_src2_value = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_124_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_125_op1_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_124_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_125_op2_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_124_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_125_alu_sel = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_124_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_125_branch_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_124_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_125_mem_type = _issue1_func_code_T_2 ? reservation_station_2_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_124_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_126_pc = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_pc :
    _io_o_issue_packs_0_T_125_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_0_T_126_inst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_inst :
    _io_o_issue_packs_0_T_125_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_func_code = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_func_code :
    _io_o_issue_packs_0_T_125_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_branch_predict_pack_valid = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_125_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_branch_predict_pack_target = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_125_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_126_branch_predict_pack_branch_type = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_125_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_branch_predict_pack_select = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_125_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_branch_predict_pack_taken = _issue1_func_code_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_125_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_phy_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_125_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_stale_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_125_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_arch_dst = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_125_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_126_inst_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_125_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_regWen = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_regWen :
    _io_o_issue_packs_0_T_125_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_src1_valid = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_125_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_phy_rs1 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_125_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_arch_rs1 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_125_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_0_T_126_src2_valid = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_125_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_phy_rs2 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_125_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_arch_rs2 = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_125_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_0_T_126_rob_idx = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_125_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_imm = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_imm :
    _io_o_issue_packs_0_T_125_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_src1_value = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src1_value
     : _io_o_issue_packs_0_T_125_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_0_T_126_src2_value = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_src2_value
     : _io_o_issue_packs_0_T_125_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_126_op1_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_125_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_0_T_126_op2_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_125_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_0_T_126_alu_sel = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_125_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_0_T_126_branch_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_branch_type
     : _io_o_issue_packs_0_T_125_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_0_T_126_mem_type = _issue1_func_code_T_1 ? reservation_station_1_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_125_mem_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T = 6'h0 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_1 = 6'h1 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_2 = 6'h2 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_3 = 6'h3 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_4 = 6'h4 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_5 = 6'h5 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_6 = 6'h6 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_7 = 6'h7 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_8 = 6'h8 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_9 = 6'h9 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_10 = 6'ha == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_11 = 6'hb == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_12 = 6'hc == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_13 = 6'hd == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_14 = 6'he == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_15 = 6'hf == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_16 = 6'h10 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_17 = 6'h11 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_18 = 6'h12 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_19 = 6'h13 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_20 = 6'h14 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_21 = 6'h15 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_22 = 6'h16 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_23 = 6'h17 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_24 = 6'h18 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_25 = 6'h19 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_26 = 6'h1a == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_27 = 6'h1b == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_28 = 6'h1c == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_29 = 6'h1d == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_30 = 6'h1e == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_31 = 6'h1f == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_32 = 6'h20 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_33 = 6'h21 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_34 = 6'h22 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_35 = 6'h23 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_36 = 6'h24 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_37 = 6'h25 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_38 = 6'h26 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_39 = 6'h27 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_40 = 6'h28 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_41 = 6'h29 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_42 = 6'h2a == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_43 = 6'h2b == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_44 = 6'h2c == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_45 = 6'h2d == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_46 = 6'h2e == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_47 = 6'h2f == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_48 = 6'h30 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_49 = 6'h31 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_50 = 6'h32 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_51 = 6'h33 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_52 = 6'h34 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_53 = 6'h35 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_54 = 6'h36 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_55 = 6'h37 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_56 = 6'h38 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_57 = 6'h39 == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_58 = 6'h3a == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_59 = 6'h3b == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_60 = 6'h3c == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_61 = 6'h3d == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_62 = 6'h3e == issue2_idx; // @[reservation_station.scala 107:94]
  wire  _io_o_issue_packs_1_T_63 = 6'h3f == issue2_idx; // @[reservation_station.scala 107:94]
  wire [31:0] _io_o_issue_packs_1_T_64_pc = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_pc :
    reservation_station_0_io_o_uop_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_64_inst = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_inst :
    reservation_station_0_io_o_uop_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_func_code = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_func_code
     : reservation_station_0_io_o_uop_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_branch_predict_pack_valid = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_valid : reservation_station_0_io_o_uop_branch_predict_pack_valid
    ; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_branch_predict_pack_target = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_target :
    reservation_station_0_io_o_uop_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_64_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_branch_type :
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_branch_predict_pack_select = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_select :
    reservation_station_0_io_o_uop_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_branch_predict_pack_taken = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_branch_predict_pack_taken : reservation_station_0_io_o_uop_branch_predict_pack_taken
    ; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_phy_dst = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_phy_dst :
    reservation_station_0_io_o_uop_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_stale_dst = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_stale_dst
     : reservation_station_0_io_o_uop_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_arch_dst = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_arch_dst :
    reservation_station_0_io_o_uop_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_64_inst_type = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_inst_type
     : reservation_station_0_io_o_uop_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_regWen = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_regWen :
    reservation_station_0_io_o_uop_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_src1_valid = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_src1_valid :
    reservation_station_0_io_o_uop_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_phy_rs1 = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_phy_rs1 :
    reservation_station_0_io_o_uop_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_arch_rs1 = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_arch_rs1 :
    reservation_station_0_io_o_uop_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_64_src2_valid = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_src2_valid :
    reservation_station_0_io_o_uop_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_phy_rs2 = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_phy_rs2 :
    reservation_station_0_io_o_uop_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_arch_rs2 = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_arch_rs2 :
    reservation_station_0_io_o_uop_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_64_rob_idx = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_rob_idx :
    reservation_station_0_io_o_uop_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_imm = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_imm :
    reservation_station_0_io_o_uop_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_src1_value = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_src1_value : reservation_station_0_io_o_uop_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_64_src2_value = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_src2_value : reservation_station_0_io_o_uop_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_64_op1_sel = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_op1_sel :
    reservation_station_0_io_o_uop_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_64_op2_sel = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_op2_sel :
    reservation_station_0_io_o_uop_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_64_alu_sel = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_alu_sel :
    reservation_station_0_io_o_uop_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_64_branch_type = _io_o_issue_packs_1_T_63 ?
    reservation_station_63_io_o_uop_branch_type : reservation_station_0_io_o_uop_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_64_mem_type = _io_o_issue_packs_1_T_63 ? reservation_station_63_io_o_uop_mem_type :
    reservation_station_0_io_o_uop_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_65_pc = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_pc :
    _io_o_issue_packs_1_T_64_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_65_inst = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_inst :
    _io_o_issue_packs_1_T_64_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_func_code = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_func_code
     : _io_o_issue_packs_1_T_64_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_branch_predict_pack_valid = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_64_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_branch_predict_pack_target = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_64_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_65_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_64_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_branch_predict_pack_select = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_64_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_branch_predict_pack_taken = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_64_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_phy_dst = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_64_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_stale_dst = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_64_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_arch_dst = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_64_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_65_inst_type = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_64_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_regWen = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_regWen :
    _io_o_issue_packs_1_T_64_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_src1_valid = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_64_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_phy_rs1 = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_64_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_arch_rs1 = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_64_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_65_src2_valid = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_64_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_phy_rs2 = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_64_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_arch_rs2 = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_64_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_65_rob_idx = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_64_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_imm = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_imm :
    _io_o_issue_packs_1_T_64_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_src1_value = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_src1_value : _io_o_issue_packs_1_T_64_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_65_src2_value = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_src2_value : _io_o_issue_packs_1_T_64_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_65_op1_sel = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_64_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_65_op2_sel = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_64_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_65_alu_sel = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_64_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_65_branch_type = _io_o_issue_packs_1_T_62 ?
    reservation_station_62_io_o_uop_branch_type : _io_o_issue_packs_1_T_64_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_65_mem_type = _io_o_issue_packs_1_T_62 ? reservation_station_62_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_64_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_66_pc = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_pc :
    _io_o_issue_packs_1_T_65_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_66_inst = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_inst :
    _io_o_issue_packs_1_T_65_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_func_code = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_func_code
     : _io_o_issue_packs_1_T_65_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_branch_predict_pack_valid = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_65_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_branch_predict_pack_target = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_65_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_66_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_65_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_branch_predict_pack_select = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_65_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_branch_predict_pack_taken = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_65_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_phy_dst = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_65_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_stale_dst = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_65_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_arch_dst = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_65_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_66_inst_type = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_65_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_regWen = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_regWen :
    _io_o_issue_packs_1_T_65_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_src1_valid = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_65_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_phy_rs1 = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_65_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_arch_rs1 = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_65_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_66_src2_valid = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_65_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_phy_rs2 = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_65_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_arch_rs2 = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_65_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_66_rob_idx = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_65_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_imm = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_imm :
    _io_o_issue_packs_1_T_65_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_src1_value = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_src1_value : _io_o_issue_packs_1_T_65_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_66_src2_value = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_src2_value : _io_o_issue_packs_1_T_65_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_66_op1_sel = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_65_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_66_op2_sel = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_65_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_66_alu_sel = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_65_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_66_branch_type = _io_o_issue_packs_1_T_61 ?
    reservation_station_61_io_o_uop_branch_type : _io_o_issue_packs_1_T_65_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_66_mem_type = _io_o_issue_packs_1_T_61 ? reservation_station_61_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_65_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_67_pc = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_pc :
    _io_o_issue_packs_1_T_66_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_67_inst = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_inst :
    _io_o_issue_packs_1_T_66_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_func_code = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_func_code
     : _io_o_issue_packs_1_T_66_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_branch_predict_pack_valid = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_66_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_branch_predict_pack_target = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_66_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_67_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_66_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_branch_predict_pack_select = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_66_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_branch_predict_pack_taken = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_66_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_phy_dst = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_66_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_stale_dst = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_66_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_arch_dst = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_66_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_67_inst_type = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_66_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_regWen = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_regWen :
    _io_o_issue_packs_1_T_66_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_src1_valid = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_66_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_phy_rs1 = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_66_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_arch_rs1 = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_66_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_67_src2_valid = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_66_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_phy_rs2 = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_66_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_arch_rs2 = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_66_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_67_rob_idx = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_66_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_imm = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_imm :
    _io_o_issue_packs_1_T_66_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_src1_value = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_src1_value : _io_o_issue_packs_1_T_66_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_67_src2_value = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_src2_value : _io_o_issue_packs_1_T_66_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_67_op1_sel = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_66_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_67_op2_sel = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_66_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_67_alu_sel = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_66_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_67_branch_type = _io_o_issue_packs_1_T_60 ?
    reservation_station_60_io_o_uop_branch_type : _io_o_issue_packs_1_T_66_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_67_mem_type = _io_o_issue_packs_1_T_60 ? reservation_station_60_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_66_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_68_pc = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_pc :
    _io_o_issue_packs_1_T_67_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_68_inst = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_inst :
    _io_o_issue_packs_1_T_67_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_func_code = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_func_code
     : _io_o_issue_packs_1_T_67_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_branch_predict_pack_valid = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_67_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_branch_predict_pack_target = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_67_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_68_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_67_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_branch_predict_pack_select = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_67_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_branch_predict_pack_taken = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_67_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_phy_dst = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_67_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_stale_dst = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_67_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_arch_dst = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_67_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_68_inst_type = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_67_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_regWen = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_regWen :
    _io_o_issue_packs_1_T_67_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_src1_valid = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_67_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_phy_rs1 = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_67_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_arch_rs1 = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_67_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_68_src2_valid = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_67_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_phy_rs2 = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_67_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_arch_rs2 = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_67_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_68_rob_idx = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_67_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_imm = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_imm :
    _io_o_issue_packs_1_T_67_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_src1_value = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_src1_value : _io_o_issue_packs_1_T_67_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_68_src2_value = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_src2_value : _io_o_issue_packs_1_T_67_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_68_op1_sel = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_67_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_68_op2_sel = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_67_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_68_alu_sel = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_67_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_68_branch_type = _io_o_issue_packs_1_T_59 ?
    reservation_station_59_io_o_uop_branch_type : _io_o_issue_packs_1_T_67_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_68_mem_type = _io_o_issue_packs_1_T_59 ? reservation_station_59_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_67_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_69_pc = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_pc :
    _io_o_issue_packs_1_T_68_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_69_inst = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_inst :
    _io_o_issue_packs_1_T_68_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_func_code = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_func_code
     : _io_o_issue_packs_1_T_68_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_branch_predict_pack_valid = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_68_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_branch_predict_pack_target = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_68_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_69_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_68_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_branch_predict_pack_select = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_68_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_branch_predict_pack_taken = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_68_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_phy_dst = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_68_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_stale_dst = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_68_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_arch_dst = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_68_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_69_inst_type = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_68_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_regWen = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_regWen :
    _io_o_issue_packs_1_T_68_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_src1_valid = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_68_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_phy_rs1 = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_68_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_arch_rs1 = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_68_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_69_src2_valid = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_68_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_phy_rs2 = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_68_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_arch_rs2 = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_68_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_69_rob_idx = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_68_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_imm = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_imm :
    _io_o_issue_packs_1_T_68_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_src1_value = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_src1_value : _io_o_issue_packs_1_T_68_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_69_src2_value = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_src2_value : _io_o_issue_packs_1_T_68_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_69_op1_sel = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_68_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_69_op2_sel = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_68_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_69_alu_sel = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_68_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_69_branch_type = _io_o_issue_packs_1_T_58 ?
    reservation_station_58_io_o_uop_branch_type : _io_o_issue_packs_1_T_68_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_69_mem_type = _io_o_issue_packs_1_T_58 ? reservation_station_58_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_68_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_70_pc = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_pc :
    _io_o_issue_packs_1_T_69_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_70_inst = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_inst :
    _io_o_issue_packs_1_T_69_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_func_code = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_func_code
     : _io_o_issue_packs_1_T_69_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_branch_predict_pack_valid = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_69_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_branch_predict_pack_target = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_69_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_70_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_69_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_branch_predict_pack_select = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_69_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_branch_predict_pack_taken = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_69_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_phy_dst = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_69_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_stale_dst = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_69_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_arch_dst = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_69_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_70_inst_type = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_69_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_regWen = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_regWen :
    _io_o_issue_packs_1_T_69_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_src1_valid = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_69_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_phy_rs1 = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_69_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_arch_rs1 = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_69_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_70_src2_valid = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_69_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_phy_rs2 = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_69_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_arch_rs2 = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_69_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_70_rob_idx = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_69_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_imm = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_imm :
    _io_o_issue_packs_1_T_69_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_src1_value = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_src1_value : _io_o_issue_packs_1_T_69_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_70_src2_value = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_src2_value : _io_o_issue_packs_1_T_69_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_70_op1_sel = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_69_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_70_op2_sel = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_69_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_70_alu_sel = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_69_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_70_branch_type = _io_o_issue_packs_1_T_57 ?
    reservation_station_57_io_o_uop_branch_type : _io_o_issue_packs_1_T_69_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_70_mem_type = _io_o_issue_packs_1_T_57 ? reservation_station_57_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_69_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_71_pc = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_pc :
    _io_o_issue_packs_1_T_70_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_71_inst = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_inst :
    _io_o_issue_packs_1_T_70_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_func_code = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_func_code
     : _io_o_issue_packs_1_T_70_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_branch_predict_pack_valid = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_70_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_branch_predict_pack_target = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_70_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_71_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_70_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_branch_predict_pack_select = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_70_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_branch_predict_pack_taken = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_70_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_phy_dst = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_70_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_stale_dst = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_70_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_arch_dst = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_70_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_71_inst_type = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_70_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_regWen = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_regWen :
    _io_o_issue_packs_1_T_70_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_src1_valid = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_70_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_phy_rs1 = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_70_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_arch_rs1 = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_70_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_71_src2_valid = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_70_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_phy_rs2 = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_70_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_arch_rs2 = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_70_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_71_rob_idx = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_70_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_imm = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_imm :
    _io_o_issue_packs_1_T_70_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_src1_value = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_src1_value : _io_o_issue_packs_1_T_70_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_71_src2_value = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_src2_value : _io_o_issue_packs_1_T_70_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_71_op1_sel = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_70_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_71_op2_sel = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_70_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_71_alu_sel = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_70_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_71_branch_type = _io_o_issue_packs_1_T_56 ?
    reservation_station_56_io_o_uop_branch_type : _io_o_issue_packs_1_T_70_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_71_mem_type = _io_o_issue_packs_1_T_56 ? reservation_station_56_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_70_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_72_pc = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_pc :
    _io_o_issue_packs_1_T_71_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_72_inst = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_inst :
    _io_o_issue_packs_1_T_71_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_func_code = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_func_code
     : _io_o_issue_packs_1_T_71_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_branch_predict_pack_valid = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_71_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_branch_predict_pack_target = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_71_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_72_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_71_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_branch_predict_pack_select = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_71_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_branch_predict_pack_taken = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_71_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_phy_dst = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_71_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_stale_dst = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_71_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_arch_dst = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_71_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_72_inst_type = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_71_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_regWen = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_regWen :
    _io_o_issue_packs_1_T_71_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_src1_valid = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_71_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_phy_rs1 = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_71_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_arch_rs1 = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_71_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_72_src2_valid = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_71_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_phy_rs2 = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_71_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_arch_rs2 = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_71_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_72_rob_idx = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_71_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_imm = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_imm :
    _io_o_issue_packs_1_T_71_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_src1_value = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_src1_value : _io_o_issue_packs_1_T_71_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_72_src2_value = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_src2_value : _io_o_issue_packs_1_T_71_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_72_op1_sel = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_71_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_72_op2_sel = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_71_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_72_alu_sel = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_71_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_72_branch_type = _io_o_issue_packs_1_T_55 ?
    reservation_station_55_io_o_uop_branch_type : _io_o_issue_packs_1_T_71_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_72_mem_type = _io_o_issue_packs_1_T_55 ? reservation_station_55_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_71_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_73_pc = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_pc :
    _io_o_issue_packs_1_T_72_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_73_inst = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_inst :
    _io_o_issue_packs_1_T_72_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_func_code = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_func_code
     : _io_o_issue_packs_1_T_72_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_branch_predict_pack_valid = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_72_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_branch_predict_pack_target = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_72_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_73_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_72_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_branch_predict_pack_select = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_72_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_branch_predict_pack_taken = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_72_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_phy_dst = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_72_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_stale_dst = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_72_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_arch_dst = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_72_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_73_inst_type = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_72_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_regWen = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_regWen :
    _io_o_issue_packs_1_T_72_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_src1_valid = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_72_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_phy_rs1 = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_72_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_arch_rs1 = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_72_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_73_src2_valid = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_72_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_phy_rs2 = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_72_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_arch_rs2 = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_72_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_73_rob_idx = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_72_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_imm = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_imm :
    _io_o_issue_packs_1_T_72_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_src1_value = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_src1_value : _io_o_issue_packs_1_T_72_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_73_src2_value = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_src2_value : _io_o_issue_packs_1_T_72_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_73_op1_sel = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_72_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_73_op2_sel = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_72_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_73_alu_sel = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_72_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_73_branch_type = _io_o_issue_packs_1_T_54 ?
    reservation_station_54_io_o_uop_branch_type : _io_o_issue_packs_1_T_72_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_73_mem_type = _io_o_issue_packs_1_T_54 ? reservation_station_54_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_72_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_74_pc = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_pc :
    _io_o_issue_packs_1_T_73_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_74_inst = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_inst :
    _io_o_issue_packs_1_T_73_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_func_code = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_func_code
     : _io_o_issue_packs_1_T_73_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_branch_predict_pack_valid = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_73_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_branch_predict_pack_target = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_73_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_74_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_73_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_branch_predict_pack_select = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_73_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_branch_predict_pack_taken = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_73_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_phy_dst = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_73_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_stale_dst = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_73_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_arch_dst = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_73_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_74_inst_type = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_73_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_regWen = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_regWen :
    _io_o_issue_packs_1_T_73_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_src1_valid = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_73_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_phy_rs1 = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_73_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_arch_rs1 = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_73_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_74_src2_valid = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_73_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_phy_rs2 = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_73_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_arch_rs2 = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_73_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_74_rob_idx = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_73_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_imm = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_imm :
    _io_o_issue_packs_1_T_73_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_src1_value = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_src1_value : _io_o_issue_packs_1_T_73_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_74_src2_value = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_src2_value : _io_o_issue_packs_1_T_73_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_74_op1_sel = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_73_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_74_op2_sel = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_73_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_74_alu_sel = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_73_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_74_branch_type = _io_o_issue_packs_1_T_53 ?
    reservation_station_53_io_o_uop_branch_type : _io_o_issue_packs_1_T_73_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_74_mem_type = _io_o_issue_packs_1_T_53 ? reservation_station_53_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_73_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_75_pc = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_pc :
    _io_o_issue_packs_1_T_74_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_75_inst = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_inst :
    _io_o_issue_packs_1_T_74_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_func_code = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_func_code
     : _io_o_issue_packs_1_T_74_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_branch_predict_pack_valid = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_74_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_branch_predict_pack_target = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_74_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_75_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_74_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_branch_predict_pack_select = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_74_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_branch_predict_pack_taken = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_74_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_phy_dst = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_74_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_stale_dst = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_74_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_arch_dst = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_74_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_75_inst_type = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_74_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_regWen = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_regWen :
    _io_o_issue_packs_1_T_74_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_src1_valid = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_74_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_phy_rs1 = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_74_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_arch_rs1 = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_74_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_75_src2_valid = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_74_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_phy_rs2 = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_74_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_arch_rs2 = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_74_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_75_rob_idx = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_74_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_imm = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_imm :
    _io_o_issue_packs_1_T_74_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_src1_value = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_src1_value : _io_o_issue_packs_1_T_74_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_75_src2_value = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_src2_value : _io_o_issue_packs_1_T_74_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_75_op1_sel = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_74_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_75_op2_sel = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_74_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_75_alu_sel = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_74_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_75_branch_type = _io_o_issue_packs_1_T_52 ?
    reservation_station_52_io_o_uop_branch_type : _io_o_issue_packs_1_T_74_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_75_mem_type = _io_o_issue_packs_1_T_52 ? reservation_station_52_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_74_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_76_pc = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_pc :
    _io_o_issue_packs_1_T_75_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_76_inst = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_inst :
    _io_o_issue_packs_1_T_75_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_func_code = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_func_code
     : _io_o_issue_packs_1_T_75_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_branch_predict_pack_valid = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_75_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_branch_predict_pack_target = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_75_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_76_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_75_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_branch_predict_pack_select = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_75_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_branch_predict_pack_taken = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_75_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_phy_dst = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_75_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_stale_dst = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_75_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_arch_dst = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_75_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_76_inst_type = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_75_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_regWen = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_regWen :
    _io_o_issue_packs_1_T_75_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_src1_valid = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_75_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_phy_rs1 = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_75_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_arch_rs1 = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_75_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_76_src2_valid = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_75_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_phy_rs2 = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_75_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_arch_rs2 = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_75_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_76_rob_idx = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_75_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_imm = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_imm :
    _io_o_issue_packs_1_T_75_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_src1_value = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_src1_value : _io_o_issue_packs_1_T_75_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_76_src2_value = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_src2_value : _io_o_issue_packs_1_T_75_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_76_op1_sel = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_75_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_76_op2_sel = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_75_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_76_alu_sel = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_75_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_76_branch_type = _io_o_issue_packs_1_T_51 ?
    reservation_station_51_io_o_uop_branch_type : _io_o_issue_packs_1_T_75_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_76_mem_type = _io_o_issue_packs_1_T_51 ? reservation_station_51_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_75_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_77_pc = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_pc :
    _io_o_issue_packs_1_T_76_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_77_inst = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_inst :
    _io_o_issue_packs_1_T_76_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_func_code = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_func_code
     : _io_o_issue_packs_1_T_76_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_branch_predict_pack_valid = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_76_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_branch_predict_pack_target = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_76_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_77_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_76_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_branch_predict_pack_select = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_76_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_branch_predict_pack_taken = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_76_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_phy_dst = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_76_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_stale_dst = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_76_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_arch_dst = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_76_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_77_inst_type = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_76_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_regWen = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_regWen :
    _io_o_issue_packs_1_T_76_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_src1_valid = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_76_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_phy_rs1 = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_76_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_arch_rs1 = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_76_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_77_src2_valid = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_76_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_phy_rs2 = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_76_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_arch_rs2 = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_76_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_77_rob_idx = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_76_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_imm = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_imm :
    _io_o_issue_packs_1_T_76_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_src1_value = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_src1_value : _io_o_issue_packs_1_T_76_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_77_src2_value = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_src2_value : _io_o_issue_packs_1_T_76_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_77_op1_sel = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_76_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_77_op2_sel = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_76_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_77_alu_sel = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_76_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_77_branch_type = _io_o_issue_packs_1_T_50 ?
    reservation_station_50_io_o_uop_branch_type : _io_o_issue_packs_1_T_76_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_77_mem_type = _io_o_issue_packs_1_T_50 ? reservation_station_50_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_76_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_78_pc = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_pc :
    _io_o_issue_packs_1_T_77_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_78_inst = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_inst :
    _io_o_issue_packs_1_T_77_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_func_code = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_func_code
     : _io_o_issue_packs_1_T_77_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_branch_predict_pack_valid = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_77_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_branch_predict_pack_target = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_77_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_78_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_77_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_branch_predict_pack_select = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_77_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_branch_predict_pack_taken = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_77_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_phy_dst = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_77_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_stale_dst = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_77_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_arch_dst = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_77_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_78_inst_type = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_77_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_regWen = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_regWen :
    _io_o_issue_packs_1_T_77_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_src1_valid = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_77_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_phy_rs1 = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_77_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_arch_rs1 = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_77_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_78_src2_valid = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_77_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_phy_rs2 = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_77_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_arch_rs2 = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_77_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_78_rob_idx = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_77_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_imm = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_imm :
    _io_o_issue_packs_1_T_77_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_src1_value = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_src1_value : _io_o_issue_packs_1_T_77_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_78_src2_value = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_src2_value : _io_o_issue_packs_1_T_77_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_78_op1_sel = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_77_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_78_op2_sel = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_77_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_78_alu_sel = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_77_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_78_branch_type = _io_o_issue_packs_1_T_49 ?
    reservation_station_49_io_o_uop_branch_type : _io_o_issue_packs_1_T_77_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_78_mem_type = _io_o_issue_packs_1_T_49 ? reservation_station_49_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_77_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_79_pc = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_pc :
    _io_o_issue_packs_1_T_78_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_79_inst = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_inst :
    _io_o_issue_packs_1_T_78_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_func_code = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_func_code
     : _io_o_issue_packs_1_T_78_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_branch_predict_pack_valid = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_78_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_branch_predict_pack_target = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_78_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_79_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_78_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_branch_predict_pack_select = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_78_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_branch_predict_pack_taken = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_78_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_phy_dst = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_78_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_stale_dst = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_78_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_arch_dst = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_78_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_79_inst_type = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_78_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_regWen = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_regWen :
    _io_o_issue_packs_1_T_78_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_src1_valid = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_78_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_phy_rs1 = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_78_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_arch_rs1 = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_78_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_79_src2_valid = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_78_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_phy_rs2 = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_78_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_arch_rs2 = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_78_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_79_rob_idx = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_78_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_imm = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_imm :
    _io_o_issue_packs_1_T_78_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_src1_value = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_src1_value : _io_o_issue_packs_1_T_78_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_79_src2_value = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_src2_value : _io_o_issue_packs_1_T_78_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_79_op1_sel = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_78_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_79_op2_sel = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_78_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_79_alu_sel = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_78_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_79_branch_type = _io_o_issue_packs_1_T_48 ?
    reservation_station_48_io_o_uop_branch_type : _io_o_issue_packs_1_T_78_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_79_mem_type = _io_o_issue_packs_1_T_48 ? reservation_station_48_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_78_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_80_pc = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_pc :
    _io_o_issue_packs_1_T_79_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_80_inst = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_inst :
    _io_o_issue_packs_1_T_79_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_func_code = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_func_code
     : _io_o_issue_packs_1_T_79_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_branch_predict_pack_valid = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_79_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_branch_predict_pack_target = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_79_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_80_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_79_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_branch_predict_pack_select = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_79_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_branch_predict_pack_taken = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_79_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_phy_dst = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_79_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_stale_dst = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_79_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_arch_dst = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_79_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_80_inst_type = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_79_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_regWen = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_regWen :
    _io_o_issue_packs_1_T_79_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_src1_valid = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_79_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_phy_rs1 = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_79_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_arch_rs1 = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_79_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_80_src2_valid = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_79_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_phy_rs2 = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_79_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_arch_rs2 = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_79_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_80_rob_idx = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_79_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_imm = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_imm :
    _io_o_issue_packs_1_T_79_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_src1_value = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_src1_value : _io_o_issue_packs_1_T_79_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_80_src2_value = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_src2_value : _io_o_issue_packs_1_T_79_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_80_op1_sel = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_79_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_80_op2_sel = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_79_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_80_alu_sel = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_79_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_80_branch_type = _io_o_issue_packs_1_T_47 ?
    reservation_station_47_io_o_uop_branch_type : _io_o_issue_packs_1_T_79_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_80_mem_type = _io_o_issue_packs_1_T_47 ? reservation_station_47_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_79_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_81_pc = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_pc :
    _io_o_issue_packs_1_T_80_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_81_inst = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_inst :
    _io_o_issue_packs_1_T_80_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_func_code = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_func_code
     : _io_o_issue_packs_1_T_80_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_branch_predict_pack_valid = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_80_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_branch_predict_pack_target = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_80_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_81_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_80_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_branch_predict_pack_select = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_80_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_branch_predict_pack_taken = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_80_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_phy_dst = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_80_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_stale_dst = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_80_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_arch_dst = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_80_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_81_inst_type = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_80_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_regWen = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_regWen :
    _io_o_issue_packs_1_T_80_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_src1_valid = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_80_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_phy_rs1 = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_80_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_arch_rs1 = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_80_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_81_src2_valid = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_80_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_phy_rs2 = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_80_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_arch_rs2 = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_80_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_81_rob_idx = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_80_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_imm = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_imm :
    _io_o_issue_packs_1_T_80_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_src1_value = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_src1_value : _io_o_issue_packs_1_T_80_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_81_src2_value = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_src2_value : _io_o_issue_packs_1_T_80_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_81_op1_sel = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_80_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_81_op2_sel = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_80_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_81_alu_sel = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_80_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_81_branch_type = _io_o_issue_packs_1_T_46 ?
    reservation_station_46_io_o_uop_branch_type : _io_o_issue_packs_1_T_80_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_81_mem_type = _io_o_issue_packs_1_T_46 ? reservation_station_46_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_80_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_82_pc = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_pc :
    _io_o_issue_packs_1_T_81_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_82_inst = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_inst :
    _io_o_issue_packs_1_T_81_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_func_code = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_func_code
     : _io_o_issue_packs_1_T_81_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_branch_predict_pack_valid = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_81_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_branch_predict_pack_target = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_81_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_82_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_81_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_branch_predict_pack_select = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_81_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_branch_predict_pack_taken = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_81_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_phy_dst = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_81_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_stale_dst = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_81_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_arch_dst = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_81_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_82_inst_type = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_81_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_regWen = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_regWen :
    _io_o_issue_packs_1_T_81_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_src1_valid = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_81_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_phy_rs1 = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_81_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_arch_rs1 = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_81_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_82_src2_valid = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_81_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_phy_rs2 = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_81_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_arch_rs2 = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_81_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_82_rob_idx = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_81_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_imm = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_imm :
    _io_o_issue_packs_1_T_81_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_src1_value = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_src1_value : _io_o_issue_packs_1_T_81_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_82_src2_value = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_src2_value : _io_o_issue_packs_1_T_81_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_82_op1_sel = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_81_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_82_op2_sel = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_81_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_82_alu_sel = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_81_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_82_branch_type = _io_o_issue_packs_1_T_45 ?
    reservation_station_45_io_o_uop_branch_type : _io_o_issue_packs_1_T_81_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_82_mem_type = _io_o_issue_packs_1_T_45 ? reservation_station_45_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_81_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_83_pc = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_pc :
    _io_o_issue_packs_1_T_82_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_83_inst = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_inst :
    _io_o_issue_packs_1_T_82_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_func_code = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_func_code
     : _io_o_issue_packs_1_T_82_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_branch_predict_pack_valid = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_82_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_branch_predict_pack_target = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_82_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_83_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_82_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_branch_predict_pack_select = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_82_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_branch_predict_pack_taken = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_82_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_phy_dst = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_82_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_stale_dst = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_82_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_arch_dst = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_82_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_83_inst_type = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_82_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_regWen = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_regWen :
    _io_o_issue_packs_1_T_82_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_src1_valid = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_82_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_phy_rs1 = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_82_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_arch_rs1 = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_82_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_83_src2_valid = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_82_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_phy_rs2 = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_82_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_arch_rs2 = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_82_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_83_rob_idx = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_82_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_imm = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_imm :
    _io_o_issue_packs_1_T_82_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_src1_value = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_src1_value : _io_o_issue_packs_1_T_82_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_83_src2_value = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_src2_value : _io_o_issue_packs_1_T_82_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_83_op1_sel = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_82_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_83_op2_sel = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_82_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_83_alu_sel = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_82_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_83_branch_type = _io_o_issue_packs_1_T_44 ?
    reservation_station_44_io_o_uop_branch_type : _io_o_issue_packs_1_T_82_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_83_mem_type = _io_o_issue_packs_1_T_44 ? reservation_station_44_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_82_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_84_pc = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_pc :
    _io_o_issue_packs_1_T_83_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_84_inst = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_inst :
    _io_o_issue_packs_1_T_83_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_func_code = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_func_code
     : _io_o_issue_packs_1_T_83_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_branch_predict_pack_valid = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_83_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_branch_predict_pack_target = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_83_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_84_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_83_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_branch_predict_pack_select = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_83_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_branch_predict_pack_taken = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_83_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_phy_dst = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_83_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_stale_dst = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_83_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_arch_dst = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_83_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_84_inst_type = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_83_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_regWen = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_regWen :
    _io_o_issue_packs_1_T_83_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_src1_valid = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_83_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_phy_rs1 = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_83_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_arch_rs1 = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_83_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_84_src2_valid = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_83_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_phy_rs2 = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_83_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_arch_rs2 = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_83_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_84_rob_idx = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_83_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_imm = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_imm :
    _io_o_issue_packs_1_T_83_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_src1_value = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_src1_value : _io_o_issue_packs_1_T_83_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_84_src2_value = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_src2_value : _io_o_issue_packs_1_T_83_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_84_op1_sel = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_83_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_84_op2_sel = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_83_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_84_alu_sel = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_83_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_84_branch_type = _io_o_issue_packs_1_T_43 ?
    reservation_station_43_io_o_uop_branch_type : _io_o_issue_packs_1_T_83_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_84_mem_type = _io_o_issue_packs_1_T_43 ? reservation_station_43_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_83_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_85_pc = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_pc :
    _io_o_issue_packs_1_T_84_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_85_inst = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_inst :
    _io_o_issue_packs_1_T_84_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_func_code = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_func_code
     : _io_o_issue_packs_1_T_84_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_branch_predict_pack_valid = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_84_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_branch_predict_pack_target = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_84_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_85_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_84_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_branch_predict_pack_select = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_84_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_branch_predict_pack_taken = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_84_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_phy_dst = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_84_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_stale_dst = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_84_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_arch_dst = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_84_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_85_inst_type = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_84_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_regWen = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_regWen :
    _io_o_issue_packs_1_T_84_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_src1_valid = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_84_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_phy_rs1 = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_84_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_arch_rs1 = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_84_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_85_src2_valid = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_84_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_phy_rs2 = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_84_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_arch_rs2 = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_84_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_85_rob_idx = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_84_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_imm = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_imm :
    _io_o_issue_packs_1_T_84_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_src1_value = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_src1_value : _io_o_issue_packs_1_T_84_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_85_src2_value = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_src2_value : _io_o_issue_packs_1_T_84_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_85_op1_sel = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_84_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_85_op2_sel = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_84_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_85_alu_sel = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_84_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_85_branch_type = _io_o_issue_packs_1_T_42 ?
    reservation_station_42_io_o_uop_branch_type : _io_o_issue_packs_1_T_84_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_85_mem_type = _io_o_issue_packs_1_T_42 ? reservation_station_42_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_84_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_86_pc = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_pc :
    _io_o_issue_packs_1_T_85_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_86_inst = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_inst :
    _io_o_issue_packs_1_T_85_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_func_code = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_func_code
     : _io_o_issue_packs_1_T_85_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_branch_predict_pack_valid = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_85_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_branch_predict_pack_target = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_85_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_86_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_85_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_branch_predict_pack_select = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_85_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_branch_predict_pack_taken = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_85_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_phy_dst = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_85_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_stale_dst = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_85_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_arch_dst = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_85_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_86_inst_type = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_85_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_regWen = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_regWen :
    _io_o_issue_packs_1_T_85_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_src1_valid = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_85_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_phy_rs1 = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_85_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_arch_rs1 = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_85_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_86_src2_valid = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_85_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_phy_rs2 = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_85_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_arch_rs2 = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_85_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_86_rob_idx = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_85_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_imm = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_imm :
    _io_o_issue_packs_1_T_85_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_src1_value = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_src1_value : _io_o_issue_packs_1_T_85_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_86_src2_value = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_src2_value : _io_o_issue_packs_1_T_85_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_86_op1_sel = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_85_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_86_op2_sel = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_85_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_86_alu_sel = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_85_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_86_branch_type = _io_o_issue_packs_1_T_41 ?
    reservation_station_41_io_o_uop_branch_type : _io_o_issue_packs_1_T_85_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_86_mem_type = _io_o_issue_packs_1_T_41 ? reservation_station_41_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_85_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_87_pc = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_pc :
    _io_o_issue_packs_1_T_86_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_87_inst = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_inst :
    _io_o_issue_packs_1_T_86_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_func_code = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_func_code
     : _io_o_issue_packs_1_T_86_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_branch_predict_pack_valid = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_86_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_branch_predict_pack_target = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_86_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_87_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_86_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_branch_predict_pack_select = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_86_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_branch_predict_pack_taken = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_86_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_phy_dst = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_86_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_stale_dst = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_86_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_arch_dst = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_86_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_87_inst_type = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_86_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_regWen = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_regWen :
    _io_o_issue_packs_1_T_86_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_src1_valid = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_86_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_phy_rs1 = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_86_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_arch_rs1 = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_86_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_87_src2_valid = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_86_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_phy_rs2 = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_86_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_arch_rs2 = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_86_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_87_rob_idx = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_86_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_imm = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_imm :
    _io_o_issue_packs_1_T_86_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_src1_value = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_src1_value : _io_o_issue_packs_1_T_86_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_87_src2_value = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_src2_value : _io_o_issue_packs_1_T_86_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_87_op1_sel = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_86_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_87_op2_sel = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_86_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_87_alu_sel = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_86_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_87_branch_type = _io_o_issue_packs_1_T_40 ?
    reservation_station_40_io_o_uop_branch_type : _io_o_issue_packs_1_T_86_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_87_mem_type = _io_o_issue_packs_1_T_40 ? reservation_station_40_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_86_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_88_pc = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_pc :
    _io_o_issue_packs_1_T_87_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_88_inst = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_inst :
    _io_o_issue_packs_1_T_87_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_func_code = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_func_code
     : _io_o_issue_packs_1_T_87_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_branch_predict_pack_valid = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_87_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_branch_predict_pack_target = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_87_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_88_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_87_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_branch_predict_pack_select = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_87_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_branch_predict_pack_taken = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_87_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_phy_dst = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_87_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_stale_dst = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_87_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_arch_dst = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_87_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_88_inst_type = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_87_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_regWen = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_regWen :
    _io_o_issue_packs_1_T_87_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_src1_valid = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_87_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_phy_rs1 = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_87_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_arch_rs1 = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_87_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_88_src2_valid = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_87_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_phy_rs2 = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_87_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_arch_rs2 = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_87_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_88_rob_idx = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_87_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_imm = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_imm :
    _io_o_issue_packs_1_T_87_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_src1_value = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_src1_value : _io_o_issue_packs_1_T_87_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_88_src2_value = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_src2_value : _io_o_issue_packs_1_T_87_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_88_op1_sel = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_87_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_88_op2_sel = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_87_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_88_alu_sel = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_87_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_88_branch_type = _io_o_issue_packs_1_T_39 ?
    reservation_station_39_io_o_uop_branch_type : _io_o_issue_packs_1_T_87_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_88_mem_type = _io_o_issue_packs_1_T_39 ? reservation_station_39_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_87_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_89_pc = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_pc :
    _io_o_issue_packs_1_T_88_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_89_inst = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_inst :
    _io_o_issue_packs_1_T_88_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_func_code = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_func_code
     : _io_o_issue_packs_1_T_88_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_branch_predict_pack_valid = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_88_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_branch_predict_pack_target = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_88_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_89_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_88_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_branch_predict_pack_select = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_88_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_branch_predict_pack_taken = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_88_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_phy_dst = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_88_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_stale_dst = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_88_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_arch_dst = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_88_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_89_inst_type = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_88_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_regWen = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_regWen :
    _io_o_issue_packs_1_T_88_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_src1_valid = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_88_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_phy_rs1 = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_88_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_arch_rs1 = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_88_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_89_src2_valid = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_88_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_phy_rs2 = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_88_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_arch_rs2 = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_88_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_89_rob_idx = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_88_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_imm = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_imm :
    _io_o_issue_packs_1_T_88_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_src1_value = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_src1_value : _io_o_issue_packs_1_T_88_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_89_src2_value = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_src2_value : _io_o_issue_packs_1_T_88_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_89_op1_sel = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_88_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_89_op2_sel = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_88_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_89_alu_sel = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_88_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_89_branch_type = _io_o_issue_packs_1_T_38 ?
    reservation_station_38_io_o_uop_branch_type : _io_o_issue_packs_1_T_88_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_89_mem_type = _io_o_issue_packs_1_T_38 ? reservation_station_38_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_88_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_90_pc = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_pc :
    _io_o_issue_packs_1_T_89_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_90_inst = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_inst :
    _io_o_issue_packs_1_T_89_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_func_code = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_func_code
     : _io_o_issue_packs_1_T_89_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_branch_predict_pack_valid = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_89_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_branch_predict_pack_target = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_89_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_90_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_89_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_branch_predict_pack_select = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_89_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_branch_predict_pack_taken = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_89_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_phy_dst = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_89_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_stale_dst = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_89_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_arch_dst = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_89_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_90_inst_type = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_89_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_regWen = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_regWen :
    _io_o_issue_packs_1_T_89_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_src1_valid = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_89_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_phy_rs1 = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_89_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_arch_rs1 = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_89_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_90_src2_valid = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_89_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_phy_rs2 = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_89_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_arch_rs2 = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_89_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_90_rob_idx = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_89_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_imm = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_imm :
    _io_o_issue_packs_1_T_89_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_src1_value = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_src1_value : _io_o_issue_packs_1_T_89_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_90_src2_value = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_src2_value : _io_o_issue_packs_1_T_89_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_90_op1_sel = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_89_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_90_op2_sel = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_89_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_90_alu_sel = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_89_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_90_branch_type = _io_o_issue_packs_1_T_37 ?
    reservation_station_37_io_o_uop_branch_type : _io_o_issue_packs_1_T_89_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_90_mem_type = _io_o_issue_packs_1_T_37 ? reservation_station_37_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_89_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_91_pc = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_pc :
    _io_o_issue_packs_1_T_90_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_91_inst = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_inst :
    _io_o_issue_packs_1_T_90_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_func_code = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_func_code
     : _io_o_issue_packs_1_T_90_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_branch_predict_pack_valid = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_90_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_branch_predict_pack_target = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_90_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_91_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_90_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_branch_predict_pack_select = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_90_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_branch_predict_pack_taken = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_90_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_phy_dst = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_90_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_stale_dst = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_90_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_arch_dst = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_90_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_91_inst_type = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_90_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_regWen = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_regWen :
    _io_o_issue_packs_1_T_90_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_src1_valid = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_90_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_phy_rs1 = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_90_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_arch_rs1 = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_90_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_91_src2_valid = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_90_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_phy_rs2 = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_90_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_arch_rs2 = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_90_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_91_rob_idx = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_90_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_imm = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_imm :
    _io_o_issue_packs_1_T_90_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_src1_value = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_src1_value : _io_o_issue_packs_1_T_90_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_91_src2_value = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_src2_value : _io_o_issue_packs_1_T_90_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_91_op1_sel = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_90_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_91_op2_sel = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_90_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_91_alu_sel = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_90_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_91_branch_type = _io_o_issue_packs_1_T_36 ?
    reservation_station_36_io_o_uop_branch_type : _io_o_issue_packs_1_T_90_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_91_mem_type = _io_o_issue_packs_1_T_36 ? reservation_station_36_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_90_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_92_pc = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_pc :
    _io_o_issue_packs_1_T_91_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_92_inst = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_inst :
    _io_o_issue_packs_1_T_91_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_func_code = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_func_code
     : _io_o_issue_packs_1_T_91_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_branch_predict_pack_valid = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_91_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_branch_predict_pack_target = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_91_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_92_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_91_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_branch_predict_pack_select = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_91_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_branch_predict_pack_taken = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_91_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_phy_dst = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_91_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_stale_dst = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_91_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_arch_dst = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_91_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_92_inst_type = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_91_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_regWen = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_regWen :
    _io_o_issue_packs_1_T_91_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_src1_valid = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_91_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_phy_rs1 = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_91_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_arch_rs1 = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_91_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_92_src2_valid = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_91_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_phy_rs2 = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_91_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_arch_rs2 = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_91_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_92_rob_idx = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_91_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_imm = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_imm :
    _io_o_issue_packs_1_T_91_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_src1_value = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_src1_value : _io_o_issue_packs_1_T_91_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_92_src2_value = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_src2_value : _io_o_issue_packs_1_T_91_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_92_op1_sel = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_91_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_92_op2_sel = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_91_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_92_alu_sel = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_91_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_92_branch_type = _io_o_issue_packs_1_T_35 ?
    reservation_station_35_io_o_uop_branch_type : _io_o_issue_packs_1_T_91_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_92_mem_type = _io_o_issue_packs_1_T_35 ? reservation_station_35_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_91_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_93_pc = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_pc :
    _io_o_issue_packs_1_T_92_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_93_inst = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_inst :
    _io_o_issue_packs_1_T_92_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_func_code = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_func_code
     : _io_o_issue_packs_1_T_92_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_branch_predict_pack_valid = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_92_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_branch_predict_pack_target = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_92_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_93_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_92_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_branch_predict_pack_select = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_92_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_branch_predict_pack_taken = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_92_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_phy_dst = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_92_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_stale_dst = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_92_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_arch_dst = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_92_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_93_inst_type = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_92_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_regWen = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_regWen :
    _io_o_issue_packs_1_T_92_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_src1_valid = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_92_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_phy_rs1 = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_92_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_arch_rs1 = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_92_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_93_src2_valid = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_92_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_phy_rs2 = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_92_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_arch_rs2 = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_92_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_93_rob_idx = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_92_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_imm = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_imm :
    _io_o_issue_packs_1_T_92_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_src1_value = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_src1_value : _io_o_issue_packs_1_T_92_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_93_src2_value = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_src2_value : _io_o_issue_packs_1_T_92_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_93_op1_sel = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_92_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_93_op2_sel = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_92_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_93_alu_sel = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_92_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_93_branch_type = _io_o_issue_packs_1_T_34 ?
    reservation_station_34_io_o_uop_branch_type : _io_o_issue_packs_1_T_92_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_93_mem_type = _io_o_issue_packs_1_T_34 ? reservation_station_34_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_92_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_94_pc = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_pc :
    _io_o_issue_packs_1_T_93_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_94_inst = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_inst :
    _io_o_issue_packs_1_T_93_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_func_code = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_func_code
     : _io_o_issue_packs_1_T_93_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_branch_predict_pack_valid = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_93_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_branch_predict_pack_target = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_93_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_94_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_93_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_branch_predict_pack_select = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_93_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_branch_predict_pack_taken = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_93_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_phy_dst = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_93_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_stale_dst = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_93_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_arch_dst = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_93_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_94_inst_type = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_93_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_regWen = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_regWen :
    _io_o_issue_packs_1_T_93_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_src1_valid = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_93_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_phy_rs1 = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_93_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_arch_rs1 = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_93_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_94_src2_valid = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_93_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_phy_rs2 = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_93_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_arch_rs2 = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_93_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_94_rob_idx = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_93_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_imm = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_imm :
    _io_o_issue_packs_1_T_93_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_src1_value = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_src1_value : _io_o_issue_packs_1_T_93_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_94_src2_value = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_src2_value : _io_o_issue_packs_1_T_93_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_94_op1_sel = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_93_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_94_op2_sel = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_93_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_94_alu_sel = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_93_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_94_branch_type = _io_o_issue_packs_1_T_33 ?
    reservation_station_33_io_o_uop_branch_type : _io_o_issue_packs_1_T_93_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_94_mem_type = _io_o_issue_packs_1_T_33 ? reservation_station_33_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_93_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_95_pc = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_pc :
    _io_o_issue_packs_1_T_94_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_95_inst = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_inst :
    _io_o_issue_packs_1_T_94_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_func_code = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_func_code
     : _io_o_issue_packs_1_T_94_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_branch_predict_pack_valid = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_94_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_branch_predict_pack_target = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_94_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_95_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_94_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_branch_predict_pack_select = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_94_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_branch_predict_pack_taken = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_94_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_phy_dst = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_94_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_stale_dst = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_94_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_arch_dst = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_94_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_95_inst_type = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_94_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_regWen = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_regWen :
    _io_o_issue_packs_1_T_94_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_src1_valid = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_94_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_phy_rs1 = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_94_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_arch_rs1 = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_94_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_95_src2_valid = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_94_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_phy_rs2 = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_94_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_arch_rs2 = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_94_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_95_rob_idx = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_94_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_imm = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_imm :
    _io_o_issue_packs_1_T_94_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_src1_value = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_src1_value : _io_o_issue_packs_1_T_94_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_95_src2_value = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_src2_value : _io_o_issue_packs_1_T_94_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_95_op1_sel = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_94_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_95_op2_sel = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_94_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_95_alu_sel = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_94_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_95_branch_type = _io_o_issue_packs_1_T_32 ?
    reservation_station_32_io_o_uop_branch_type : _io_o_issue_packs_1_T_94_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_95_mem_type = _io_o_issue_packs_1_T_32 ? reservation_station_32_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_94_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_96_pc = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_pc :
    _io_o_issue_packs_1_T_95_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_96_inst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_inst :
    _io_o_issue_packs_1_T_95_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_func_code = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_func_code
     : _io_o_issue_packs_1_T_95_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_branch_predict_pack_valid = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_95_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_branch_predict_pack_target = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_95_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_96_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_95_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_branch_predict_pack_select = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_95_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_branch_predict_pack_taken = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_95_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_phy_dst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_95_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_stale_dst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_95_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_arch_dst = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_95_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_96_inst_type = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_95_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_regWen = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_regWen :
    _io_o_issue_packs_1_T_95_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_src1_valid = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_95_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_phy_rs1 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_95_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_arch_rs1 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_95_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_96_src2_valid = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_95_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_phy_rs2 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_95_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_arch_rs2 = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_95_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_96_rob_idx = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_95_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_imm = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_imm :
    _io_o_issue_packs_1_T_95_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_src1_value = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_src1_value : _io_o_issue_packs_1_T_95_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_96_src2_value = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_src2_value : _io_o_issue_packs_1_T_95_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_96_op1_sel = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_95_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_96_op2_sel = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_95_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_96_alu_sel = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_95_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_96_branch_type = _io_o_issue_packs_1_T_31 ?
    reservation_station_31_io_o_uop_branch_type : _io_o_issue_packs_1_T_95_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_96_mem_type = _io_o_issue_packs_1_T_31 ? reservation_station_31_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_95_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_97_pc = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_pc :
    _io_o_issue_packs_1_T_96_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_97_inst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_inst :
    _io_o_issue_packs_1_T_96_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_func_code = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_func_code
     : _io_o_issue_packs_1_T_96_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_branch_predict_pack_valid = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_96_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_branch_predict_pack_target = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_96_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_97_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_96_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_branch_predict_pack_select = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_96_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_branch_predict_pack_taken = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_96_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_phy_dst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_96_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_stale_dst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_96_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_arch_dst = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_96_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_97_inst_type = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_96_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_regWen = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_regWen :
    _io_o_issue_packs_1_T_96_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_src1_valid = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_96_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_phy_rs1 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_96_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_arch_rs1 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_96_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_97_src2_valid = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_96_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_phy_rs2 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_96_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_arch_rs2 = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_96_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_97_rob_idx = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_96_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_imm = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_imm :
    _io_o_issue_packs_1_T_96_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_src1_value = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_src1_value : _io_o_issue_packs_1_T_96_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_97_src2_value = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_src2_value : _io_o_issue_packs_1_T_96_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_97_op1_sel = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_96_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_97_op2_sel = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_96_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_97_alu_sel = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_96_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_97_branch_type = _io_o_issue_packs_1_T_30 ?
    reservation_station_30_io_o_uop_branch_type : _io_o_issue_packs_1_T_96_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_97_mem_type = _io_o_issue_packs_1_T_30 ? reservation_station_30_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_96_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_98_pc = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_pc :
    _io_o_issue_packs_1_T_97_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_98_inst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_inst :
    _io_o_issue_packs_1_T_97_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_func_code = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_func_code
     : _io_o_issue_packs_1_T_97_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_branch_predict_pack_valid = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_97_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_branch_predict_pack_target = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_97_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_98_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_97_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_branch_predict_pack_select = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_97_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_branch_predict_pack_taken = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_97_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_phy_dst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_97_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_stale_dst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_97_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_arch_dst = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_97_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_98_inst_type = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_97_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_regWen = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_regWen :
    _io_o_issue_packs_1_T_97_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_src1_valid = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_97_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_phy_rs1 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_97_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_arch_rs1 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_97_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_98_src2_valid = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_97_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_phy_rs2 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_97_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_arch_rs2 = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_97_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_98_rob_idx = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_97_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_imm = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_imm :
    _io_o_issue_packs_1_T_97_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_src1_value = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_src1_value : _io_o_issue_packs_1_T_97_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_98_src2_value = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_src2_value : _io_o_issue_packs_1_T_97_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_98_op1_sel = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_97_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_98_op2_sel = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_97_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_98_alu_sel = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_97_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_98_branch_type = _io_o_issue_packs_1_T_29 ?
    reservation_station_29_io_o_uop_branch_type : _io_o_issue_packs_1_T_97_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_98_mem_type = _io_o_issue_packs_1_T_29 ? reservation_station_29_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_97_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_99_pc = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_pc :
    _io_o_issue_packs_1_T_98_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_99_inst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_inst :
    _io_o_issue_packs_1_T_98_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_func_code = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_func_code
     : _io_o_issue_packs_1_T_98_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_branch_predict_pack_valid = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_98_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_branch_predict_pack_target = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_98_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_99_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_98_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_branch_predict_pack_select = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_98_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_branch_predict_pack_taken = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_98_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_phy_dst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_98_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_stale_dst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_98_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_arch_dst = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_98_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_99_inst_type = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_98_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_regWen = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_regWen :
    _io_o_issue_packs_1_T_98_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_src1_valid = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_98_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_phy_rs1 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_98_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_arch_rs1 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_98_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_99_src2_valid = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_98_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_phy_rs2 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_98_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_arch_rs2 = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_98_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_99_rob_idx = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_98_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_imm = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_imm :
    _io_o_issue_packs_1_T_98_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_src1_value = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_src1_value : _io_o_issue_packs_1_T_98_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_99_src2_value = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_src2_value : _io_o_issue_packs_1_T_98_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_99_op1_sel = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_98_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_99_op2_sel = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_98_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_99_alu_sel = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_98_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_99_branch_type = _io_o_issue_packs_1_T_28 ?
    reservation_station_28_io_o_uop_branch_type : _io_o_issue_packs_1_T_98_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_99_mem_type = _io_o_issue_packs_1_T_28 ? reservation_station_28_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_98_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_100_pc = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_pc :
    _io_o_issue_packs_1_T_99_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_100_inst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_inst :
    _io_o_issue_packs_1_T_99_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_func_code = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_func_code
     : _io_o_issue_packs_1_T_99_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_branch_predict_pack_valid = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_99_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_branch_predict_pack_target = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_99_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_100_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_99_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_branch_predict_pack_select = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_99_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_branch_predict_pack_taken = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_99_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_phy_dst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_99_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_stale_dst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_99_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_arch_dst = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_99_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_100_inst_type = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_99_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_regWen = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_regWen :
    _io_o_issue_packs_1_T_99_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_src1_valid = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_99_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_phy_rs1 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_99_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_arch_rs1 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_99_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_100_src2_valid = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_99_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_phy_rs2 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_99_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_arch_rs2 = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_99_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_100_rob_idx = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_99_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_imm = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_imm :
    _io_o_issue_packs_1_T_99_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_src1_value = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_src1_value : _io_o_issue_packs_1_T_99_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_100_src2_value = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_src2_value : _io_o_issue_packs_1_T_99_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_100_op1_sel = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_99_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_100_op2_sel = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_99_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_100_alu_sel = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_99_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_100_branch_type = _io_o_issue_packs_1_T_27 ?
    reservation_station_27_io_o_uop_branch_type : _io_o_issue_packs_1_T_99_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_100_mem_type = _io_o_issue_packs_1_T_27 ? reservation_station_27_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_99_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_101_pc = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_pc :
    _io_o_issue_packs_1_T_100_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_101_inst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_inst :
    _io_o_issue_packs_1_T_100_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_func_code = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_func_code
     : _io_o_issue_packs_1_T_100_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_branch_predict_pack_valid = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_100_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_branch_predict_pack_target = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_100_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_101_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_100_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_branch_predict_pack_select = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_100_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_branch_predict_pack_taken = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_100_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_phy_dst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_100_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_stale_dst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_100_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_arch_dst = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_100_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_101_inst_type = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_100_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_regWen = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_regWen :
    _io_o_issue_packs_1_T_100_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_src1_valid = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_100_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_phy_rs1 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_100_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_arch_rs1 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_100_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_101_src2_valid = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_100_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_phy_rs2 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_100_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_arch_rs2 = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_100_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_101_rob_idx = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_100_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_imm = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_imm :
    _io_o_issue_packs_1_T_100_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_src1_value = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_src1_value : _io_o_issue_packs_1_T_100_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_101_src2_value = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_src2_value : _io_o_issue_packs_1_T_100_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_101_op1_sel = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_100_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_101_op2_sel = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_100_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_101_alu_sel = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_100_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_101_branch_type = _io_o_issue_packs_1_T_26 ?
    reservation_station_26_io_o_uop_branch_type : _io_o_issue_packs_1_T_100_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_101_mem_type = _io_o_issue_packs_1_T_26 ? reservation_station_26_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_100_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_102_pc = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_pc :
    _io_o_issue_packs_1_T_101_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_102_inst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_inst :
    _io_o_issue_packs_1_T_101_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_func_code = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_func_code
     : _io_o_issue_packs_1_T_101_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_branch_predict_pack_valid = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_101_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_branch_predict_pack_target = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_101_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_102_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_101_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_branch_predict_pack_select = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_101_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_branch_predict_pack_taken = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_101_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_phy_dst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_101_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_stale_dst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_101_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_arch_dst = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_101_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_102_inst_type = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_101_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_regWen = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_regWen :
    _io_o_issue_packs_1_T_101_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_src1_valid = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_101_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_phy_rs1 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_101_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_arch_rs1 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_101_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_102_src2_valid = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_101_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_phy_rs2 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_101_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_arch_rs2 = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_101_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_102_rob_idx = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_101_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_imm = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_imm :
    _io_o_issue_packs_1_T_101_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_src1_value = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_src1_value : _io_o_issue_packs_1_T_101_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_102_src2_value = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_src2_value : _io_o_issue_packs_1_T_101_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_102_op1_sel = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_101_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_102_op2_sel = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_101_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_102_alu_sel = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_101_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_102_branch_type = _io_o_issue_packs_1_T_25 ?
    reservation_station_25_io_o_uop_branch_type : _io_o_issue_packs_1_T_101_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_102_mem_type = _io_o_issue_packs_1_T_25 ? reservation_station_25_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_101_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_103_pc = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_pc :
    _io_o_issue_packs_1_T_102_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_103_inst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_inst :
    _io_o_issue_packs_1_T_102_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_func_code = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_func_code
     : _io_o_issue_packs_1_T_102_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_branch_predict_pack_valid = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_102_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_branch_predict_pack_target = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_102_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_103_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_102_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_branch_predict_pack_select = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_102_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_branch_predict_pack_taken = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_102_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_phy_dst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_102_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_stale_dst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_102_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_arch_dst = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_102_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_103_inst_type = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_102_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_regWen = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_regWen :
    _io_o_issue_packs_1_T_102_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_src1_valid = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_102_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_phy_rs1 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_102_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_arch_rs1 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_102_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_103_src2_valid = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_102_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_phy_rs2 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_102_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_arch_rs2 = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_102_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_103_rob_idx = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_102_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_imm = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_imm :
    _io_o_issue_packs_1_T_102_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_src1_value = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_src1_value : _io_o_issue_packs_1_T_102_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_103_src2_value = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_src2_value : _io_o_issue_packs_1_T_102_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_103_op1_sel = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_102_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_103_op2_sel = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_102_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_103_alu_sel = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_102_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_103_branch_type = _io_o_issue_packs_1_T_24 ?
    reservation_station_24_io_o_uop_branch_type : _io_o_issue_packs_1_T_102_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_103_mem_type = _io_o_issue_packs_1_T_24 ? reservation_station_24_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_102_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_104_pc = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_pc :
    _io_o_issue_packs_1_T_103_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_104_inst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_inst :
    _io_o_issue_packs_1_T_103_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_func_code = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_func_code
     : _io_o_issue_packs_1_T_103_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_branch_predict_pack_valid = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_103_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_branch_predict_pack_target = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_103_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_104_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_103_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_branch_predict_pack_select = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_103_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_branch_predict_pack_taken = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_103_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_phy_dst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_103_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_stale_dst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_103_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_arch_dst = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_103_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_104_inst_type = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_103_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_regWen = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_regWen :
    _io_o_issue_packs_1_T_103_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_src1_valid = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_103_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_phy_rs1 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_103_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_arch_rs1 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_103_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_104_src2_valid = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_103_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_phy_rs2 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_103_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_arch_rs2 = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_103_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_104_rob_idx = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_103_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_imm = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_imm :
    _io_o_issue_packs_1_T_103_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_src1_value = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_src1_value : _io_o_issue_packs_1_T_103_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_104_src2_value = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_src2_value : _io_o_issue_packs_1_T_103_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_104_op1_sel = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_103_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_104_op2_sel = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_103_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_104_alu_sel = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_103_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_104_branch_type = _io_o_issue_packs_1_T_23 ?
    reservation_station_23_io_o_uop_branch_type : _io_o_issue_packs_1_T_103_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_104_mem_type = _io_o_issue_packs_1_T_23 ? reservation_station_23_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_103_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_105_pc = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_pc :
    _io_o_issue_packs_1_T_104_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_105_inst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_inst :
    _io_o_issue_packs_1_T_104_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_func_code = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_func_code
     : _io_o_issue_packs_1_T_104_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_branch_predict_pack_valid = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_104_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_branch_predict_pack_target = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_104_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_105_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_104_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_branch_predict_pack_select = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_104_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_branch_predict_pack_taken = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_104_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_phy_dst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_104_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_stale_dst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_104_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_arch_dst = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_104_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_105_inst_type = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_104_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_regWen = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_regWen :
    _io_o_issue_packs_1_T_104_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_src1_valid = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_104_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_phy_rs1 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_104_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_arch_rs1 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_104_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_105_src2_valid = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_104_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_phy_rs2 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_104_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_arch_rs2 = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_104_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_105_rob_idx = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_104_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_imm = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_imm :
    _io_o_issue_packs_1_T_104_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_src1_value = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_src1_value : _io_o_issue_packs_1_T_104_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_105_src2_value = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_src2_value : _io_o_issue_packs_1_T_104_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_105_op1_sel = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_104_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_105_op2_sel = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_104_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_105_alu_sel = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_104_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_105_branch_type = _io_o_issue_packs_1_T_22 ?
    reservation_station_22_io_o_uop_branch_type : _io_o_issue_packs_1_T_104_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_105_mem_type = _io_o_issue_packs_1_T_22 ? reservation_station_22_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_104_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_106_pc = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_pc :
    _io_o_issue_packs_1_T_105_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_106_inst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_inst :
    _io_o_issue_packs_1_T_105_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_func_code = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_func_code
     : _io_o_issue_packs_1_T_105_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_branch_predict_pack_valid = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_105_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_branch_predict_pack_target = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_105_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_106_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_105_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_branch_predict_pack_select = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_105_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_branch_predict_pack_taken = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_105_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_phy_dst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_105_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_stale_dst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_105_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_arch_dst = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_105_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_106_inst_type = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_105_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_regWen = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_regWen :
    _io_o_issue_packs_1_T_105_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_src1_valid = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_105_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_phy_rs1 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_105_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_arch_rs1 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_105_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_106_src2_valid = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_105_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_phy_rs2 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_105_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_arch_rs2 = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_105_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_106_rob_idx = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_105_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_imm = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_imm :
    _io_o_issue_packs_1_T_105_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_src1_value = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_src1_value : _io_o_issue_packs_1_T_105_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_106_src2_value = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_src2_value : _io_o_issue_packs_1_T_105_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_106_op1_sel = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_105_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_106_op2_sel = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_105_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_106_alu_sel = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_105_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_106_branch_type = _io_o_issue_packs_1_T_21 ?
    reservation_station_21_io_o_uop_branch_type : _io_o_issue_packs_1_T_105_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_106_mem_type = _io_o_issue_packs_1_T_21 ? reservation_station_21_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_105_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_107_pc = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_pc :
    _io_o_issue_packs_1_T_106_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_107_inst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_inst :
    _io_o_issue_packs_1_T_106_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_func_code = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_func_code
     : _io_o_issue_packs_1_T_106_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_branch_predict_pack_valid = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_106_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_branch_predict_pack_target = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_106_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_107_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_106_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_branch_predict_pack_select = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_106_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_branch_predict_pack_taken = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_106_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_phy_dst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_106_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_stale_dst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_106_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_arch_dst = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_106_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_107_inst_type = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_106_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_regWen = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_regWen :
    _io_o_issue_packs_1_T_106_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_src1_valid = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_106_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_phy_rs1 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_106_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_arch_rs1 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_106_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_107_src2_valid = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_106_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_phy_rs2 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_106_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_arch_rs2 = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_106_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_107_rob_idx = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_106_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_imm = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_imm :
    _io_o_issue_packs_1_T_106_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_src1_value = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_src1_value : _io_o_issue_packs_1_T_106_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_107_src2_value = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_src2_value : _io_o_issue_packs_1_T_106_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_107_op1_sel = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_106_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_107_op2_sel = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_106_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_107_alu_sel = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_106_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_107_branch_type = _io_o_issue_packs_1_T_20 ?
    reservation_station_20_io_o_uop_branch_type : _io_o_issue_packs_1_T_106_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_107_mem_type = _io_o_issue_packs_1_T_20 ? reservation_station_20_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_106_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_108_pc = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_pc :
    _io_o_issue_packs_1_T_107_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_108_inst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_inst :
    _io_o_issue_packs_1_T_107_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_func_code = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_func_code
     : _io_o_issue_packs_1_T_107_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_branch_predict_pack_valid = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_107_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_branch_predict_pack_target = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_107_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_108_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_107_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_branch_predict_pack_select = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_107_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_branch_predict_pack_taken = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_107_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_phy_dst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_107_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_stale_dst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_107_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_arch_dst = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_107_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_108_inst_type = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_107_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_regWen = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_regWen :
    _io_o_issue_packs_1_T_107_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_src1_valid = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_107_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_phy_rs1 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_107_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_arch_rs1 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_107_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_108_src2_valid = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_107_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_phy_rs2 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_107_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_arch_rs2 = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_107_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_108_rob_idx = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_107_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_imm = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_imm :
    _io_o_issue_packs_1_T_107_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_src1_value = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_src1_value : _io_o_issue_packs_1_T_107_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_108_src2_value = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_src2_value : _io_o_issue_packs_1_T_107_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_108_op1_sel = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_107_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_108_op2_sel = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_107_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_108_alu_sel = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_107_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_108_branch_type = _io_o_issue_packs_1_T_19 ?
    reservation_station_19_io_o_uop_branch_type : _io_o_issue_packs_1_T_107_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_108_mem_type = _io_o_issue_packs_1_T_19 ? reservation_station_19_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_107_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_109_pc = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_pc :
    _io_o_issue_packs_1_T_108_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_109_inst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_inst :
    _io_o_issue_packs_1_T_108_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_func_code = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_func_code
     : _io_o_issue_packs_1_T_108_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_branch_predict_pack_valid = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_108_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_branch_predict_pack_target = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_108_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_109_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_108_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_branch_predict_pack_select = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_108_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_branch_predict_pack_taken = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_108_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_phy_dst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_108_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_stale_dst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_108_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_arch_dst = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_108_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_109_inst_type = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_108_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_regWen = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_regWen :
    _io_o_issue_packs_1_T_108_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_src1_valid = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_108_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_phy_rs1 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_108_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_arch_rs1 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_108_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_109_src2_valid = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_108_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_phy_rs2 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_108_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_arch_rs2 = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_108_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_109_rob_idx = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_108_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_imm = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_imm :
    _io_o_issue_packs_1_T_108_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_src1_value = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_src1_value : _io_o_issue_packs_1_T_108_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_109_src2_value = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_src2_value : _io_o_issue_packs_1_T_108_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_109_op1_sel = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_108_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_109_op2_sel = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_108_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_109_alu_sel = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_108_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_109_branch_type = _io_o_issue_packs_1_T_18 ?
    reservation_station_18_io_o_uop_branch_type : _io_o_issue_packs_1_T_108_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_109_mem_type = _io_o_issue_packs_1_T_18 ? reservation_station_18_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_108_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_110_pc = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_pc :
    _io_o_issue_packs_1_T_109_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_110_inst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_inst :
    _io_o_issue_packs_1_T_109_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_func_code = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_func_code
     : _io_o_issue_packs_1_T_109_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_branch_predict_pack_valid = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_109_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_branch_predict_pack_target = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_109_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_110_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_109_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_branch_predict_pack_select = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_109_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_branch_predict_pack_taken = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_109_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_phy_dst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_109_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_stale_dst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_109_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_arch_dst = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_109_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_110_inst_type = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_109_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_regWen = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_regWen :
    _io_o_issue_packs_1_T_109_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_src1_valid = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_109_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_phy_rs1 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_109_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_arch_rs1 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_109_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_110_src2_valid = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_109_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_phy_rs2 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_109_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_arch_rs2 = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_109_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_110_rob_idx = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_109_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_imm = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_imm :
    _io_o_issue_packs_1_T_109_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_src1_value = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_src1_value : _io_o_issue_packs_1_T_109_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_110_src2_value = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_src2_value : _io_o_issue_packs_1_T_109_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_110_op1_sel = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_109_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_110_op2_sel = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_109_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_110_alu_sel = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_109_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_110_branch_type = _io_o_issue_packs_1_T_17 ?
    reservation_station_17_io_o_uop_branch_type : _io_o_issue_packs_1_T_109_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_110_mem_type = _io_o_issue_packs_1_T_17 ? reservation_station_17_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_109_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_111_pc = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_pc :
    _io_o_issue_packs_1_T_110_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_111_inst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_inst :
    _io_o_issue_packs_1_T_110_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_func_code = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_func_code
     : _io_o_issue_packs_1_T_110_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_branch_predict_pack_valid = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_110_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_branch_predict_pack_target = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_110_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_111_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_110_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_branch_predict_pack_select = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_110_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_branch_predict_pack_taken = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_110_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_phy_dst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_110_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_stale_dst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_110_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_arch_dst = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_110_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_111_inst_type = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_110_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_regWen = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_regWen :
    _io_o_issue_packs_1_T_110_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_src1_valid = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_110_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_phy_rs1 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_110_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_arch_rs1 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_110_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_111_src2_valid = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_110_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_phy_rs2 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_110_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_arch_rs2 = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_110_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_111_rob_idx = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_110_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_imm = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_imm :
    _io_o_issue_packs_1_T_110_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_src1_value = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_src1_value : _io_o_issue_packs_1_T_110_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_111_src2_value = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_src2_value : _io_o_issue_packs_1_T_110_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_111_op1_sel = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_110_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_111_op2_sel = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_110_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_111_alu_sel = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_110_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_111_branch_type = _io_o_issue_packs_1_T_16 ?
    reservation_station_16_io_o_uop_branch_type : _io_o_issue_packs_1_T_110_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_111_mem_type = _io_o_issue_packs_1_T_16 ? reservation_station_16_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_110_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_112_pc = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_pc :
    _io_o_issue_packs_1_T_111_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_112_inst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_inst :
    _io_o_issue_packs_1_T_111_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_func_code = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_func_code
     : _io_o_issue_packs_1_T_111_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_branch_predict_pack_valid = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_111_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_branch_predict_pack_target = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_111_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_112_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_111_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_branch_predict_pack_select = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_111_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_branch_predict_pack_taken = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_111_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_phy_dst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_111_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_stale_dst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_111_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_arch_dst = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_111_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_112_inst_type = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_111_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_regWen = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_regWen :
    _io_o_issue_packs_1_T_111_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_src1_valid = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_111_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_phy_rs1 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_111_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_arch_rs1 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_111_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_112_src2_valid = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_111_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_phy_rs2 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_111_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_arch_rs2 = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_111_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_112_rob_idx = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_111_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_imm = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_imm :
    _io_o_issue_packs_1_T_111_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_src1_value = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_src1_value : _io_o_issue_packs_1_T_111_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_112_src2_value = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_src2_value : _io_o_issue_packs_1_T_111_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_112_op1_sel = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_111_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_112_op2_sel = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_111_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_112_alu_sel = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_111_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_112_branch_type = _io_o_issue_packs_1_T_15 ?
    reservation_station_15_io_o_uop_branch_type : _io_o_issue_packs_1_T_111_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_112_mem_type = _io_o_issue_packs_1_T_15 ? reservation_station_15_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_111_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_113_pc = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_pc :
    _io_o_issue_packs_1_T_112_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_113_inst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_inst :
    _io_o_issue_packs_1_T_112_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_func_code = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_func_code
     : _io_o_issue_packs_1_T_112_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_branch_predict_pack_valid = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_112_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_branch_predict_pack_target = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_112_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_113_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_112_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_branch_predict_pack_select = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_112_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_branch_predict_pack_taken = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_112_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_phy_dst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_112_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_stale_dst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_112_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_arch_dst = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_112_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_113_inst_type = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_112_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_regWen = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_regWen :
    _io_o_issue_packs_1_T_112_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_src1_valid = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_112_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_phy_rs1 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_112_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_arch_rs1 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_112_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_113_src2_valid = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_112_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_phy_rs2 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_112_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_arch_rs2 = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_112_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_113_rob_idx = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_112_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_imm = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_imm :
    _io_o_issue_packs_1_T_112_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_src1_value = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_src1_value : _io_o_issue_packs_1_T_112_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_113_src2_value = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_src2_value : _io_o_issue_packs_1_T_112_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_113_op1_sel = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_112_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_113_op2_sel = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_112_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_113_alu_sel = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_112_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_113_branch_type = _io_o_issue_packs_1_T_14 ?
    reservation_station_14_io_o_uop_branch_type : _io_o_issue_packs_1_T_112_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_113_mem_type = _io_o_issue_packs_1_T_14 ? reservation_station_14_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_112_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_114_pc = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_pc :
    _io_o_issue_packs_1_T_113_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_114_inst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_inst :
    _io_o_issue_packs_1_T_113_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_func_code = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_func_code
     : _io_o_issue_packs_1_T_113_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_branch_predict_pack_valid = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_113_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_branch_predict_pack_target = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_113_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_114_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_113_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_branch_predict_pack_select = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_113_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_branch_predict_pack_taken = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_113_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_phy_dst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_113_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_stale_dst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_113_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_arch_dst = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_113_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_114_inst_type = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_113_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_regWen = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_regWen :
    _io_o_issue_packs_1_T_113_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_src1_valid = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_113_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_phy_rs1 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_113_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_arch_rs1 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_113_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_114_src2_valid = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_113_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_phy_rs2 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_113_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_arch_rs2 = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_113_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_114_rob_idx = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_113_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_imm = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_imm :
    _io_o_issue_packs_1_T_113_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_src1_value = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_src1_value : _io_o_issue_packs_1_T_113_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_114_src2_value = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_src2_value : _io_o_issue_packs_1_T_113_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_114_op1_sel = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_113_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_114_op2_sel = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_113_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_114_alu_sel = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_113_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_114_branch_type = _io_o_issue_packs_1_T_13 ?
    reservation_station_13_io_o_uop_branch_type : _io_o_issue_packs_1_T_113_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_114_mem_type = _io_o_issue_packs_1_T_13 ? reservation_station_13_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_113_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_115_pc = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_pc :
    _io_o_issue_packs_1_T_114_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_115_inst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_inst :
    _io_o_issue_packs_1_T_114_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_func_code = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_func_code
     : _io_o_issue_packs_1_T_114_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_branch_predict_pack_valid = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_114_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_branch_predict_pack_target = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_114_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_115_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_114_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_branch_predict_pack_select = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_114_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_branch_predict_pack_taken = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_114_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_phy_dst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_114_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_stale_dst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_114_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_arch_dst = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_114_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_115_inst_type = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_114_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_regWen = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_regWen :
    _io_o_issue_packs_1_T_114_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_src1_valid = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_114_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_phy_rs1 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_114_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_arch_rs1 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_114_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_115_src2_valid = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_114_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_phy_rs2 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_114_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_arch_rs2 = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_114_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_115_rob_idx = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_114_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_imm = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_imm :
    _io_o_issue_packs_1_T_114_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_src1_value = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_src1_value : _io_o_issue_packs_1_T_114_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_115_src2_value = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_src2_value : _io_o_issue_packs_1_T_114_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_115_op1_sel = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_114_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_115_op2_sel = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_114_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_115_alu_sel = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_114_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_115_branch_type = _io_o_issue_packs_1_T_12 ?
    reservation_station_12_io_o_uop_branch_type : _io_o_issue_packs_1_T_114_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_115_mem_type = _io_o_issue_packs_1_T_12 ? reservation_station_12_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_114_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_116_pc = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_pc :
    _io_o_issue_packs_1_T_115_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_116_inst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_inst :
    _io_o_issue_packs_1_T_115_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_func_code = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_func_code
     : _io_o_issue_packs_1_T_115_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_branch_predict_pack_valid = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_115_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_branch_predict_pack_target = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_115_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_116_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_115_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_branch_predict_pack_select = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_115_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_branch_predict_pack_taken = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_115_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_phy_dst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_115_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_stale_dst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_115_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_arch_dst = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_115_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_116_inst_type = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_115_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_regWen = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_regWen :
    _io_o_issue_packs_1_T_115_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_src1_valid = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_115_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_phy_rs1 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_115_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_arch_rs1 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_115_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_116_src2_valid = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_115_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_phy_rs2 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_115_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_arch_rs2 = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_115_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_116_rob_idx = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_115_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_imm = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_imm :
    _io_o_issue_packs_1_T_115_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_src1_value = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_src1_value : _io_o_issue_packs_1_T_115_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_116_src2_value = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_src2_value : _io_o_issue_packs_1_T_115_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_116_op1_sel = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_115_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_116_op2_sel = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_115_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_116_alu_sel = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_115_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_116_branch_type = _io_o_issue_packs_1_T_11 ?
    reservation_station_11_io_o_uop_branch_type : _io_o_issue_packs_1_T_115_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_116_mem_type = _io_o_issue_packs_1_T_11 ? reservation_station_11_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_115_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_117_pc = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_pc :
    _io_o_issue_packs_1_T_116_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_117_inst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_inst :
    _io_o_issue_packs_1_T_116_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_func_code = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_func_code
     : _io_o_issue_packs_1_T_116_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_branch_predict_pack_valid = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_116_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_branch_predict_pack_target = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_116_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_117_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_116_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_branch_predict_pack_select = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_116_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_branch_predict_pack_taken = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_116_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_phy_dst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_116_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_stale_dst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_stale_dst
     : _io_o_issue_packs_1_T_116_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_arch_dst = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_116_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_117_inst_type = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_inst_type
     : _io_o_issue_packs_1_T_116_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_regWen = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_regWen :
    _io_o_issue_packs_1_T_116_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_src1_valid = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_116_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_phy_rs1 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_116_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_arch_rs1 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_116_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_117_src2_valid = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_116_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_phy_rs2 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_116_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_arch_rs2 = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_116_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_117_rob_idx = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_116_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_imm = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_imm :
    _io_o_issue_packs_1_T_116_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_src1_value = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_src1_value : _io_o_issue_packs_1_T_116_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_117_src2_value = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_src2_value : _io_o_issue_packs_1_T_116_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_117_op1_sel = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_116_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_117_op2_sel = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_116_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_117_alu_sel = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_116_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_117_branch_type = _io_o_issue_packs_1_T_10 ?
    reservation_station_10_io_o_uop_branch_type : _io_o_issue_packs_1_T_116_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_117_mem_type = _io_o_issue_packs_1_T_10 ? reservation_station_10_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_116_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_118_pc = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_pc :
    _io_o_issue_packs_1_T_117_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_118_inst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_inst :
    _io_o_issue_packs_1_T_117_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_func_code = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_func_code :
    _io_o_issue_packs_1_T_117_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_branch_predict_pack_valid = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_117_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_branch_predict_pack_target = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_117_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_118_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_117_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_branch_predict_pack_select = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_117_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_branch_predict_pack_taken = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_117_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_phy_dst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_117_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_stale_dst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_117_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_arch_dst = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_117_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_118_inst_type = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_117_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_regWen = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_regWen :
    _io_o_issue_packs_1_T_117_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_src1_valid = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_117_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_phy_rs1 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_117_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_arch_rs1 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_117_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_118_src2_valid = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_117_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_phy_rs2 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_117_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_arch_rs2 = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_117_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_118_rob_idx = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_117_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_imm = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_imm :
    _io_o_issue_packs_1_T_117_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_src1_value = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_117_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_118_src2_value = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_117_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_118_op1_sel = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_117_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_118_op2_sel = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_117_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_118_alu_sel = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_117_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_118_branch_type = _io_o_issue_packs_1_T_9 ?
    reservation_station_9_io_o_uop_branch_type : _io_o_issue_packs_1_T_117_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_118_mem_type = _io_o_issue_packs_1_T_9 ? reservation_station_9_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_117_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_119_pc = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_pc :
    _io_o_issue_packs_1_T_118_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_119_inst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_inst :
    _io_o_issue_packs_1_T_118_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_func_code = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_func_code :
    _io_o_issue_packs_1_T_118_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_branch_predict_pack_valid = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_118_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_branch_predict_pack_target = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_118_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_119_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_118_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_branch_predict_pack_select = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_118_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_branch_predict_pack_taken = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_118_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_phy_dst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_118_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_stale_dst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_118_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_arch_dst = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_118_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_119_inst_type = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_118_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_regWen = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_regWen :
    _io_o_issue_packs_1_T_118_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_src1_valid = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_118_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_phy_rs1 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_118_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_arch_rs1 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_118_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_119_src2_valid = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_118_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_phy_rs2 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_118_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_arch_rs2 = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_118_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_119_rob_idx = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_118_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_imm = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_imm :
    _io_o_issue_packs_1_T_118_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_src1_value = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_118_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_119_src2_value = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_118_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_119_op1_sel = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_118_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_119_op2_sel = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_118_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_119_alu_sel = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_118_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_119_branch_type = _io_o_issue_packs_1_T_8 ?
    reservation_station_8_io_o_uop_branch_type : _io_o_issue_packs_1_T_118_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_119_mem_type = _io_o_issue_packs_1_T_8 ? reservation_station_8_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_118_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_120_pc = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_pc :
    _io_o_issue_packs_1_T_119_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_120_inst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_inst :
    _io_o_issue_packs_1_T_119_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_func_code = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_func_code :
    _io_o_issue_packs_1_T_119_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_branch_predict_pack_valid = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_119_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_branch_predict_pack_target = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_119_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_120_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_119_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_branch_predict_pack_select = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_119_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_branch_predict_pack_taken = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_119_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_phy_dst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_119_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_stale_dst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_119_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_arch_dst = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_119_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_120_inst_type = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_119_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_regWen = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_regWen :
    _io_o_issue_packs_1_T_119_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_src1_valid = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_119_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_phy_rs1 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_119_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_arch_rs1 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_119_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_120_src2_valid = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_119_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_phy_rs2 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_119_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_arch_rs2 = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_119_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_120_rob_idx = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_119_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_imm = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_imm :
    _io_o_issue_packs_1_T_119_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_src1_value = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_119_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_120_src2_value = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_119_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_120_op1_sel = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_119_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_120_op2_sel = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_119_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_120_alu_sel = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_119_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_120_branch_type = _io_o_issue_packs_1_T_7 ?
    reservation_station_7_io_o_uop_branch_type : _io_o_issue_packs_1_T_119_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_120_mem_type = _io_o_issue_packs_1_T_7 ? reservation_station_7_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_119_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_121_pc = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_pc :
    _io_o_issue_packs_1_T_120_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_121_inst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_inst :
    _io_o_issue_packs_1_T_120_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_func_code = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_func_code :
    _io_o_issue_packs_1_T_120_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_branch_predict_pack_valid = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_120_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_branch_predict_pack_target = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_120_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_121_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_120_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_branch_predict_pack_select = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_120_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_branch_predict_pack_taken = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_120_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_phy_dst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_120_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_stale_dst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_120_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_arch_dst = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_120_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_121_inst_type = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_120_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_regWen = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_regWen :
    _io_o_issue_packs_1_T_120_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_src1_valid = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_120_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_phy_rs1 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_120_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_arch_rs1 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_120_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_121_src2_valid = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_120_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_phy_rs2 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_120_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_arch_rs2 = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_120_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_121_rob_idx = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_120_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_imm = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_imm :
    _io_o_issue_packs_1_T_120_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_src1_value = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_120_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_121_src2_value = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_120_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_121_op1_sel = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_120_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_121_op2_sel = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_120_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_121_alu_sel = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_120_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_121_branch_type = _io_o_issue_packs_1_T_6 ?
    reservation_station_6_io_o_uop_branch_type : _io_o_issue_packs_1_T_120_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_121_mem_type = _io_o_issue_packs_1_T_6 ? reservation_station_6_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_120_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_122_pc = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_pc :
    _io_o_issue_packs_1_T_121_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_122_inst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_inst :
    _io_o_issue_packs_1_T_121_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_func_code = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_func_code :
    _io_o_issue_packs_1_T_121_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_branch_predict_pack_valid = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_121_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_branch_predict_pack_target = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_121_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_122_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_121_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_branch_predict_pack_select = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_121_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_branch_predict_pack_taken = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_121_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_phy_dst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_121_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_stale_dst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_121_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_arch_dst = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_121_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_122_inst_type = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_121_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_regWen = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_regWen :
    _io_o_issue_packs_1_T_121_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_src1_valid = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_121_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_phy_rs1 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_121_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_arch_rs1 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_121_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_122_src2_valid = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_121_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_phy_rs2 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_121_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_arch_rs2 = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_121_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_122_rob_idx = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_121_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_imm = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_imm :
    _io_o_issue_packs_1_T_121_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_src1_value = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_121_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_122_src2_value = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_121_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_122_op1_sel = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_121_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_122_op2_sel = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_121_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_122_alu_sel = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_121_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_122_branch_type = _io_o_issue_packs_1_T_5 ?
    reservation_station_5_io_o_uop_branch_type : _io_o_issue_packs_1_T_121_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_122_mem_type = _io_o_issue_packs_1_T_5 ? reservation_station_5_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_121_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_123_pc = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_pc :
    _io_o_issue_packs_1_T_122_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_123_inst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_inst :
    _io_o_issue_packs_1_T_122_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_func_code = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_func_code :
    _io_o_issue_packs_1_T_122_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_branch_predict_pack_valid = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_122_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_branch_predict_pack_target = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_122_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_123_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_122_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_branch_predict_pack_select = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_122_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_branch_predict_pack_taken = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_122_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_phy_dst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_122_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_stale_dst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_122_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_arch_dst = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_122_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_123_inst_type = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_122_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_regWen = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_regWen :
    _io_o_issue_packs_1_T_122_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_src1_valid = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_122_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_phy_rs1 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_122_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_arch_rs1 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_122_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_123_src2_valid = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_122_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_phy_rs2 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_122_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_arch_rs2 = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_122_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_123_rob_idx = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_122_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_imm = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_imm :
    _io_o_issue_packs_1_T_122_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_src1_value = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_122_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_123_src2_value = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_122_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_123_op1_sel = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_122_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_123_op2_sel = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_122_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_123_alu_sel = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_122_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_123_branch_type = _io_o_issue_packs_1_T_4 ?
    reservation_station_4_io_o_uop_branch_type : _io_o_issue_packs_1_T_122_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_123_mem_type = _io_o_issue_packs_1_T_4 ? reservation_station_4_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_122_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_124_pc = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_pc :
    _io_o_issue_packs_1_T_123_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_124_inst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_inst :
    _io_o_issue_packs_1_T_123_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_func_code = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_func_code :
    _io_o_issue_packs_1_T_123_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_branch_predict_pack_valid = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_123_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_branch_predict_pack_target = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_123_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_124_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_123_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_branch_predict_pack_select = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_123_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_branch_predict_pack_taken = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_123_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_phy_dst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_123_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_stale_dst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_123_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_arch_dst = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_123_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_124_inst_type = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_123_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_regWen = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_regWen :
    _io_o_issue_packs_1_T_123_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_src1_valid = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_123_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_phy_rs1 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_123_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_arch_rs1 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_123_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_124_src2_valid = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_123_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_phy_rs2 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_123_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_arch_rs2 = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_123_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_124_rob_idx = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_123_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_imm = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_imm :
    _io_o_issue_packs_1_T_123_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_src1_value = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_123_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_124_src2_value = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_123_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_124_op1_sel = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_123_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_124_op2_sel = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_123_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_124_alu_sel = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_123_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_124_branch_type = _io_o_issue_packs_1_T_3 ?
    reservation_station_3_io_o_uop_branch_type : _io_o_issue_packs_1_T_123_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_124_mem_type = _io_o_issue_packs_1_T_3 ? reservation_station_3_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_123_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_125_pc = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_pc :
    _io_o_issue_packs_1_T_124_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_125_inst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_inst :
    _io_o_issue_packs_1_T_124_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_func_code = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_func_code :
    _io_o_issue_packs_1_T_124_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_branch_predict_pack_valid = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_124_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_branch_predict_pack_target = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_124_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_125_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_124_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_branch_predict_pack_select = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_124_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_branch_predict_pack_taken = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_124_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_phy_dst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_124_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_stale_dst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_124_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_arch_dst = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_124_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_125_inst_type = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_124_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_regWen = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_regWen :
    _io_o_issue_packs_1_T_124_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_src1_valid = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_124_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_phy_rs1 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_124_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_arch_rs1 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_124_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_125_src2_valid = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_124_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_phy_rs2 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_124_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_arch_rs2 = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_124_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_125_rob_idx = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_124_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_imm = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_imm :
    _io_o_issue_packs_1_T_124_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_src1_value = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_124_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_125_src2_value = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_124_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_125_op1_sel = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_124_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_125_op2_sel = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_124_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_125_alu_sel = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_124_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_125_branch_type = _io_o_issue_packs_1_T_2 ?
    reservation_station_2_io_o_uop_branch_type : _io_o_issue_packs_1_T_124_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_125_mem_type = _io_o_issue_packs_1_T_2 ? reservation_station_2_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_124_mem_type; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_126_pc = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_pc :
    _io_o_issue_packs_1_T_125_pc; // @[Mux.scala 101:16]
  wire [31:0] _io_o_issue_packs_1_T_126_inst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_inst :
    _io_o_issue_packs_1_T_125_inst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_func_code = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_func_code :
    _io_o_issue_packs_1_T_125_func_code; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_branch_predict_pack_valid = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_125_branch_predict_pack_valid; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_branch_predict_pack_target = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_125_branch_predict_pack_target; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_126_branch_predict_pack_branch_type = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_125_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_branch_predict_pack_select = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_125_branch_predict_pack_select; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_branch_predict_pack_taken = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_125_branch_predict_pack_taken; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_phy_dst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_125_phy_dst; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_stale_dst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_125_stale_dst; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_arch_dst = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_125_arch_dst; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_126_inst_type = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_125_inst_type; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_regWen = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_regWen :
    _io_o_issue_packs_1_T_125_regWen; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_src1_valid = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_125_src1_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_phy_rs1 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_125_phy_rs1; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_arch_rs1 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_125_arch_rs1; // @[Mux.scala 101:16]
  wire  _io_o_issue_packs_1_T_126_src2_valid = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_125_src2_valid; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_phy_rs2 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_125_phy_rs2; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_arch_rs2 = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_125_arch_rs2; // @[Mux.scala 101:16]
  wire [6:0] _io_o_issue_packs_1_T_126_rob_idx = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_125_rob_idx; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_imm = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_imm :
    _io_o_issue_packs_1_T_125_imm; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_src1_value = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src1_value
     : _io_o_issue_packs_1_T_125_src1_value; // @[Mux.scala 101:16]
  wire [63:0] _io_o_issue_packs_1_T_126_src2_value = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_src2_value
     : _io_o_issue_packs_1_T_125_src2_value; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_126_op1_sel = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_125_op1_sel; // @[Mux.scala 101:16]
  wire [2:0] _io_o_issue_packs_1_T_126_op2_sel = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_125_op2_sel; // @[Mux.scala 101:16]
  wire [4:0] _io_o_issue_packs_1_T_126_alu_sel = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_125_alu_sel; // @[Mux.scala 101:16]
  wire [3:0] _io_o_issue_packs_1_T_126_branch_type = _io_o_issue_packs_1_T_1 ?
    reservation_station_1_io_o_uop_branch_type : _io_o_issue_packs_1_T_125_branch_type; // @[Mux.scala 101:16]
  wire [1:0] _io_o_issue_packs_1_T_126_mem_type = _io_o_issue_packs_1_T_1 ? reservation_station_1_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_125_mem_type; // @[Mux.scala 101:16]
  wire  _reservation_station_0_io_i_write_slot_T = 6'h0 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_0_io_i_write_slot_T_2 = 6'h0 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_0_io_i_write_slot_T_5 = 6'h0 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_1_io_i_write_slot_T = 6'h1 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_1_io_i_write_slot_T_2 = 6'h1 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_1_io_i_write_slot_T_5 = 6'h1 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_2_io_i_write_slot_T = 6'h2 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_2_io_i_write_slot_T_2 = 6'h2 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_2_io_i_write_slot_T_5 = 6'h2 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_3_io_i_write_slot_T = 6'h3 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_3_io_i_write_slot_T_2 = 6'h3 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_3_io_i_write_slot_T_5 = 6'h3 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_4_io_i_write_slot_T = 6'h4 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_4_io_i_write_slot_T_2 = 6'h4 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_4_io_i_write_slot_T_5 = 6'h4 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_5_io_i_write_slot_T = 6'h5 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_5_io_i_write_slot_T_2 = 6'h5 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_5_io_i_write_slot_T_5 = 6'h5 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_6_io_i_write_slot_T = 6'h6 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_6_io_i_write_slot_T_2 = 6'h6 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_6_io_i_write_slot_T_5 = 6'h6 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_7_io_i_write_slot_T = 6'h7 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_7_io_i_write_slot_T_2 = 6'h7 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_7_io_i_write_slot_T_5 = 6'h7 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_8_io_i_write_slot_T = 6'h8 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_8_io_i_write_slot_T_2 = 6'h8 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_8_io_i_write_slot_T_5 = 6'h8 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_9_io_i_write_slot_T = 6'h9 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_9_io_i_write_slot_T_2 = 6'h9 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_9_io_i_write_slot_T_5 = 6'h9 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_10_io_i_write_slot_T = 6'ha == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_10_io_i_write_slot_T_2 = 6'ha == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_10_io_i_write_slot_T_5 = 6'ha == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_11_io_i_write_slot_T = 6'hb == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_11_io_i_write_slot_T_2 = 6'hb == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_11_io_i_write_slot_T_5 = 6'hb == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_12_io_i_write_slot_T = 6'hc == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_12_io_i_write_slot_T_2 = 6'hc == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_12_io_i_write_slot_T_5 = 6'hc == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_13_io_i_write_slot_T = 6'hd == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_13_io_i_write_slot_T_2 = 6'hd == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_13_io_i_write_slot_T_5 = 6'hd == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_14_io_i_write_slot_T = 6'he == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_14_io_i_write_slot_T_2 = 6'he == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_14_io_i_write_slot_T_5 = 6'he == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_15_io_i_write_slot_T = 6'hf == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_15_io_i_write_slot_T_2 = 6'hf == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_15_io_i_write_slot_T_5 = 6'hf == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_16_io_i_write_slot_T = 6'h10 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_16_io_i_write_slot_T_2 = 6'h10 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_16_io_i_write_slot_T_5 = 6'h10 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_17_io_i_write_slot_T = 6'h11 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_17_io_i_write_slot_T_2 = 6'h11 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_17_io_i_write_slot_T_5 = 6'h11 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_18_io_i_write_slot_T = 6'h12 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_18_io_i_write_slot_T_2 = 6'h12 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_18_io_i_write_slot_T_5 = 6'h12 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_19_io_i_write_slot_T = 6'h13 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_19_io_i_write_slot_T_2 = 6'h13 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_19_io_i_write_slot_T_5 = 6'h13 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_20_io_i_write_slot_T = 6'h14 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_20_io_i_write_slot_T_2 = 6'h14 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_20_io_i_write_slot_T_5 = 6'h14 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_21_io_i_write_slot_T = 6'h15 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_21_io_i_write_slot_T_2 = 6'h15 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_21_io_i_write_slot_T_5 = 6'h15 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_22_io_i_write_slot_T = 6'h16 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_22_io_i_write_slot_T_2 = 6'h16 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_22_io_i_write_slot_T_5 = 6'h16 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_23_io_i_write_slot_T = 6'h17 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_23_io_i_write_slot_T_2 = 6'h17 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_23_io_i_write_slot_T_5 = 6'h17 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_24_io_i_write_slot_T = 6'h18 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_24_io_i_write_slot_T_2 = 6'h18 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_24_io_i_write_slot_T_5 = 6'h18 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_25_io_i_write_slot_T = 6'h19 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_25_io_i_write_slot_T_2 = 6'h19 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_25_io_i_write_slot_T_5 = 6'h19 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_26_io_i_write_slot_T = 6'h1a == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_26_io_i_write_slot_T_2 = 6'h1a == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_26_io_i_write_slot_T_5 = 6'h1a == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_27_io_i_write_slot_T = 6'h1b == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_27_io_i_write_slot_T_2 = 6'h1b == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_27_io_i_write_slot_T_5 = 6'h1b == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_28_io_i_write_slot_T = 6'h1c == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_28_io_i_write_slot_T_2 = 6'h1c == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_28_io_i_write_slot_T_5 = 6'h1c == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_29_io_i_write_slot_T = 6'h1d == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_29_io_i_write_slot_T_2 = 6'h1d == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_29_io_i_write_slot_T_5 = 6'h1d == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_30_io_i_write_slot_T = 6'h1e == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_30_io_i_write_slot_T_2 = 6'h1e == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_30_io_i_write_slot_T_5 = 6'h1e == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_31_io_i_write_slot_T = 6'h1f == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_31_io_i_write_slot_T_2 = 6'h1f == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_31_io_i_write_slot_T_5 = 6'h1f == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_32_io_i_write_slot_T = 6'h20 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_32_io_i_write_slot_T_2 = 6'h20 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_32_io_i_write_slot_T_5 = 6'h20 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_33_io_i_write_slot_T = 6'h21 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_33_io_i_write_slot_T_2 = 6'h21 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_33_io_i_write_slot_T_5 = 6'h21 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_34_io_i_write_slot_T = 6'h22 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_34_io_i_write_slot_T_2 = 6'h22 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_34_io_i_write_slot_T_5 = 6'h22 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_35_io_i_write_slot_T = 6'h23 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_35_io_i_write_slot_T_2 = 6'h23 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_35_io_i_write_slot_T_5 = 6'h23 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_36_io_i_write_slot_T = 6'h24 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_36_io_i_write_slot_T_2 = 6'h24 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_36_io_i_write_slot_T_5 = 6'h24 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_37_io_i_write_slot_T = 6'h25 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_37_io_i_write_slot_T_2 = 6'h25 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_37_io_i_write_slot_T_5 = 6'h25 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_38_io_i_write_slot_T = 6'h26 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_38_io_i_write_slot_T_2 = 6'h26 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_38_io_i_write_slot_T_5 = 6'h26 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_39_io_i_write_slot_T = 6'h27 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_39_io_i_write_slot_T_2 = 6'h27 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_39_io_i_write_slot_T_5 = 6'h27 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_40_io_i_write_slot_T = 6'h28 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_40_io_i_write_slot_T_2 = 6'h28 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_40_io_i_write_slot_T_5 = 6'h28 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_41_io_i_write_slot_T = 6'h29 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_41_io_i_write_slot_T_2 = 6'h29 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_41_io_i_write_slot_T_5 = 6'h29 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_42_io_i_write_slot_T = 6'h2a == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_42_io_i_write_slot_T_2 = 6'h2a == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_42_io_i_write_slot_T_5 = 6'h2a == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_43_io_i_write_slot_T = 6'h2b == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_43_io_i_write_slot_T_2 = 6'h2b == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_43_io_i_write_slot_T_5 = 6'h2b == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_44_io_i_write_slot_T = 6'h2c == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_44_io_i_write_slot_T_2 = 6'h2c == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_44_io_i_write_slot_T_5 = 6'h2c == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_45_io_i_write_slot_T = 6'h2d == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_45_io_i_write_slot_T_2 = 6'h2d == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_45_io_i_write_slot_T_5 = 6'h2d == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_46_io_i_write_slot_T = 6'h2e == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_46_io_i_write_slot_T_2 = 6'h2e == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_46_io_i_write_slot_T_5 = 6'h2e == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_47_io_i_write_slot_T = 6'h2f == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_47_io_i_write_slot_T_2 = 6'h2f == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_47_io_i_write_slot_T_5 = 6'h2f == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_48_io_i_write_slot_T = 6'h30 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_48_io_i_write_slot_T_2 = 6'h30 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_48_io_i_write_slot_T_5 = 6'h30 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_49_io_i_write_slot_T = 6'h31 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_49_io_i_write_slot_T_2 = 6'h31 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_49_io_i_write_slot_T_5 = 6'h31 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_50_io_i_write_slot_T = 6'h32 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_50_io_i_write_slot_T_2 = 6'h32 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_50_io_i_write_slot_T_5 = 6'h32 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_51_io_i_write_slot_T = 6'h33 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_51_io_i_write_slot_T_2 = 6'h33 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_51_io_i_write_slot_T_5 = 6'h33 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_52_io_i_write_slot_T = 6'h34 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_52_io_i_write_slot_T_2 = 6'h34 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_52_io_i_write_slot_T_5 = 6'h34 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_53_io_i_write_slot_T = 6'h35 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_53_io_i_write_slot_T_2 = 6'h35 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_53_io_i_write_slot_T_5 = 6'h35 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_54_io_i_write_slot_T = 6'h36 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_54_io_i_write_slot_T_2 = 6'h36 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_54_io_i_write_slot_T_5 = 6'h36 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_55_io_i_write_slot_T = 6'h37 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_55_io_i_write_slot_T_2 = 6'h37 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_55_io_i_write_slot_T_5 = 6'h37 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_56_io_i_write_slot_T = 6'h38 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_56_io_i_write_slot_T_2 = 6'h38 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_56_io_i_write_slot_T_5 = 6'h38 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_57_io_i_write_slot_T = 6'h39 == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_57_io_i_write_slot_T_2 = 6'h39 == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_57_io_i_write_slot_T_5 = 6'h39 == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_58_io_i_write_slot_T = 6'h3a == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_58_io_i_write_slot_T_2 = 6'h3a == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_58_io_i_write_slot_T_5 = 6'h3a == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_59_io_i_write_slot_T = 6'h3b == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_59_io_i_write_slot_T_2 = 6'h3b == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_59_io_i_write_slot_T_5 = 6'h3b == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_60_io_i_write_slot_T = 6'h3c == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_60_io_i_write_slot_T_2 = 6'h3c == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_60_io_i_write_slot_T_5 = 6'h3c == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_61_io_i_write_slot_T = 6'h3d == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_61_io_i_write_slot_T_2 = 6'h3d == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_61_io_i_write_slot_T_5 = 6'h3d == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_62_io_i_write_slot_T = 6'h3e == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_62_io_i_write_slot_T_2 = 6'h3e == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_62_io_i_write_slot_T_5 = 6'h3e == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  wire  _reservation_station_63_io_i_write_slot_T = 6'h3f == write_idx1; // @[reservation_station.scala 118:14]
  wire  _reservation_station_63_io_i_write_slot_T_2 = 6'h3f == write_idx1 & write_idx1 != 6'h3f; // @[reservation_station.scala 118:29]
  wire  _reservation_station_63_io_i_write_slot_T_5 = 6'h3f == write_idx2 & write_idx2 != 6'h3f; // @[reservation_station.scala 119:29]
  Reservation_Station_Slot reservation_station_0 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_0_clock),
    .reset(reservation_station_0_reset),
    .io_o_valid(reservation_station_0_io_o_valid),
    .io_o_ready_to_issue(reservation_station_0_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_0_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_0_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_0_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_0_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_0_io_i_exception),
    .io_i_write_slot(reservation_station_0_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_0_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_0_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_0_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_0_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_0_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_0_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_0_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_0_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_0_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_0_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_0_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_0_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_0_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_0_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_0_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_0_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_0_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_0_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_0_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_0_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_0_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_0_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_0_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_0_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_0_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_0_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_0_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_0_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_0_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_0_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_0_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_0_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_0_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_0_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_0_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_0_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_0_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_0_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_0_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_0_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_0_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_0_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_0_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_0_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_0_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_0_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_0_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_0_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_0_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_0_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_0_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_0_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_0_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_0_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_0_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_0_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_0_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_0_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_0_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_0_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_0_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_0_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_0_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_1 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_1_clock),
    .reset(reservation_station_1_reset),
    .io_o_valid(reservation_station_1_io_o_valid),
    .io_o_ready_to_issue(reservation_station_1_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_1_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_1_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_1_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_1_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_1_io_i_exception),
    .io_i_write_slot(reservation_station_1_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_1_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_1_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_1_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_1_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_1_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_1_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_1_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_1_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_1_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_1_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_1_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_1_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_1_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_1_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_1_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_1_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_1_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_1_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_1_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_1_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_1_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_1_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_1_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_1_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_1_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_1_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_1_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_1_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_1_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_1_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_1_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_1_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_1_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_1_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_1_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_1_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_1_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_1_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_1_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_1_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_1_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_1_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_1_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_1_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_1_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_1_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_1_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_1_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_1_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_1_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_1_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_1_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_1_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_1_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_1_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_1_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_1_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_1_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_1_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_1_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_1_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_1_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_1_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_2 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_2_clock),
    .reset(reservation_station_2_reset),
    .io_o_valid(reservation_station_2_io_o_valid),
    .io_o_ready_to_issue(reservation_station_2_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_2_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_2_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_2_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_2_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_2_io_i_exception),
    .io_i_write_slot(reservation_station_2_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_2_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_2_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_2_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_2_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_2_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_2_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_2_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_2_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_2_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_2_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_2_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_2_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_2_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_2_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_2_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_2_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_2_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_2_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_2_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_2_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_2_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_2_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_2_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_2_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_2_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_2_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_2_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_2_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_2_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_2_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_2_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_2_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_2_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_2_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_2_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_2_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_2_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_2_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_2_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_2_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_2_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_2_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_2_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_2_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_2_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_2_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_2_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_2_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_2_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_2_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_2_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_2_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_2_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_2_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_2_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_2_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_2_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_2_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_2_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_2_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_2_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_2_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_2_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_3 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_3_clock),
    .reset(reservation_station_3_reset),
    .io_o_valid(reservation_station_3_io_o_valid),
    .io_o_ready_to_issue(reservation_station_3_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_3_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_3_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_3_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_3_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_3_io_i_exception),
    .io_i_write_slot(reservation_station_3_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_3_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_3_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_3_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_3_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_3_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_3_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_3_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_3_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_3_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_3_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_3_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_3_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_3_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_3_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_3_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_3_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_3_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_3_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_3_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_3_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_3_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_3_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_3_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_3_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_3_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_3_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_3_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_3_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_3_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_3_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_3_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_3_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_3_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_3_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_3_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_3_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_3_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_3_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_3_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_3_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_3_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_3_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_3_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_3_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_3_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_3_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_3_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_3_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_3_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_3_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_3_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_3_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_3_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_3_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_3_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_3_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_3_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_3_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_3_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_3_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_3_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_3_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_3_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_4 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_4_clock),
    .reset(reservation_station_4_reset),
    .io_o_valid(reservation_station_4_io_o_valid),
    .io_o_ready_to_issue(reservation_station_4_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_4_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_4_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_4_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_4_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_4_io_i_exception),
    .io_i_write_slot(reservation_station_4_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_4_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_4_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_4_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_4_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_4_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_4_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_4_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_4_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_4_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_4_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_4_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_4_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_4_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_4_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_4_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_4_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_4_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_4_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_4_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_4_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_4_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_4_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_4_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_4_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_4_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_4_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_4_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_4_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_4_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_4_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_4_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_4_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_4_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_4_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_4_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_4_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_4_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_4_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_4_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_4_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_4_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_4_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_4_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_4_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_4_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_4_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_4_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_4_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_4_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_4_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_4_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_4_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_4_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_4_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_4_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_4_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_4_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_4_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_4_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_4_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_4_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_4_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_4_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_5 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_5_clock),
    .reset(reservation_station_5_reset),
    .io_o_valid(reservation_station_5_io_o_valid),
    .io_o_ready_to_issue(reservation_station_5_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_5_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_5_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_5_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_5_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_5_io_i_exception),
    .io_i_write_slot(reservation_station_5_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_5_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_5_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_5_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_5_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_5_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_5_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_5_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_5_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_5_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_5_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_5_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_5_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_5_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_5_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_5_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_5_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_5_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_5_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_5_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_5_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_5_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_5_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_5_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_5_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_5_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_5_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_5_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_5_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_5_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_5_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_5_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_5_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_5_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_5_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_5_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_5_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_5_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_5_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_5_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_5_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_5_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_5_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_5_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_5_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_5_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_5_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_5_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_5_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_5_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_5_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_5_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_5_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_5_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_5_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_5_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_5_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_5_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_5_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_5_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_5_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_5_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_5_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_5_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_6 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_6_clock),
    .reset(reservation_station_6_reset),
    .io_o_valid(reservation_station_6_io_o_valid),
    .io_o_ready_to_issue(reservation_station_6_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_6_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_6_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_6_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_6_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_6_io_i_exception),
    .io_i_write_slot(reservation_station_6_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_6_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_6_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_6_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_6_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_6_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_6_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_6_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_6_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_6_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_6_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_6_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_6_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_6_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_6_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_6_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_6_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_6_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_6_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_6_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_6_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_6_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_6_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_6_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_6_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_6_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_6_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_6_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_6_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_6_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_6_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_6_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_6_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_6_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_6_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_6_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_6_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_6_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_6_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_6_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_6_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_6_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_6_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_6_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_6_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_6_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_6_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_6_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_6_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_6_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_6_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_6_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_6_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_6_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_6_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_6_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_6_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_6_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_6_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_6_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_6_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_6_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_6_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_6_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_7 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_7_clock),
    .reset(reservation_station_7_reset),
    .io_o_valid(reservation_station_7_io_o_valid),
    .io_o_ready_to_issue(reservation_station_7_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_7_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_7_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_7_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_7_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_7_io_i_exception),
    .io_i_write_slot(reservation_station_7_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_7_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_7_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_7_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_7_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_7_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_7_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_7_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_7_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_7_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_7_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_7_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_7_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_7_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_7_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_7_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_7_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_7_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_7_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_7_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_7_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_7_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_7_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_7_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_7_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_7_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_7_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_7_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_7_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_7_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_7_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_7_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_7_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_7_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_7_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_7_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_7_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_7_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_7_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_7_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_7_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_7_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_7_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_7_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_7_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_7_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_7_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_7_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_7_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_7_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_7_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_7_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_7_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_7_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_7_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_7_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_7_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_7_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_7_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_7_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_7_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_7_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_7_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_7_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_8 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_8_clock),
    .reset(reservation_station_8_reset),
    .io_o_valid(reservation_station_8_io_o_valid),
    .io_o_ready_to_issue(reservation_station_8_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_8_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_8_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_8_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_8_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_8_io_i_exception),
    .io_i_write_slot(reservation_station_8_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_8_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_8_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_8_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_8_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_8_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_8_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_8_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_8_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_8_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_8_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_8_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_8_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_8_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_8_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_8_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_8_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_8_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_8_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_8_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_8_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_8_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_8_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_8_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_8_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_8_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_8_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_8_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_8_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_8_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_8_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_8_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_8_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_8_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_8_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_8_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_8_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_8_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_8_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_8_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_8_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_8_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_8_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_8_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_8_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_8_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_8_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_8_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_8_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_8_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_8_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_8_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_8_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_8_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_8_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_8_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_8_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_8_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_8_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_8_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_8_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_8_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_8_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_8_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_9 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_9_clock),
    .reset(reservation_station_9_reset),
    .io_o_valid(reservation_station_9_io_o_valid),
    .io_o_ready_to_issue(reservation_station_9_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_9_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_9_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_9_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_9_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_9_io_i_exception),
    .io_i_write_slot(reservation_station_9_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_9_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_9_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_9_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_9_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_9_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_9_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_9_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_9_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_9_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_9_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_9_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_9_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_9_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_9_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_9_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_9_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_9_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_9_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_9_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_9_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_9_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_9_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_9_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_9_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_9_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_9_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_9_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_9_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_9_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_9_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_9_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_9_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_9_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_9_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_9_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_9_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_9_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_9_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_9_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_9_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_9_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_9_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_9_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_9_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_9_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_9_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_9_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_9_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_9_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_9_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_9_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_9_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_9_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_9_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_9_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_9_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_9_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_9_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_9_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_9_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_9_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_9_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_9_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_10 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_10_clock),
    .reset(reservation_station_10_reset),
    .io_o_valid(reservation_station_10_io_o_valid),
    .io_o_ready_to_issue(reservation_station_10_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_10_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_10_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_10_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_10_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_10_io_i_exception),
    .io_i_write_slot(reservation_station_10_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_10_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_10_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_10_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_10_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_10_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_10_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_10_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_10_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_10_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_10_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_10_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_10_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_10_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_10_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_10_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_10_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_10_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_10_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_10_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_10_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_10_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_10_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_10_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_10_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_10_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_10_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_10_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_10_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_10_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_10_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_10_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_10_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_10_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_10_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_10_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_10_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_10_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_10_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_10_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_10_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_10_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_10_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_10_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_10_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_10_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_10_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_10_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_10_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_10_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_10_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_10_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_10_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_10_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_10_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_10_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_10_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_10_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_10_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_10_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_10_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_10_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_10_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_10_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_11 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_11_clock),
    .reset(reservation_station_11_reset),
    .io_o_valid(reservation_station_11_io_o_valid),
    .io_o_ready_to_issue(reservation_station_11_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_11_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_11_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_11_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_11_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_11_io_i_exception),
    .io_i_write_slot(reservation_station_11_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_11_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_11_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_11_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_11_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_11_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_11_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_11_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_11_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_11_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_11_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_11_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_11_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_11_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_11_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_11_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_11_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_11_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_11_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_11_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_11_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_11_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_11_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_11_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_11_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_11_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_11_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_11_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_11_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_11_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_11_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_11_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_11_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_11_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_11_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_11_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_11_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_11_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_11_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_11_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_11_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_11_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_11_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_11_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_11_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_11_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_11_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_11_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_11_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_11_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_11_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_11_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_11_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_11_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_11_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_11_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_11_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_11_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_11_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_11_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_11_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_11_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_11_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_11_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_12 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_12_clock),
    .reset(reservation_station_12_reset),
    .io_o_valid(reservation_station_12_io_o_valid),
    .io_o_ready_to_issue(reservation_station_12_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_12_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_12_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_12_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_12_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_12_io_i_exception),
    .io_i_write_slot(reservation_station_12_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_12_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_12_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_12_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_12_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_12_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_12_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_12_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_12_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_12_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_12_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_12_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_12_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_12_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_12_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_12_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_12_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_12_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_12_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_12_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_12_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_12_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_12_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_12_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_12_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_12_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_12_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_12_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_12_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_12_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_12_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_12_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_12_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_12_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_12_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_12_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_12_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_12_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_12_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_12_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_12_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_12_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_12_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_12_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_12_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_12_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_12_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_12_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_12_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_12_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_12_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_12_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_12_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_12_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_12_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_12_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_12_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_12_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_12_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_12_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_12_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_12_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_12_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_12_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_13 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_13_clock),
    .reset(reservation_station_13_reset),
    .io_o_valid(reservation_station_13_io_o_valid),
    .io_o_ready_to_issue(reservation_station_13_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_13_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_13_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_13_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_13_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_13_io_i_exception),
    .io_i_write_slot(reservation_station_13_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_13_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_13_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_13_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_13_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_13_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_13_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_13_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_13_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_13_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_13_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_13_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_13_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_13_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_13_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_13_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_13_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_13_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_13_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_13_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_13_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_13_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_13_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_13_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_13_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_13_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_13_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_13_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_13_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_13_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_13_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_13_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_13_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_13_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_13_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_13_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_13_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_13_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_13_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_13_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_13_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_13_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_13_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_13_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_13_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_13_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_13_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_13_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_13_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_13_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_13_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_13_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_13_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_13_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_13_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_13_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_13_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_13_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_13_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_13_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_13_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_13_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_13_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_13_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_14 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_14_clock),
    .reset(reservation_station_14_reset),
    .io_o_valid(reservation_station_14_io_o_valid),
    .io_o_ready_to_issue(reservation_station_14_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_14_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_14_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_14_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_14_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_14_io_i_exception),
    .io_i_write_slot(reservation_station_14_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_14_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_14_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_14_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_14_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_14_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_14_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_14_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_14_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_14_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_14_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_14_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_14_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_14_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_14_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_14_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_14_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_14_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_14_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_14_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_14_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_14_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_14_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_14_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_14_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_14_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_14_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_14_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_14_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_14_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_14_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_14_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_14_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_14_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_14_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_14_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_14_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_14_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_14_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_14_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_14_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_14_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_14_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_14_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_14_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_14_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_14_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_14_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_14_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_14_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_14_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_14_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_14_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_14_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_14_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_14_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_14_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_14_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_14_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_14_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_14_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_14_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_14_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_14_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_15 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_15_clock),
    .reset(reservation_station_15_reset),
    .io_o_valid(reservation_station_15_io_o_valid),
    .io_o_ready_to_issue(reservation_station_15_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_15_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_15_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_15_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_15_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_15_io_i_exception),
    .io_i_write_slot(reservation_station_15_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_15_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_15_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_15_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_15_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_15_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_15_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_15_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_15_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_15_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_15_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_15_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_15_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_15_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_15_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_15_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_15_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_15_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_15_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_15_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_15_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_15_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_15_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_15_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_15_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_15_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_15_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_15_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_15_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_15_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_15_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_15_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_15_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_15_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_15_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_15_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_15_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_15_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_15_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_15_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_15_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_15_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_15_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_15_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_15_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_15_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_15_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_15_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_15_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_15_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_15_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_15_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_15_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_15_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_15_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_15_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_15_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_15_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_15_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_15_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_15_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_15_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_15_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_15_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_16 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_16_clock),
    .reset(reservation_station_16_reset),
    .io_o_valid(reservation_station_16_io_o_valid),
    .io_o_ready_to_issue(reservation_station_16_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_16_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_16_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_16_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_16_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_16_io_i_exception),
    .io_i_write_slot(reservation_station_16_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_16_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_16_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_16_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_16_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_16_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_16_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_16_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_16_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_16_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_16_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_16_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_16_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_16_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_16_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_16_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_16_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_16_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_16_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_16_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_16_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_16_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_16_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_16_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_16_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_16_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_16_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_16_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_16_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_16_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_16_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_16_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_16_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_16_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_16_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_16_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_16_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_16_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_16_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_16_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_16_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_16_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_16_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_16_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_16_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_16_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_16_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_16_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_16_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_16_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_16_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_16_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_16_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_16_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_16_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_16_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_16_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_16_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_16_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_16_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_16_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_16_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_16_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_16_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_17 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_17_clock),
    .reset(reservation_station_17_reset),
    .io_o_valid(reservation_station_17_io_o_valid),
    .io_o_ready_to_issue(reservation_station_17_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_17_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_17_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_17_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_17_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_17_io_i_exception),
    .io_i_write_slot(reservation_station_17_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_17_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_17_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_17_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_17_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_17_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_17_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_17_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_17_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_17_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_17_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_17_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_17_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_17_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_17_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_17_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_17_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_17_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_17_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_17_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_17_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_17_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_17_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_17_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_17_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_17_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_17_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_17_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_17_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_17_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_17_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_17_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_17_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_17_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_17_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_17_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_17_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_17_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_17_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_17_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_17_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_17_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_17_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_17_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_17_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_17_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_17_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_17_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_17_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_17_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_17_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_17_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_17_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_17_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_17_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_17_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_17_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_17_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_17_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_17_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_17_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_17_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_17_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_17_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_18 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_18_clock),
    .reset(reservation_station_18_reset),
    .io_o_valid(reservation_station_18_io_o_valid),
    .io_o_ready_to_issue(reservation_station_18_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_18_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_18_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_18_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_18_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_18_io_i_exception),
    .io_i_write_slot(reservation_station_18_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_18_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_18_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_18_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_18_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_18_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_18_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_18_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_18_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_18_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_18_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_18_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_18_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_18_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_18_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_18_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_18_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_18_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_18_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_18_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_18_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_18_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_18_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_18_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_18_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_18_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_18_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_18_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_18_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_18_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_18_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_18_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_18_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_18_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_18_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_18_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_18_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_18_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_18_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_18_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_18_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_18_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_18_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_18_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_18_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_18_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_18_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_18_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_18_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_18_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_18_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_18_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_18_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_18_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_18_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_18_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_18_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_18_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_18_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_18_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_18_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_18_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_18_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_18_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_19 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_19_clock),
    .reset(reservation_station_19_reset),
    .io_o_valid(reservation_station_19_io_o_valid),
    .io_o_ready_to_issue(reservation_station_19_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_19_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_19_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_19_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_19_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_19_io_i_exception),
    .io_i_write_slot(reservation_station_19_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_19_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_19_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_19_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_19_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_19_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_19_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_19_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_19_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_19_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_19_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_19_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_19_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_19_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_19_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_19_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_19_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_19_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_19_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_19_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_19_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_19_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_19_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_19_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_19_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_19_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_19_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_19_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_19_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_19_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_19_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_19_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_19_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_19_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_19_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_19_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_19_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_19_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_19_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_19_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_19_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_19_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_19_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_19_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_19_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_19_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_19_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_19_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_19_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_19_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_19_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_19_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_19_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_19_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_19_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_19_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_19_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_19_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_19_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_19_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_19_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_19_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_19_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_19_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_20 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_20_clock),
    .reset(reservation_station_20_reset),
    .io_o_valid(reservation_station_20_io_o_valid),
    .io_o_ready_to_issue(reservation_station_20_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_20_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_20_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_20_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_20_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_20_io_i_exception),
    .io_i_write_slot(reservation_station_20_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_20_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_20_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_20_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_20_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_20_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_20_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_20_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_20_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_20_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_20_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_20_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_20_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_20_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_20_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_20_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_20_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_20_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_20_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_20_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_20_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_20_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_20_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_20_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_20_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_20_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_20_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_20_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_20_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_20_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_20_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_20_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_20_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_20_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_20_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_20_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_20_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_20_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_20_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_20_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_20_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_20_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_20_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_20_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_20_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_20_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_20_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_20_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_20_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_20_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_20_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_20_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_20_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_20_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_20_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_20_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_20_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_20_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_20_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_20_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_20_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_20_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_20_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_20_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_21 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_21_clock),
    .reset(reservation_station_21_reset),
    .io_o_valid(reservation_station_21_io_o_valid),
    .io_o_ready_to_issue(reservation_station_21_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_21_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_21_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_21_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_21_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_21_io_i_exception),
    .io_i_write_slot(reservation_station_21_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_21_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_21_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_21_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_21_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_21_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_21_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_21_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_21_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_21_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_21_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_21_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_21_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_21_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_21_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_21_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_21_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_21_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_21_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_21_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_21_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_21_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_21_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_21_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_21_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_21_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_21_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_21_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_21_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_21_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_21_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_21_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_21_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_21_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_21_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_21_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_21_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_21_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_21_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_21_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_21_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_21_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_21_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_21_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_21_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_21_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_21_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_21_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_21_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_21_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_21_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_21_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_21_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_21_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_21_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_21_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_21_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_21_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_21_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_21_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_21_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_21_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_21_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_21_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_22 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_22_clock),
    .reset(reservation_station_22_reset),
    .io_o_valid(reservation_station_22_io_o_valid),
    .io_o_ready_to_issue(reservation_station_22_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_22_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_22_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_22_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_22_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_22_io_i_exception),
    .io_i_write_slot(reservation_station_22_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_22_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_22_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_22_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_22_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_22_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_22_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_22_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_22_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_22_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_22_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_22_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_22_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_22_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_22_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_22_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_22_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_22_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_22_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_22_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_22_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_22_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_22_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_22_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_22_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_22_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_22_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_22_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_22_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_22_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_22_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_22_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_22_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_22_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_22_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_22_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_22_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_22_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_22_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_22_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_22_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_22_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_22_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_22_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_22_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_22_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_22_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_22_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_22_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_22_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_22_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_22_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_22_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_22_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_22_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_22_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_22_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_22_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_22_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_22_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_22_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_22_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_22_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_22_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_23 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_23_clock),
    .reset(reservation_station_23_reset),
    .io_o_valid(reservation_station_23_io_o_valid),
    .io_o_ready_to_issue(reservation_station_23_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_23_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_23_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_23_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_23_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_23_io_i_exception),
    .io_i_write_slot(reservation_station_23_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_23_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_23_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_23_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_23_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_23_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_23_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_23_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_23_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_23_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_23_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_23_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_23_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_23_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_23_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_23_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_23_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_23_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_23_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_23_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_23_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_23_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_23_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_23_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_23_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_23_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_23_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_23_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_23_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_23_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_23_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_23_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_23_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_23_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_23_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_23_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_23_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_23_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_23_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_23_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_23_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_23_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_23_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_23_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_23_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_23_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_23_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_23_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_23_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_23_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_23_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_23_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_23_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_23_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_23_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_23_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_23_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_23_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_23_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_23_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_23_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_23_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_23_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_23_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_24 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_24_clock),
    .reset(reservation_station_24_reset),
    .io_o_valid(reservation_station_24_io_o_valid),
    .io_o_ready_to_issue(reservation_station_24_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_24_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_24_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_24_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_24_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_24_io_i_exception),
    .io_i_write_slot(reservation_station_24_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_24_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_24_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_24_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_24_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_24_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_24_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_24_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_24_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_24_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_24_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_24_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_24_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_24_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_24_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_24_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_24_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_24_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_24_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_24_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_24_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_24_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_24_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_24_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_24_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_24_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_24_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_24_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_24_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_24_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_24_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_24_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_24_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_24_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_24_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_24_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_24_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_24_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_24_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_24_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_24_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_24_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_24_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_24_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_24_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_24_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_24_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_24_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_24_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_24_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_24_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_24_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_24_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_24_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_24_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_24_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_24_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_24_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_24_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_24_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_24_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_24_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_24_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_24_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_25 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_25_clock),
    .reset(reservation_station_25_reset),
    .io_o_valid(reservation_station_25_io_o_valid),
    .io_o_ready_to_issue(reservation_station_25_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_25_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_25_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_25_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_25_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_25_io_i_exception),
    .io_i_write_slot(reservation_station_25_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_25_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_25_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_25_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_25_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_25_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_25_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_25_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_25_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_25_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_25_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_25_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_25_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_25_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_25_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_25_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_25_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_25_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_25_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_25_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_25_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_25_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_25_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_25_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_25_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_25_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_25_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_25_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_25_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_25_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_25_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_25_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_25_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_25_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_25_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_25_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_25_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_25_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_25_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_25_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_25_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_25_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_25_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_25_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_25_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_25_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_25_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_25_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_25_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_25_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_25_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_25_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_25_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_25_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_25_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_25_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_25_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_25_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_25_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_25_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_25_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_25_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_25_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_25_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_26 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_26_clock),
    .reset(reservation_station_26_reset),
    .io_o_valid(reservation_station_26_io_o_valid),
    .io_o_ready_to_issue(reservation_station_26_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_26_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_26_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_26_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_26_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_26_io_i_exception),
    .io_i_write_slot(reservation_station_26_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_26_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_26_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_26_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_26_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_26_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_26_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_26_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_26_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_26_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_26_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_26_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_26_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_26_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_26_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_26_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_26_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_26_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_26_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_26_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_26_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_26_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_26_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_26_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_26_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_26_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_26_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_26_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_26_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_26_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_26_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_26_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_26_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_26_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_26_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_26_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_26_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_26_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_26_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_26_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_26_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_26_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_26_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_26_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_26_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_26_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_26_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_26_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_26_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_26_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_26_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_26_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_26_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_26_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_26_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_26_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_26_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_26_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_26_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_26_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_26_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_26_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_26_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_26_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_27 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_27_clock),
    .reset(reservation_station_27_reset),
    .io_o_valid(reservation_station_27_io_o_valid),
    .io_o_ready_to_issue(reservation_station_27_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_27_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_27_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_27_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_27_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_27_io_i_exception),
    .io_i_write_slot(reservation_station_27_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_27_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_27_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_27_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_27_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_27_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_27_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_27_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_27_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_27_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_27_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_27_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_27_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_27_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_27_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_27_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_27_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_27_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_27_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_27_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_27_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_27_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_27_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_27_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_27_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_27_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_27_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_27_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_27_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_27_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_27_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_27_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_27_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_27_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_27_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_27_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_27_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_27_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_27_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_27_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_27_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_27_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_27_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_27_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_27_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_27_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_27_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_27_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_27_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_27_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_27_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_27_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_27_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_27_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_27_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_27_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_27_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_27_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_27_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_27_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_27_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_27_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_27_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_27_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_28 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_28_clock),
    .reset(reservation_station_28_reset),
    .io_o_valid(reservation_station_28_io_o_valid),
    .io_o_ready_to_issue(reservation_station_28_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_28_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_28_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_28_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_28_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_28_io_i_exception),
    .io_i_write_slot(reservation_station_28_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_28_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_28_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_28_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_28_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_28_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_28_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_28_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_28_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_28_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_28_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_28_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_28_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_28_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_28_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_28_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_28_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_28_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_28_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_28_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_28_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_28_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_28_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_28_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_28_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_28_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_28_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_28_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_28_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_28_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_28_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_28_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_28_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_28_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_28_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_28_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_28_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_28_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_28_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_28_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_28_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_28_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_28_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_28_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_28_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_28_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_28_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_28_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_28_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_28_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_28_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_28_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_28_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_28_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_28_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_28_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_28_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_28_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_28_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_28_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_28_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_28_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_28_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_28_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_29 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_29_clock),
    .reset(reservation_station_29_reset),
    .io_o_valid(reservation_station_29_io_o_valid),
    .io_o_ready_to_issue(reservation_station_29_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_29_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_29_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_29_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_29_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_29_io_i_exception),
    .io_i_write_slot(reservation_station_29_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_29_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_29_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_29_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_29_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_29_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_29_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_29_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_29_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_29_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_29_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_29_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_29_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_29_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_29_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_29_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_29_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_29_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_29_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_29_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_29_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_29_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_29_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_29_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_29_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_29_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_29_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_29_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_29_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_29_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_29_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_29_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_29_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_29_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_29_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_29_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_29_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_29_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_29_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_29_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_29_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_29_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_29_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_29_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_29_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_29_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_29_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_29_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_29_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_29_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_29_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_29_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_29_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_29_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_29_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_29_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_29_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_29_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_29_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_29_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_29_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_29_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_29_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_29_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_30 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_30_clock),
    .reset(reservation_station_30_reset),
    .io_o_valid(reservation_station_30_io_o_valid),
    .io_o_ready_to_issue(reservation_station_30_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_30_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_30_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_30_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_30_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_30_io_i_exception),
    .io_i_write_slot(reservation_station_30_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_30_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_30_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_30_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_30_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_30_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_30_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_30_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_30_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_30_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_30_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_30_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_30_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_30_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_30_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_30_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_30_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_30_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_30_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_30_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_30_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_30_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_30_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_30_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_30_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_30_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_30_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_30_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_30_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_30_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_30_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_30_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_30_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_30_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_30_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_30_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_30_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_30_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_30_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_30_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_30_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_30_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_30_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_30_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_30_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_30_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_30_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_30_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_30_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_30_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_30_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_30_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_30_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_30_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_30_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_30_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_30_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_30_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_30_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_30_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_30_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_30_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_30_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_30_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_31 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_31_clock),
    .reset(reservation_station_31_reset),
    .io_o_valid(reservation_station_31_io_o_valid),
    .io_o_ready_to_issue(reservation_station_31_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_31_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_31_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_31_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_31_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_31_io_i_exception),
    .io_i_write_slot(reservation_station_31_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_31_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_31_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_31_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_31_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_31_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_31_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_31_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_31_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_31_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_31_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_31_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_31_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_31_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_31_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_31_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_31_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_31_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_31_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_31_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_31_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_31_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_31_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_31_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_31_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_31_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_31_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_31_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_31_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_31_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_31_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_31_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_31_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_31_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_31_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_31_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_31_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_31_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_31_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_31_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_31_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_31_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_31_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_31_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_31_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_31_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_31_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_31_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_31_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_31_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_31_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_31_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_31_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_31_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_31_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_31_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_31_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_31_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_31_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_31_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_31_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_31_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_31_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_31_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_32 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_32_clock),
    .reset(reservation_station_32_reset),
    .io_o_valid(reservation_station_32_io_o_valid),
    .io_o_ready_to_issue(reservation_station_32_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_32_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_32_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_32_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_32_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_32_io_i_exception),
    .io_i_write_slot(reservation_station_32_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_32_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_32_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_32_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_32_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_32_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_32_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_32_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_32_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_32_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_32_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_32_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_32_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_32_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_32_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_32_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_32_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_32_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_32_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_32_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_32_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_32_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_32_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_32_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_32_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_32_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_32_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_32_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_32_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_32_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_32_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_32_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_32_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_32_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_32_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_32_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_32_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_32_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_32_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_32_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_32_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_32_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_32_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_32_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_32_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_32_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_32_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_32_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_32_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_32_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_32_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_32_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_32_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_32_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_32_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_32_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_32_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_32_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_32_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_32_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_32_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_32_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_32_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_32_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_33 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_33_clock),
    .reset(reservation_station_33_reset),
    .io_o_valid(reservation_station_33_io_o_valid),
    .io_o_ready_to_issue(reservation_station_33_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_33_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_33_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_33_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_33_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_33_io_i_exception),
    .io_i_write_slot(reservation_station_33_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_33_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_33_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_33_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_33_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_33_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_33_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_33_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_33_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_33_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_33_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_33_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_33_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_33_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_33_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_33_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_33_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_33_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_33_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_33_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_33_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_33_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_33_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_33_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_33_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_33_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_33_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_33_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_33_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_33_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_33_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_33_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_33_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_33_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_33_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_33_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_33_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_33_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_33_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_33_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_33_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_33_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_33_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_33_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_33_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_33_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_33_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_33_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_33_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_33_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_33_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_33_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_33_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_33_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_33_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_33_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_33_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_33_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_33_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_33_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_33_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_33_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_33_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_33_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_34 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_34_clock),
    .reset(reservation_station_34_reset),
    .io_o_valid(reservation_station_34_io_o_valid),
    .io_o_ready_to_issue(reservation_station_34_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_34_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_34_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_34_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_34_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_34_io_i_exception),
    .io_i_write_slot(reservation_station_34_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_34_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_34_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_34_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_34_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_34_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_34_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_34_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_34_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_34_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_34_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_34_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_34_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_34_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_34_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_34_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_34_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_34_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_34_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_34_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_34_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_34_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_34_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_34_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_34_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_34_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_34_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_34_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_34_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_34_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_34_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_34_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_34_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_34_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_34_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_34_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_34_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_34_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_34_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_34_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_34_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_34_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_34_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_34_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_34_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_34_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_34_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_34_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_34_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_34_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_34_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_34_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_34_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_34_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_34_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_34_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_34_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_34_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_34_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_34_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_34_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_34_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_34_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_34_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_35 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_35_clock),
    .reset(reservation_station_35_reset),
    .io_o_valid(reservation_station_35_io_o_valid),
    .io_o_ready_to_issue(reservation_station_35_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_35_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_35_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_35_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_35_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_35_io_i_exception),
    .io_i_write_slot(reservation_station_35_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_35_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_35_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_35_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_35_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_35_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_35_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_35_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_35_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_35_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_35_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_35_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_35_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_35_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_35_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_35_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_35_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_35_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_35_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_35_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_35_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_35_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_35_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_35_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_35_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_35_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_35_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_35_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_35_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_35_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_35_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_35_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_35_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_35_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_35_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_35_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_35_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_35_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_35_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_35_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_35_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_35_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_35_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_35_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_35_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_35_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_35_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_35_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_35_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_35_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_35_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_35_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_35_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_35_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_35_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_35_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_35_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_35_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_35_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_35_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_35_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_35_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_35_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_35_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_36 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_36_clock),
    .reset(reservation_station_36_reset),
    .io_o_valid(reservation_station_36_io_o_valid),
    .io_o_ready_to_issue(reservation_station_36_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_36_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_36_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_36_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_36_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_36_io_i_exception),
    .io_i_write_slot(reservation_station_36_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_36_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_36_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_36_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_36_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_36_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_36_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_36_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_36_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_36_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_36_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_36_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_36_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_36_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_36_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_36_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_36_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_36_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_36_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_36_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_36_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_36_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_36_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_36_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_36_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_36_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_36_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_36_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_36_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_36_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_36_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_36_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_36_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_36_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_36_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_36_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_36_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_36_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_36_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_36_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_36_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_36_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_36_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_36_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_36_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_36_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_36_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_36_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_36_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_36_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_36_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_36_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_36_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_36_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_36_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_36_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_36_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_36_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_36_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_36_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_36_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_36_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_36_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_36_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_37 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_37_clock),
    .reset(reservation_station_37_reset),
    .io_o_valid(reservation_station_37_io_o_valid),
    .io_o_ready_to_issue(reservation_station_37_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_37_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_37_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_37_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_37_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_37_io_i_exception),
    .io_i_write_slot(reservation_station_37_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_37_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_37_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_37_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_37_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_37_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_37_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_37_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_37_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_37_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_37_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_37_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_37_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_37_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_37_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_37_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_37_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_37_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_37_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_37_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_37_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_37_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_37_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_37_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_37_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_37_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_37_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_37_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_37_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_37_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_37_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_37_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_37_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_37_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_37_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_37_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_37_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_37_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_37_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_37_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_37_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_37_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_37_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_37_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_37_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_37_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_37_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_37_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_37_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_37_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_37_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_37_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_37_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_37_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_37_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_37_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_37_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_37_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_37_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_37_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_37_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_37_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_37_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_37_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_38 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_38_clock),
    .reset(reservation_station_38_reset),
    .io_o_valid(reservation_station_38_io_o_valid),
    .io_o_ready_to_issue(reservation_station_38_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_38_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_38_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_38_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_38_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_38_io_i_exception),
    .io_i_write_slot(reservation_station_38_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_38_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_38_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_38_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_38_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_38_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_38_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_38_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_38_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_38_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_38_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_38_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_38_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_38_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_38_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_38_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_38_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_38_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_38_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_38_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_38_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_38_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_38_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_38_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_38_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_38_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_38_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_38_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_38_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_38_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_38_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_38_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_38_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_38_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_38_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_38_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_38_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_38_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_38_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_38_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_38_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_38_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_38_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_38_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_38_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_38_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_38_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_38_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_38_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_38_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_38_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_38_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_38_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_38_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_38_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_38_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_38_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_38_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_38_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_38_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_38_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_38_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_38_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_38_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_39 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_39_clock),
    .reset(reservation_station_39_reset),
    .io_o_valid(reservation_station_39_io_o_valid),
    .io_o_ready_to_issue(reservation_station_39_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_39_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_39_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_39_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_39_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_39_io_i_exception),
    .io_i_write_slot(reservation_station_39_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_39_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_39_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_39_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_39_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_39_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_39_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_39_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_39_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_39_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_39_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_39_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_39_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_39_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_39_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_39_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_39_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_39_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_39_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_39_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_39_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_39_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_39_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_39_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_39_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_39_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_39_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_39_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_39_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_39_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_39_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_39_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_39_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_39_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_39_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_39_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_39_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_39_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_39_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_39_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_39_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_39_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_39_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_39_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_39_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_39_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_39_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_39_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_39_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_39_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_39_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_39_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_39_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_39_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_39_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_39_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_39_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_39_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_39_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_39_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_39_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_39_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_39_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_39_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_40 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_40_clock),
    .reset(reservation_station_40_reset),
    .io_o_valid(reservation_station_40_io_o_valid),
    .io_o_ready_to_issue(reservation_station_40_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_40_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_40_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_40_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_40_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_40_io_i_exception),
    .io_i_write_slot(reservation_station_40_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_40_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_40_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_40_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_40_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_40_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_40_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_40_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_40_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_40_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_40_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_40_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_40_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_40_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_40_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_40_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_40_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_40_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_40_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_40_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_40_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_40_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_40_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_40_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_40_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_40_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_40_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_40_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_40_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_40_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_40_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_40_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_40_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_40_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_40_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_40_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_40_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_40_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_40_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_40_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_40_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_40_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_40_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_40_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_40_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_40_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_40_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_40_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_40_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_40_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_40_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_40_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_40_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_40_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_40_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_40_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_40_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_40_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_40_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_40_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_40_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_40_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_40_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_40_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_41 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_41_clock),
    .reset(reservation_station_41_reset),
    .io_o_valid(reservation_station_41_io_o_valid),
    .io_o_ready_to_issue(reservation_station_41_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_41_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_41_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_41_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_41_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_41_io_i_exception),
    .io_i_write_slot(reservation_station_41_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_41_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_41_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_41_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_41_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_41_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_41_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_41_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_41_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_41_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_41_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_41_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_41_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_41_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_41_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_41_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_41_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_41_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_41_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_41_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_41_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_41_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_41_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_41_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_41_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_41_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_41_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_41_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_41_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_41_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_41_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_41_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_41_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_41_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_41_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_41_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_41_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_41_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_41_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_41_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_41_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_41_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_41_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_41_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_41_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_41_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_41_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_41_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_41_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_41_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_41_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_41_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_41_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_41_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_41_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_41_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_41_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_41_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_41_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_41_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_41_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_41_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_41_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_41_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_42 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_42_clock),
    .reset(reservation_station_42_reset),
    .io_o_valid(reservation_station_42_io_o_valid),
    .io_o_ready_to_issue(reservation_station_42_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_42_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_42_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_42_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_42_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_42_io_i_exception),
    .io_i_write_slot(reservation_station_42_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_42_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_42_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_42_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_42_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_42_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_42_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_42_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_42_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_42_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_42_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_42_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_42_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_42_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_42_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_42_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_42_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_42_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_42_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_42_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_42_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_42_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_42_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_42_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_42_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_42_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_42_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_42_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_42_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_42_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_42_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_42_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_42_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_42_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_42_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_42_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_42_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_42_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_42_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_42_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_42_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_42_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_42_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_42_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_42_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_42_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_42_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_42_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_42_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_42_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_42_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_42_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_42_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_42_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_42_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_42_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_42_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_42_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_42_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_42_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_42_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_42_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_42_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_42_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_43 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_43_clock),
    .reset(reservation_station_43_reset),
    .io_o_valid(reservation_station_43_io_o_valid),
    .io_o_ready_to_issue(reservation_station_43_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_43_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_43_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_43_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_43_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_43_io_i_exception),
    .io_i_write_slot(reservation_station_43_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_43_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_43_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_43_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_43_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_43_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_43_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_43_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_43_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_43_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_43_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_43_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_43_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_43_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_43_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_43_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_43_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_43_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_43_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_43_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_43_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_43_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_43_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_43_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_43_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_43_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_43_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_43_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_43_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_43_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_43_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_43_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_43_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_43_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_43_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_43_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_43_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_43_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_43_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_43_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_43_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_43_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_43_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_43_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_43_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_43_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_43_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_43_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_43_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_43_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_43_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_43_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_43_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_43_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_43_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_43_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_43_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_43_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_43_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_43_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_43_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_43_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_43_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_43_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_44 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_44_clock),
    .reset(reservation_station_44_reset),
    .io_o_valid(reservation_station_44_io_o_valid),
    .io_o_ready_to_issue(reservation_station_44_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_44_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_44_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_44_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_44_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_44_io_i_exception),
    .io_i_write_slot(reservation_station_44_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_44_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_44_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_44_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_44_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_44_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_44_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_44_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_44_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_44_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_44_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_44_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_44_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_44_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_44_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_44_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_44_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_44_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_44_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_44_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_44_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_44_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_44_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_44_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_44_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_44_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_44_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_44_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_44_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_44_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_44_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_44_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_44_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_44_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_44_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_44_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_44_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_44_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_44_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_44_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_44_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_44_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_44_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_44_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_44_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_44_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_44_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_44_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_44_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_44_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_44_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_44_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_44_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_44_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_44_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_44_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_44_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_44_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_44_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_44_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_44_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_44_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_44_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_44_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_45 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_45_clock),
    .reset(reservation_station_45_reset),
    .io_o_valid(reservation_station_45_io_o_valid),
    .io_o_ready_to_issue(reservation_station_45_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_45_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_45_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_45_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_45_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_45_io_i_exception),
    .io_i_write_slot(reservation_station_45_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_45_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_45_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_45_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_45_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_45_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_45_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_45_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_45_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_45_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_45_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_45_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_45_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_45_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_45_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_45_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_45_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_45_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_45_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_45_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_45_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_45_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_45_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_45_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_45_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_45_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_45_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_45_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_45_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_45_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_45_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_45_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_45_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_45_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_45_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_45_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_45_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_45_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_45_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_45_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_45_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_45_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_45_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_45_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_45_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_45_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_45_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_45_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_45_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_45_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_45_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_45_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_45_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_45_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_45_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_45_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_45_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_45_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_45_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_45_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_45_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_45_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_45_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_45_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_46 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_46_clock),
    .reset(reservation_station_46_reset),
    .io_o_valid(reservation_station_46_io_o_valid),
    .io_o_ready_to_issue(reservation_station_46_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_46_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_46_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_46_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_46_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_46_io_i_exception),
    .io_i_write_slot(reservation_station_46_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_46_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_46_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_46_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_46_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_46_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_46_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_46_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_46_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_46_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_46_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_46_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_46_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_46_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_46_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_46_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_46_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_46_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_46_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_46_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_46_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_46_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_46_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_46_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_46_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_46_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_46_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_46_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_46_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_46_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_46_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_46_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_46_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_46_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_46_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_46_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_46_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_46_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_46_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_46_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_46_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_46_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_46_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_46_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_46_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_46_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_46_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_46_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_46_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_46_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_46_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_46_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_46_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_46_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_46_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_46_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_46_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_46_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_46_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_46_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_46_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_46_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_46_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_46_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_47 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_47_clock),
    .reset(reservation_station_47_reset),
    .io_o_valid(reservation_station_47_io_o_valid),
    .io_o_ready_to_issue(reservation_station_47_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_47_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_47_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_47_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_47_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_47_io_i_exception),
    .io_i_write_slot(reservation_station_47_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_47_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_47_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_47_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_47_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_47_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_47_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_47_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_47_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_47_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_47_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_47_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_47_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_47_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_47_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_47_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_47_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_47_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_47_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_47_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_47_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_47_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_47_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_47_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_47_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_47_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_47_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_47_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_47_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_47_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_47_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_47_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_47_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_47_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_47_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_47_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_47_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_47_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_47_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_47_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_47_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_47_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_47_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_47_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_47_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_47_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_47_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_47_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_47_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_47_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_47_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_47_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_47_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_47_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_47_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_47_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_47_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_47_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_47_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_47_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_47_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_47_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_47_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_47_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_48 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_48_clock),
    .reset(reservation_station_48_reset),
    .io_o_valid(reservation_station_48_io_o_valid),
    .io_o_ready_to_issue(reservation_station_48_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_48_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_48_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_48_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_48_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_48_io_i_exception),
    .io_i_write_slot(reservation_station_48_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_48_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_48_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_48_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_48_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_48_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_48_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_48_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_48_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_48_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_48_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_48_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_48_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_48_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_48_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_48_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_48_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_48_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_48_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_48_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_48_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_48_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_48_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_48_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_48_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_48_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_48_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_48_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_48_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_48_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_48_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_48_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_48_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_48_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_48_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_48_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_48_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_48_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_48_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_48_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_48_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_48_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_48_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_48_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_48_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_48_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_48_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_48_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_48_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_48_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_48_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_48_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_48_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_48_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_48_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_48_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_48_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_48_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_48_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_48_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_48_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_48_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_48_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_48_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_49 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_49_clock),
    .reset(reservation_station_49_reset),
    .io_o_valid(reservation_station_49_io_o_valid),
    .io_o_ready_to_issue(reservation_station_49_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_49_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_49_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_49_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_49_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_49_io_i_exception),
    .io_i_write_slot(reservation_station_49_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_49_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_49_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_49_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_49_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_49_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_49_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_49_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_49_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_49_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_49_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_49_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_49_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_49_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_49_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_49_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_49_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_49_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_49_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_49_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_49_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_49_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_49_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_49_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_49_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_49_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_49_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_49_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_49_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_49_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_49_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_49_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_49_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_49_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_49_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_49_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_49_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_49_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_49_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_49_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_49_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_49_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_49_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_49_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_49_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_49_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_49_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_49_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_49_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_49_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_49_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_49_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_49_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_49_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_49_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_49_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_49_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_49_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_49_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_49_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_49_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_49_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_49_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_49_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_50 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_50_clock),
    .reset(reservation_station_50_reset),
    .io_o_valid(reservation_station_50_io_o_valid),
    .io_o_ready_to_issue(reservation_station_50_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_50_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_50_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_50_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_50_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_50_io_i_exception),
    .io_i_write_slot(reservation_station_50_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_50_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_50_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_50_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_50_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_50_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_50_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_50_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_50_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_50_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_50_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_50_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_50_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_50_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_50_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_50_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_50_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_50_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_50_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_50_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_50_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_50_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_50_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_50_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_50_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_50_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_50_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_50_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_50_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_50_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_50_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_50_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_50_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_50_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_50_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_50_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_50_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_50_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_50_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_50_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_50_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_50_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_50_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_50_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_50_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_50_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_50_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_50_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_50_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_50_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_50_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_50_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_50_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_50_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_50_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_50_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_50_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_50_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_50_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_50_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_50_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_50_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_50_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_50_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_51 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_51_clock),
    .reset(reservation_station_51_reset),
    .io_o_valid(reservation_station_51_io_o_valid),
    .io_o_ready_to_issue(reservation_station_51_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_51_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_51_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_51_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_51_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_51_io_i_exception),
    .io_i_write_slot(reservation_station_51_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_51_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_51_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_51_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_51_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_51_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_51_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_51_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_51_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_51_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_51_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_51_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_51_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_51_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_51_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_51_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_51_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_51_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_51_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_51_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_51_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_51_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_51_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_51_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_51_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_51_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_51_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_51_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_51_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_51_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_51_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_51_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_51_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_51_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_51_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_51_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_51_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_51_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_51_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_51_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_51_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_51_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_51_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_51_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_51_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_51_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_51_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_51_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_51_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_51_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_51_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_51_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_51_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_51_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_51_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_51_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_51_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_51_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_51_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_51_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_51_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_51_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_51_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_51_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_52 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_52_clock),
    .reset(reservation_station_52_reset),
    .io_o_valid(reservation_station_52_io_o_valid),
    .io_o_ready_to_issue(reservation_station_52_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_52_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_52_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_52_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_52_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_52_io_i_exception),
    .io_i_write_slot(reservation_station_52_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_52_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_52_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_52_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_52_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_52_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_52_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_52_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_52_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_52_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_52_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_52_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_52_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_52_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_52_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_52_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_52_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_52_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_52_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_52_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_52_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_52_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_52_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_52_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_52_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_52_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_52_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_52_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_52_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_52_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_52_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_52_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_52_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_52_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_52_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_52_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_52_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_52_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_52_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_52_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_52_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_52_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_52_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_52_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_52_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_52_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_52_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_52_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_52_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_52_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_52_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_52_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_52_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_52_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_52_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_52_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_52_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_52_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_52_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_52_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_52_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_52_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_52_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_52_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_53 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_53_clock),
    .reset(reservation_station_53_reset),
    .io_o_valid(reservation_station_53_io_o_valid),
    .io_o_ready_to_issue(reservation_station_53_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_53_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_53_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_53_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_53_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_53_io_i_exception),
    .io_i_write_slot(reservation_station_53_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_53_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_53_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_53_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_53_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_53_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_53_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_53_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_53_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_53_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_53_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_53_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_53_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_53_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_53_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_53_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_53_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_53_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_53_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_53_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_53_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_53_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_53_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_53_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_53_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_53_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_53_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_53_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_53_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_53_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_53_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_53_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_53_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_53_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_53_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_53_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_53_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_53_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_53_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_53_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_53_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_53_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_53_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_53_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_53_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_53_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_53_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_53_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_53_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_53_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_53_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_53_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_53_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_53_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_53_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_53_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_53_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_53_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_53_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_53_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_53_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_53_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_53_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_53_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_54 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_54_clock),
    .reset(reservation_station_54_reset),
    .io_o_valid(reservation_station_54_io_o_valid),
    .io_o_ready_to_issue(reservation_station_54_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_54_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_54_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_54_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_54_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_54_io_i_exception),
    .io_i_write_slot(reservation_station_54_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_54_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_54_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_54_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_54_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_54_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_54_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_54_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_54_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_54_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_54_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_54_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_54_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_54_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_54_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_54_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_54_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_54_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_54_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_54_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_54_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_54_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_54_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_54_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_54_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_54_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_54_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_54_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_54_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_54_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_54_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_54_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_54_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_54_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_54_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_54_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_54_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_54_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_54_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_54_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_54_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_54_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_54_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_54_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_54_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_54_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_54_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_54_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_54_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_54_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_54_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_54_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_54_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_54_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_54_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_54_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_54_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_54_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_54_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_54_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_54_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_54_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_54_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_54_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_55 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_55_clock),
    .reset(reservation_station_55_reset),
    .io_o_valid(reservation_station_55_io_o_valid),
    .io_o_ready_to_issue(reservation_station_55_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_55_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_55_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_55_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_55_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_55_io_i_exception),
    .io_i_write_slot(reservation_station_55_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_55_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_55_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_55_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_55_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_55_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_55_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_55_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_55_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_55_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_55_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_55_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_55_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_55_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_55_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_55_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_55_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_55_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_55_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_55_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_55_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_55_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_55_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_55_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_55_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_55_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_55_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_55_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_55_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_55_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_55_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_55_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_55_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_55_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_55_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_55_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_55_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_55_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_55_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_55_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_55_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_55_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_55_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_55_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_55_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_55_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_55_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_55_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_55_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_55_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_55_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_55_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_55_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_55_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_55_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_55_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_55_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_55_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_55_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_55_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_55_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_55_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_55_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_55_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_56 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_56_clock),
    .reset(reservation_station_56_reset),
    .io_o_valid(reservation_station_56_io_o_valid),
    .io_o_ready_to_issue(reservation_station_56_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_56_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_56_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_56_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_56_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_56_io_i_exception),
    .io_i_write_slot(reservation_station_56_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_56_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_56_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_56_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_56_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_56_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_56_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_56_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_56_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_56_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_56_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_56_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_56_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_56_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_56_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_56_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_56_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_56_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_56_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_56_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_56_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_56_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_56_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_56_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_56_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_56_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_56_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_56_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_56_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_56_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_56_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_56_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_56_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_56_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_56_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_56_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_56_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_56_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_56_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_56_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_56_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_56_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_56_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_56_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_56_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_56_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_56_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_56_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_56_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_56_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_56_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_56_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_56_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_56_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_56_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_56_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_56_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_56_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_56_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_56_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_56_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_56_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_56_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_56_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_57 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_57_clock),
    .reset(reservation_station_57_reset),
    .io_o_valid(reservation_station_57_io_o_valid),
    .io_o_ready_to_issue(reservation_station_57_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_57_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_57_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_57_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_57_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_57_io_i_exception),
    .io_i_write_slot(reservation_station_57_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_57_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_57_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_57_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_57_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_57_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_57_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_57_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_57_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_57_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_57_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_57_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_57_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_57_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_57_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_57_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_57_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_57_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_57_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_57_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_57_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_57_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_57_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_57_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_57_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_57_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_57_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_57_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_57_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_57_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_57_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_57_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_57_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_57_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_57_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_57_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_57_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_57_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_57_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_57_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_57_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_57_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_57_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_57_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_57_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_57_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_57_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_57_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_57_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_57_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_57_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_57_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_57_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_57_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_57_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_57_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_57_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_57_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_57_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_57_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_57_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_57_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_57_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_57_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_58 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_58_clock),
    .reset(reservation_station_58_reset),
    .io_o_valid(reservation_station_58_io_o_valid),
    .io_o_ready_to_issue(reservation_station_58_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_58_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_58_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_58_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_58_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_58_io_i_exception),
    .io_i_write_slot(reservation_station_58_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_58_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_58_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_58_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_58_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_58_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_58_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_58_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_58_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_58_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_58_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_58_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_58_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_58_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_58_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_58_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_58_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_58_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_58_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_58_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_58_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_58_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_58_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_58_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_58_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_58_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_58_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_58_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_58_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_58_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_58_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_58_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_58_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_58_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_58_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_58_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_58_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_58_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_58_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_58_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_58_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_58_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_58_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_58_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_58_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_58_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_58_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_58_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_58_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_58_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_58_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_58_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_58_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_58_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_58_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_58_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_58_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_58_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_58_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_58_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_58_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_58_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_58_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_58_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_59 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_59_clock),
    .reset(reservation_station_59_reset),
    .io_o_valid(reservation_station_59_io_o_valid),
    .io_o_ready_to_issue(reservation_station_59_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_59_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_59_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_59_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_59_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_59_io_i_exception),
    .io_i_write_slot(reservation_station_59_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_59_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_59_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_59_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_59_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_59_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_59_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_59_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_59_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_59_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_59_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_59_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_59_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_59_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_59_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_59_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_59_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_59_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_59_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_59_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_59_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_59_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_59_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_59_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_59_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_59_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_59_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_59_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_59_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_59_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_59_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_59_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_59_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_59_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_59_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_59_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_59_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_59_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_59_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_59_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_59_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_59_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_59_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_59_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_59_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_59_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_59_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_59_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_59_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_59_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_59_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_59_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_59_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_59_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_59_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_59_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_59_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_59_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_59_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_59_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_59_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_59_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_59_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_59_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_60 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_60_clock),
    .reset(reservation_station_60_reset),
    .io_o_valid(reservation_station_60_io_o_valid),
    .io_o_ready_to_issue(reservation_station_60_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_60_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_60_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_60_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_60_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_60_io_i_exception),
    .io_i_write_slot(reservation_station_60_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_60_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_60_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_60_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_60_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_60_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_60_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_60_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_60_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_60_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_60_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_60_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_60_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_60_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_60_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_60_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_60_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_60_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_60_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_60_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_60_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_60_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_60_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_60_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_60_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_60_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_60_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_60_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_60_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_60_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_60_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_60_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_60_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_60_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_60_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_60_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_60_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_60_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_60_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_60_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_60_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_60_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_60_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_60_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_60_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_60_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_60_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_60_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_60_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_60_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_60_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_60_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_60_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_60_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_60_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_60_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_60_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_60_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_60_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_60_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_60_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_60_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_60_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_60_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_61 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_61_clock),
    .reset(reservation_station_61_reset),
    .io_o_valid(reservation_station_61_io_o_valid),
    .io_o_ready_to_issue(reservation_station_61_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_61_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_61_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_61_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_61_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_61_io_i_exception),
    .io_i_write_slot(reservation_station_61_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_61_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_61_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_61_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_61_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_61_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_61_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_61_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_61_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_61_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_61_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_61_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_61_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_61_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_61_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_61_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_61_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_61_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_61_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_61_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_61_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_61_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_61_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_61_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_61_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_61_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_61_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_61_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_61_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_61_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_61_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_61_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_61_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_61_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_61_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_61_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_61_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_61_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_61_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_61_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_61_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_61_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_61_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_61_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_61_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_61_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_61_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_61_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_61_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_61_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_61_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_61_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_61_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_61_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_61_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_61_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_61_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_61_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_61_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_61_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_61_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_61_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_61_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_61_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_62 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_62_clock),
    .reset(reservation_station_62_reset),
    .io_o_valid(reservation_station_62_io_o_valid),
    .io_o_ready_to_issue(reservation_station_62_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_62_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_62_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_62_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_62_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_62_io_i_exception),
    .io_i_write_slot(reservation_station_62_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_62_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_62_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_62_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_62_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_62_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_62_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_62_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_62_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_62_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_62_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_62_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_62_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_62_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_62_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_62_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_62_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_62_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_62_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_62_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_62_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_62_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_62_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_62_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_62_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_62_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_62_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_62_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_62_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_62_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_62_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_62_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_62_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_62_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_62_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_62_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_62_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_62_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_62_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_62_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_62_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_62_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_62_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_62_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_62_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_62_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_62_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_62_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_62_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_62_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_62_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_62_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_62_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_62_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_62_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_62_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_62_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_62_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_62_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_62_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_62_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_62_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_62_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_62_io_i_ROB_first_entry)
  );
  Reservation_Station_Slot reservation_station_63 ( // @[reservation_station.scala 38:51]
    .clock(reservation_station_63_clock),
    .reset(reservation_station_63_reset),
    .io_o_valid(reservation_station_63_io_o_valid),
    .io_o_ready_to_issue(reservation_station_63_io_o_ready_to_issue),
    .io_i_issue_granted(reservation_station_63_io_i_issue_granted),
    .io_i_branch_resolve_pack_valid(reservation_station_63_io_i_branch_resolve_pack_valid),
    .io_i_branch_resolve_pack_mispred(reservation_station_63_io_i_branch_resolve_pack_mispred),
    .io_i_branch_resolve_pack_rob_idx(reservation_station_63_io_i_branch_resolve_pack_rob_idx),
    .io_i_exception(reservation_station_63_io_i_exception),
    .io_i_write_slot(reservation_station_63_io_i_write_slot),
    .io_i_wakeup_port(reservation_station_63_io_i_wakeup_port),
    .io_i_uop_valid(reservation_station_63_io_i_uop_valid),
    .io_i_uop_pc(reservation_station_63_io_i_uop_pc),
    .io_i_uop_inst(reservation_station_63_io_i_uop_inst),
    .io_i_uop_func_code(reservation_station_63_io_i_uop_func_code),
    .io_i_uop_branch_predict_pack_valid(reservation_station_63_io_i_uop_branch_predict_pack_valid),
    .io_i_uop_branch_predict_pack_target(reservation_station_63_io_i_uop_branch_predict_pack_target),
    .io_i_uop_branch_predict_pack_branch_type(reservation_station_63_io_i_uop_branch_predict_pack_branch_type),
    .io_i_uop_branch_predict_pack_select(reservation_station_63_io_i_uop_branch_predict_pack_select),
    .io_i_uop_branch_predict_pack_taken(reservation_station_63_io_i_uop_branch_predict_pack_taken),
    .io_i_uop_phy_dst(reservation_station_63_io_i_uop_phy_dst),
    .io_i_uop_stale_dst(reservation_station_63_io_i_uop_stale_dst),
    .io_i_uop_arch_dst(reservation_station_63_io_i_uop_arch_dst),
    .io_i_uop_inst_type(reservation_station_63_io_i_uop_inst_type),
    .io_i_uop_regWen(reservation_station_63_io_i_uop_regWen),
    .io_i_uop_src1_valid(reservation_station_63_io_i_uop_src1_valid),
    .io_i_uop_phy_rs1(reservation_station_63_io_i_uop_phy_rs1),
    .io_i_uop_arch_rs1(reservation_station_63_io_i_uop_arch_rs1),
    .io_i_uop_src2_valid(reservation_station_63_io_i_uop_src2_valid),
    .io_i_uop_phy_rs2(reservation_station_63_io_i_uop_phy_rs2),
    .io_i_uop_arch_rs2(reservation_station_63_io_i_uop_arch_rs2),
    .io_i_uop_rob_idx(reservation_station_63_io_i_uop_rob_idx),
    .io_i_uop_imm(reservation_station_63_io_i_uop_imm),
    .io_i_uop_src1_value(reservation_station_63_io_i_uop_src1_value),
    .io_i_uop_src2_value(reservation_station_63_io_i_uop_src2_value),
    .io_i_uop_op1_sel(reservation_station_63_io_i_uop_op1_sel),
    .io_i_uop_op2_sel(reservation_station_63_io_i_uop_op2_sel),
    .io_i_uop_alu_sel(reservation_station_63_io_i_uop_alu_sel),
    .io_i_uop_branch_type(reservation_station_63_io_i_uop_branch_type),
    .io_i_uop_mem_type(reservation_station_63_io_i_uop_mem_type),
    .io_o_uop_pc(reservation_station_63_io_o_uop_pc),
    .io_o_uop_inst(reservation_station_63_io_o_uop_inst),
    .io_o_uop_func_code(reservation_station_63_io_o_uop_func_code),
    .io_o_uop_branch_predict_pack_valid(reservation_station_63_io_o_uop_branch_predict_pack_valid),
    .io_o_uop_branch_predict_pack_target(reservation_station_63_io_o_uop_branch_predict_pack_target),
    .io_o_uop_branch_predict_pack_branch_type(reservation_station_63_io_o_uop_branch_predict_pack_branch_type),
    .io_o_uop_branch_predict_pack_select(reservation_station_63_io_o_uop_branch_predict_pack_select),
    .io_o_uop_branch_predict_pack_taken(reservation_station_63_io_o_uop_branch_predict_pack_taken),
    .io_o_uop_phy_dst(reservation_station_63_io_o_uop_phy_dst),
    .io_o_uop_stale_dst(reservation_station_63_io_o_uop_stale_dst),
    .io_o_uop_arch_dst(reservation_station_63_io_o_uop_arch_dst),
    .io_o_uop_inst_type(reservation_station_63_io_o_uop_inst_type),
    .io_o_uop_regWen(reservation_station_63_io_o_uop_regWen),
    .io_o_uop_src1_valid(reservation_station_63_io_o_uop_src1_valid),
    .io_o_uop_phy_rs1(reservation_station_63_io_o_uop_phy_rs1),
    .io_o_uop_arch_rs1(reservation_station_63_io_o_uop_arch_rs1),
    .io_o_uop_src2_valid(reservation_station_63_io_o_uop_src2_valid),
    .io_o_uop_phy_rs2(reservation_station_63_io_o_uop_phy_rs2),
    .io_o_uop_arch_rs2(reservation_station_63_io_o_uop_arch_rs2),
    .io_o_uop_rob_idx(reservation_station_63_io_o_uop_rob_idx),
    .io_o_uop_imm(reservation_station_63_io_o_uop_imm),
    .io_o_uop_src1_value(reservation_station_63_io_o_uop_src1_value),
    .io_o_uop_src2_value(reservation_station_63_io_o_uop_src2_value),
    .io_o_uop_op1_sel(reservation_station_63_io_o_uop_op1_sel),
    .io_o_uop_op2_sel(reservation_station_63_io_o_uop_op2_sel),
    .io_o_uop_alu_sel(reservation_station_63_io_o_uop_alu_sel),
    .io_o_uop_branch_type(reservation_station_63_io_o_uop_branch_type),
    .io_o_uop_mem_type(reservation_station_63_io_o_uop_mem_type),
    .io_i_exe_dst1(reservation_station_63_io_i_exe_dst1),
    .io_i_exe_dst2(reservation_station_63_io_i_exe_dst2),
    .io_i_exe_value1(reservation_station_63_io_i_exe_value1),
    .io_i_exe_value2(reservation_station_63_io_i_exe_value2),
    .io_i_ROB_first_entry(reservation_station_63_io_i_ROB_first_entry)
  );
  assign io_o_issue_packs_0_valid = issue_num == 2'h1 | issue_num == 2'h2; // @[reservation_station.scala 93:38]
  assign io_o_issue_packs_0_pc = _issue1_func_code_T ? reservation_station_0_io_o_uop_pc : _io_o_issue_packs_0_T_126_pc; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_inst = _issue1_func_code_T ? reservation_station_0_io_o_uop_inst :
    _io_o_issue_packs_0_T_126_inst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_func_code = _issue1_func_code_T ? reservation_station_0_io_o_uop_func_code :
    _io_o_issue_packs_0_T_126_func_code; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_valid = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_0_T_126_branch_predict_pack_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_target = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_0_T_126_branch_predict_pack_target; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_branch_type = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_0_T_126_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_select = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_0_T_126_branch_predict_pack_select; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_predict_pack_taken = _issue1_func_code_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_0_T_126_branch_predict_pack_taken; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_dst :
    _io_o_issue_packs_0_T_126_phy_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_stale_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_stale_dst :
    _io_o_issue_packs_0_T_126_stale_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_dst = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_dst :
    _io_o_issue_packs_0_T_126_arch_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_inst_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_inst_type :
    _io_o_issue_packs_0_T_126_inst_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_regWen = _issue1_func_code_T ? reservation_station_0_io_o_uop_regWen :
    _io_o_issue_packs_0_T_126_regWen; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src1_valid = _issue1_func_code_T ? reservation_station_0_io_o_uop_src1_valid :
    _io_o_issue_packs_0_T_126_src1_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_rs1 = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_rs1 :
    _io_o_issue_packs_0_T_126_phy_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_rs1 = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_rs1 :
    _io_o_issue_packs_0_T_126_arch_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src2_valid = _issue1_func_code_T ? reservation_station_0_io_o_uop_src2_valid :
    _io_o_issue_packs_0_T_126_src2_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_phy_rs2 = _issue1_func_code_T ? reservation_station_0_io_o_uop_phy_rs2 :
    _io_o_issue_packs_0_T_126_phy_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_arch_rs2 = _issue1_func_code_T ? reservation_station_0_io_o_uop_arch_rs2 :
    _io_o_issue_packs_0_T_126_arch_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_rob_idx = _issue1_func_code_T ? reservation_station_0_io_o_uop_rob_idx :
    _io_o_issue_packs_0_T_126_rob_idx; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_imm = _issue1_func_code_T ? reservation_station_0_io_o_uop_imm :
    _io_o_issue_packs_0_T_126_imm; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src1_value = _issue1_func_code_T ? reservation_station_0_io_o_uop_src1_value :
    _io_o_issue_packs_0_T_126_src1_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_src2_value = _issue1_func_code_T ? reservation_station_0_io_o_uop_src2_value :
    _io_o_issue_packs_0_T_126_src2_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_op1_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_op1_sel :
    _io_o_issue_packs_0_T_126_op1_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_op2_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_op2_sel :
    _io_o_issue_packs_0_T_126_op2_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_alu_sel = _issue1_func_code_T ? reservation_station_0_io_o_uop_alu_sel :
    _io_o_issue_packs_0_T_126_alu_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_branch_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_branch_type :
    _io_o_issue_packs_0_T_126_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_0_mem_type = _issue1_func_code_T ? reservation_station_0_io_o_uop_mem_type :
    _io_o_issue_packs_0_T_126_mem_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_valid = issue_num == 2'h2; // @[reservation_station.scala 94:31]
  assign io_o_issue_packs_1_pc = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_pc :
    _io_o_issue_packs_1_T_126_pc; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_inst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_inst :
    _io_o_issue_packs_1_T_126_inst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_func_code = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_func_code :
    _io_o_issue_packs_1_T_126_func_code; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_valid = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_valid : _io_o_issue_packs_1_T_126_branch_predict_pack_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_target = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_target : _io_o_issue_packs_1_T_126_branch_predict_pack_target; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_branch_type = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_branch_type :
    _io_o_issue_packs_1_T_126_branch_predict_pack_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_select = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_select : _io_o_issue_packs_1_T_126_branch_predict_pack_select; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_predict_pack_taken = _io_o_issue_packs_1_T ?
    reservation_station_0_io_o_uop_branch_predict_pack_taken : _io_o_issue_packs_1_T_126_branch_predict_pack_taken; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_dst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_phy_dst :
    _io_o_issue_packs_1_T_126_phy_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_stale_dst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_stale_dst :
    _io_o_issue_packs_1_T_126_stale_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_dst = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_arch_dst :
    _io_o_issue_packs_1_T_126_arch_dst; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_inst_type = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_inst_type :
    _io_o_issue_packs_1_T_126_inst_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_regWen = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_regWen :
    _io_o_issue_packs_1_T_126_regWen; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src1_valid = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src1_valid :
    _io_o_issue_packs_1_T_126_src1_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_rs1 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_phy_rs1 :
    _io_o_issue_packs_1_T_126_phy_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_rs1 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_arch_rs1 :
    _io_o_issue_packs_1_T_126_arch_rs1; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src2_valid = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src2_valid :
    _io_o_issue_packs_1_T_126_src2_valid; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_phy_rs2 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_phy_rs2 :
    _io_o_issue_packs_1_T_126_phy_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_arch_rs2 = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_arch_rs2 :
    _io_o_issue_packs_1_T_126_arch_rs2; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_rob_idx = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_rob_idx :
    _io_o_issue_packs_1_T_126_rob_idx; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_imm = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_imm :
    _io_o_issue_packs_1_T_126_imm; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src1_value = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src1_value :
    _io_o_issue_packs_1_T_126_src1_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_src2_value = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_src2_value :
    _io_o_issue_packs_1_T_126_src2_value; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_op1_sel = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_op1_sel :
    _io_o_issue_packs_1_T_126_op1_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_op2_sel = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_op2_sel :
    _io_o_issue_packs_1_T_126_op2_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_alu_sel = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_alu_sel :
    _io_o_issue_packs_1_T_126_alu_sel; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_branch_type = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_branch_type :
    _io_o_issue_packs_1_T_126_branch_type; // @[Mux.scala 101:16]
  assign io_o_issue_packs_1_mem_type = _io_o_issue_packs_1_T ? reservation_station_0_io_o_uop_mem_type :
    _io_o_issue_packs_1_T_126_mem_type; // @[Mux.scala 101:16]
  assign io_o_full = _write_num_T | _write_num_T_1; // @[reservation_station.scala 104:38]
  assign reservation_station_0_clock = clock;
  assign reservation_station_0_reset = reset;
  assign reservation_station_0_io_i_issue_granted = (_issue1_func_code_T | _io_o_issue_packs_1_T) & ~(io_i_exception |
    io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_0_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_0_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_0_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_0_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_0_io_i_write_slot = _reservation_station_0_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_0_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_0_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_0_io_i_uop_valid = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_pc = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_inst = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_func_code = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_target = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_branch_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_select = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_predict_pack_taken = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_phy_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_stale_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_arch_dst = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_inst_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_regWen = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src1_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_phy_rs1 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_arch_rs1 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src2_valid = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_phy_rs2 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_arch_rs2 = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_rob_idx = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_imm = _reservation_station_0_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src1_value = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_src2_value = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_op1_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_op2_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_alu_sel = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_branch_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_uop_mem_type = _reservation_station_0_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_0_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_0_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_0_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_0_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_0_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_1_clock = clock;
  assign reservation_station_1_reset = reset;
  assign reservation_station_1_io_i_issue_granted = (_issue1_func_code_T_1 | _io_o_issue_packs_1_T_1) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_1_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_1_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_1_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_1_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_1_io_i_write_slot = _reservation_station_1_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_1_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_1_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_1_io_i_uop_valid = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_pc = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_inst = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_func_code = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_target = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_branch_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_select = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_predict_pack_taken = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_phy_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_stale_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_arch_dst = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_inst_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_regWen = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src1_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_phy_rs1 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_arch_rs1 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src2_valid = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_phy_rs2 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_arch_rs2 = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_rob_idx = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_imm = _reservation_station_1_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src1_value = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_src2_value = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_op1_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_op2_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_alu_sel = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_branch_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_uop_mem_type = _reservation_station_1_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_1_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_1_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_1_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_1_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_1_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_2_clock = clock;
  assign reservation_station_2_reset = reset;
  assign reservation_station_2_io_i_issue_granted = (_issue1_func_code_T_2 | _io_o_issue_packs_1_T_2) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_2_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_2_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_2_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_2_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_2_io_i_write_slot = _reservation_station_2_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_2_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_2_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_2_io_i_uop_valid = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_pc = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_inst = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_func_code = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_target = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_branch_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_select = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_predict_pack_taken = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_phy_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_stale_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_arch_dst = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_inst_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_regWen = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src1_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_phy_rs1 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_arch_rs1 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src2_valid = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_phy_rs2 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_arch_rs2 = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_rob_idx = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_imm = _reservation_station_2_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src1_value = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_src2_value = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_op1_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_op2_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_alu_sel = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_branch_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_uop_mem_type = _reservation_station_2_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_2_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_2_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_2_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_2_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_2_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_3_clock = clock;
  assign reservation_station_3_reset = reset;
  assign reservation_station_3_io_i_issue_granted = (_issue1_func_code_T_3 | _io_o_issue_packs_1_T_3) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_3_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_3_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_3_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_3_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_3_io_i_write_slot = _reservation_station_3_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_3_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_3_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_3_io_i_uop_valid = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_pc = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_inst = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_func_code = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_target = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_branch_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_select = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_predict_pack_taken = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_phy_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_stale_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_arch_dst = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_inst_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_regWen = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src1_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_phy_rs1 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_arch_rs1 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src2_valid = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_phy_rs2 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_arch_rs2 = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_rob_idx = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_imm = _reservation_station_3_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src1_value = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_src2_value = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_op1_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_op2_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_alu_sel = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_branch_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_uop_mem_type = _reservation_station_3_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_3_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_3_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_3_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_3_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_3_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_4_clock = clock;
  assign reservation_station_4_reset = reset;
  assign reservation_station_4_io_i_issue_granted = (_issue1_func_code_T_4 | _io_o_issue_packs_1_T_4) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_4_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_4_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_4_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_4_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_4_io_i_write_slot = _reservation_station_4_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_4_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_4_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_4_io_i_uop_valid = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_pc = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_inst = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_func_code = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_target = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_branch_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_select = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_predict_pack_taken = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_phy_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_stale_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_arch_dst = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_inst_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_regWen = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src1_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_phy_rs1 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_arch_rs1 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src2_valid = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_phy_rs2 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_arch_rs2 = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_rob_idx = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_imm = _reservation_station_4_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src1_value = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_src2_value = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_op1_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_op2_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_alu_sel = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_branch_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_uop_mem_type = _reservation_station_4_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_4_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_4_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_4_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_4_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_4_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_5_clock = clock;
  assign reservation_station_5_reset = reset;
  assign reservation_station_5_io_i_issue_granted = (_issue1_func_code_T_5 | _io_o_issue_packs_1_T_5) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_5_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_5_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_5_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_5_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_5_io_i_write_slot = _reservation_station_5_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_5_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_5_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_5_io_i_uop_valid = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_pc = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_inst = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_func_code = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_target = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_branch_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_select = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_predict_pack_taken = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_phy_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_stale_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_arch_dst = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_inst_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_regWen = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src1_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_phy_rs1 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_arch_rs1 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src2_valid = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_phy_rs2 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_arch_rs2 = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_rob_idx = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_imm = _reservation_station_5_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src1_value = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_src2_value = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_op1_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_op2_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_alu_sel = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_branch_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_uop_mem_type = _reservation_station_5_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_5_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_5_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_5_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_5_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_5_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_6_clock = clock;
  assign reservation_station_6_reset = reset;
  assign reservation_station_6_io_i_issue_granted = (_issue1_func_code_T_6 | _io_o_issue_packs_1_T_6) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_6_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_6_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_6_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_6_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_6_io_i_write_slot = _reservation_station_6_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_6_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_6_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_6_io_i_uop_valid = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_pc = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_inst = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_func_code = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_target = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_branch_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_select = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_predict_pack_taken = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_phy_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_stale_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_arch_dst = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_inst_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_regWen = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src1_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_phy_rs1 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_arch_rs1 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src2_valid = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_phy_rs2 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_arch_rs2 = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_rob_idx = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_imm = _reservation_station_6_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src1_value = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_src2_value = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_op1_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_op2_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_alu_sel = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_branch_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_uop_mem_type = _reservation_station_6_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_6_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_6_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_6_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_6_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_6_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_7_clock = clock;
  assign reservation_station_7_reset = reset;
  assign reservation_station_7_io_i_issue_granted = (_issue1_func_code_T_7 | _io_o_issue_packs_1_T_7) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_7_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_7_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_7_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_7_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_7_io_i_write_slot = _reservation_station_7_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_7_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_7_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_7_io_i_uop_valid = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_pc = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_inst = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_func_code = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_target = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_branch_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_select = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_predict_pack_taken = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_phy_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_stale_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_arch_dst = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_inst_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_regWen = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src1_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_phy_rs1 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_arch_rs1 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src2_valid = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_phy_rs2 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_arch_rs2 = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_rob_idx = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_imm = _reservation_station_7_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src1_value = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_src2_value = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_op1_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_op2_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_alu_sel = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_branch_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_uop_mem_type = _reservation_station_7_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_7_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_7_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_7_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_7_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_7_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_8_clock = clock;
  assign reservation_station_8_reset = reset;
  assign reservation_station_8_io_i_issue_granted = (_issue1_func_code_T_8 | _io_o_issue_packs_1_T_8) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_8_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_8_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_8_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_8_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_8_io_i_write_slot = _reservation_station_8_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_8_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_8_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_8_io_i_uop_valid = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_pc = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_inst = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_func_code = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_target = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_branch_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_select = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_predict_pack_taken = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_phy_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_stale_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_arch_dst = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_inst_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_regWen = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src1_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_phy_rs1 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_arch_rs1 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src2_valid = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_phy_rs2 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_arch_rs2 = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_rob_idx = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_imm = _reservation_station_8_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src1_value = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_src2_value = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_op1_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_op2_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_alu_sel = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_branch_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_uop_mem_type = _reservation_station_8_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_8_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_8_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_8_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_8_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_8_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_9_clock = clock;
  assign reservation_station_9_reset = reset;
  assign reservation_station_9_io_i_issue_granted = (_issue1_func_code_T_9 | _io_o_issue_packs_1_T_9) & ~(io_i_exception
     | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_9_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_9_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_9_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_9_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_9_io_i_write_slot = _reservation_station_9_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_9_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_9_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_9_io_i_uop_valid = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_pc = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_inst = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_inst :
    io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_func_code = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_target = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_branch_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_select = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_predict_pack_taken = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_phy_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_stale_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_arch_dst = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_inst_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_regWen = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_regWen
     : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src1_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_phy_rs1 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_arch_rs1 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src2_valid = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_phy_rs2 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_arch_rs2 = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_rob_idx = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_imm = _reservation_station_9_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src1_value = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_src2_value = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_op1_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_op2_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_alu_sel = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_branch_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_uop_mem_type = _reservation_station_9_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_9_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_9_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20 ?
    io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_9_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_9_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_9_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_10_clock = clock;
  assign reservation_station_10_reset = reset;
  assign reservation_station_10_io_i_issue_granted = (_issue1_func_code_T_10 | _io_o_issue_packs_1_T_10) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_10_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_10_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_10_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_10_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_10_io_i_write_slot = _reservation_station_10_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_10_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_10_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_10_io_i_uop_valid = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_pc = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_inst = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_func_code = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_target = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_branch_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_select = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_predict_pack_taken = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_phy_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_stale_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_arch_dst = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_inst_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_regWen = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src1_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_phy_rs1 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_arch_rs1 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src2_valid = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_phy_rs2 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_arch_rs2 = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_rob_idx = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_imm = _reservation_station_10_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src1_value = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_src2_value = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_op1_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_op2_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_alu_sel = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_branch_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_uop_mem_type = _reservation_station_10_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_10_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_10_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_10_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_10_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_10_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_11_clock = clock;
  assign reservation_station_11_reset = reset;
  assign reservation_station_11_io_i_issue_granted = (_issue1_func_code_T_11 | _io_o_issue_packs_1_T_11) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_11_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_11_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_11_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_11_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_11_io_i_write_slot = _reservation_station_11_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_11_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_11_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_11_io_i_uop_valid = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_pc = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_inst = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_func_code = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_target = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_branch_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_select = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_predict_pack_taken = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_phy_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_stale_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_arch_dst = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_inst_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_regWen = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src1_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_phy_rs1 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_arch_rs1 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src2_valid = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_phy_rs2 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_arch_rs2 = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_rob_idx = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_imm = _reservation_station_11_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src1_value = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_src2_value = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_op1_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_op2_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_alu_sel = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_branch_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_uop_mem_type = _reservation_station_11_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_11_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_11_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_11_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_11_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_11_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_12_clock = clock;
  assign reservation_station_12_reset = reset;
  assign reservation_station_12_io_i_issue_granted = (_issue1_func_code_T_12 | _io_o_issue_packs_1_T_12) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_12_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_12_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_12_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_12_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_12_io_i_write_slot = _reservation_station_12_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_12_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_12_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_12_io_i_uop_valid = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_pc = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_inst = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_func_code = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_target = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_branch_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_select = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_predict_pack_taken = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_phy_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_stale_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_arch_dst = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_inst_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_regWen = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src1_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_phy_rs1 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_arch_rs1 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src2_valid = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_phy_rs2 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_arch_rs2 = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_rob_idx = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_imm = _reservation_station_12_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src1_value = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_src2_value = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_op1_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_op2_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_alu_sel = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_branch_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_uop_mem_type = _reservation_station_12_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_12_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_12_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_12_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_12_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_12_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_13_clock = clock;
  assign reservation_station_13_reset = reset;
  assign reservation_station_13_io_i_issue_granted = (_issue1_func_code_T_13 | _io_o_issue_packs_1_T_13) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_13_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_13_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_13_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_13_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_13_io_i_write_slot = _reservation_station_13_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_13_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_13_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_13_io_i_uop_valid = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_pc = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_inst = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_func_code = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_target = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_branch_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_select = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_predict_pack_taken = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_phy_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_stale_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_arch_dst = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_inst_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_regWen = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src1_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_phy_rs1 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_arch_rs1 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src2_valid = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_phy_rs2 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_arch_rs2 = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_rob_idx = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_imm = _reservation_station_13_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src1_value = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_src2_value = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_op1_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_op2_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_alu_sel = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_branch_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_uop_mem_type = _reservation_station_13_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_13_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_13_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_13_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_13_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_13_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_14_clock = clock;
  assign reservation_station_14_reset = reset;
  assign reservation_station_14_io_i_issue_granted = (_issue1_func_code_T_14 | _io_o_issue_packs_1_T_14) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_14_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_14_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_14_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_14_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_14_io_i_write_slot = _reservation_station_14_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_14_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_14_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_14_io_i_uop_valid = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_pc = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_inst = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_func_code = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_target = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_branch_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_select = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_predict_pack_taken = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_phy_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_stale_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_arch_dst = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_inst_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_regWen = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src1_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_phy_rs1 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_arch_rs1 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src2_valid = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_phy_rs2 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_arch_rs2 = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_rob_idx = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_imm = _reservation_station_14_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src1_value = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_src2_value = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_op1_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_op2_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_alu_sel = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_branch_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_uop_mem_type = _reservation_station_14_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_14_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_14_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_14_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_14_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_14_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_15_clock = clock;
  assign reservation_station_15_reset = reset;
  assign reservation_station_15_io_i_issue_granted = (_issue1_func_code_T_15 | _io_o_issue_packs_1_T_15) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_15_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_15_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_15_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_15_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_15_io_i_write_slot = _reservation_station_15_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_15_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_15_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_15_io_i_uop_valid = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_pc = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_inst = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_func_code = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_target = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_branch_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_select = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_predict_pack_taken = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_phy_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_stale_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_arch_dst = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_inst_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_regWen = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src1_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_phy_rs1 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_arch_rs1 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src2_valid = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_phy_rs2 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_arch_rs2 = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_rob_idx = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_imm = _reservation_station_15_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src1_value = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_src2_value = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_op1_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_op2_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_alu_sel = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_branch_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_uop_mem_type = _reservation_station_15_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_15_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_15_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_15_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_15_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_15_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_16_clock = clock;
  assign reservation_station_16_reset = reset;
  assign reservation_station_16_io_i_issue_granted = (_issue1_func_code_T_16 | _io_o_issue_packs_1_T_16) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_16_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_16_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_16_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_16_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_16_io_i_write_slot = _reservation_station_16_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_16_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_16_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_16_io_i_uop_valid = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_pc = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_inst = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_func_code = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_target = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_branch_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_select = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_predict_pack_taken = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_phy_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_stale_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_arch_dst = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_inst_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_regWen = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src1_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_phy_rs1 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_arch_rs1 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src2_valid = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_phy_rs2 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_arch_rs2 = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_rob_idx = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_imm = _reservation_station_16_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src1_value = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_src2_value = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_op1_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_op2_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_alu_sel = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_branch_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_uop_mem_type = _reservation_station_16_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_16_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_16_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_16_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_16_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_16_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_17_clock = clock;
  assign reservation_station_17_reset = reset;
  assign reservation_station_17_io_i_issue_granted = (_issue1_func_code_T_17 | _io_o_issue_packs_1_T_17) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_17_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_17_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_17_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_17_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_17_io_i_write_slot = _reservation_station_17_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_17_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_17_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_17_io_i_uop_valid = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_pc = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_inst = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_func_code = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_target = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_branch_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_select = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_predict_pack_taken = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_phy_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_stale_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_arch_dst = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_inst_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_regWen = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src1_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_phy_rs1 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_arch_rs1 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src2_valid = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_phy_rs2 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_arch_rs2 = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_rob_idx = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_imm = _reservation_station_17_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src1_value = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_src2_value = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_op1_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_op2_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_alu_sel = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_branch_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_uop_mem_type = _reservation_station_17_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_17_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_17_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_17_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_17_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_17_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_18_clock = clock;
  assign reservation_station_18_reset = reset;
  assign reservation_station_18_io_i_issue_granted = (_issue1_func_code_T_18 | _io_o_issue_packs_1_T_18) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_18_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_18_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_18_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_18_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_18_io_i_write_slot = _reservation_station_18_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_18_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_18_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_18_io_i_uop_valid = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_pc = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_inst = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_func_code = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_target = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_branch_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_select = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_predict_pack_taken = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_phy_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_stale_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_arch_dst = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_inst_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_regWen = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src1_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_phy_rs1 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_arch_rs1 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src2_valid = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_phy_rs2 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_arch_rs2 = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_rob_idx = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_imm = _reservation_station_18_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src1_value = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_src2_value = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_op1_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_op2_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_alu_sel = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_branch_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_uop_mem_type = _reservation_station_18_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_18_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_18_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_18_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_18_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_18_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_19_clock = clock;
  assign reservation_station_19_reset = reset;
  assign reservation_station_19_io_i_issue_granted = (_issue1_func_code_T_19 | _io_o_issue_packs_1_T_19) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_19_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_19_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_19_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_19_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_19_io_i_write_slot = _reservation_station_19_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_19_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_19_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_19_io_i_uop_valid = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_pc = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_inst = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_func_code = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_target = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_branch_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_select = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_predict_pack_taken = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_phy_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_stale_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_arch_dst = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_inst_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_regWen = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src1_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_phy_rs1 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_arch_rs1 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src2_valid = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_phy_rs2 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_arch_rs2 = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_rob_idx = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_imm = _reservation_station_19_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src1_value = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_src2_value = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_op1_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_op2_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_alu_sel = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_branch_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_uop_mem_type = _reservation_station_19_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_19_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_19_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_19_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_19_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_19_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_20_clock = clock;
  assign reservation_station_20_reset = reset;
  assign reservation_station_20_io_i_issue_granted = (_issue1_func_code_T_20 | _io_o_issue_packs_1_T_20) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_20_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_20_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_20_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_20_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_20_io_i_write_slot = _reservation_station_20_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_20_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_20_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_20_io_i_uop_valid = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_pc = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_inst = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_func_code = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_target = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_branch_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_select = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_predict_pack_taken = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_phy_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_stale_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_arch_dst = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_inst_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_regWen = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src1_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_phy_rs1 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_arch_rs1 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src2_valid = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_phy_rs2 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_arch_rs2 = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_rob_idx = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_imm = _reservation_station_20_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src1_value = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_src2_value = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_op1_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_op2_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_alu_sel = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_branch_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_uop_mem_type = _reservation_station_20_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_20_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_20_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_20_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_20_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_20_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_21_clock = clock;
  assign reservation_station_21_reset = reset;
  assign reservation_station_21_io_i_issue_granted = (_issue1_func_code_T_21 | _io_o_issue_packs_1_T_21) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_21_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_21_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_21_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_21_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_21_io_i_write_slot = _reservation_station_21_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_21_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_21_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_21_io_i_uop_valid = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_pc = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_inst = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_func_code = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_target = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_branch_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_select = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_predict_pack_taken = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_phy_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_stale_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_arch_dst = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_inst_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_regWen = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src1_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_phy_rs1 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_arch_rs1 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src2_valid = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_phy_rs2 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_arch_rs2 = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_rob_idx = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_imm = _reservation_station_21_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src1_value = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_src2_value = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_op1_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_op2_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_alu_sel = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_branch_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_uop_mem_type = _reservation_station_21_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_21_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_21_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_21_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_21_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_21_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_22_clock = clock;
  assign reservation_station_22_reset = reset;
  assign reservation_station_22_io_i_issue_granted = (_issue1_func_code_T_22 | _io_o_issue_packs_1_T_22) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_22_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_22_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_22_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_22_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_22_io_i_write_slot = _reservation_station_22_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_22_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_22_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_22_io_i_uop_valid = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_pc = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_inst = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_func_code = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_target = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_branch_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_select = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_predict_pack_taken = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_phy_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_stale_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_arch_dst = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_inst_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_regWen = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src1_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_phy_rs1 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_arch_rs1 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src2_valid = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_phy_rs2 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_arch_rs2 = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_rob_idx = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_imm = _reservation_station_22_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src1_value = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_src2_value = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_op1_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_op2_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_alu_sel = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_branch_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_uop_mem_type = _reservation_station_22_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_22_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_22_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_22_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_22_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_22_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_23_clock = clock;
  assign reservation_station_23_reset = reset;
  assign reservation_station_23_io_i_issue_granted = (_issue1_func_code_T_23 | _io_o_issue_packs_1_T_23) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_23_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_23_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_23_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_23_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_23_io_i_write_slot = _reservation_station_23_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_23_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_23_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_23_io_i_uop_valid = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_pc = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_inst = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_func_code = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_target = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_branch_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_select = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_predict_pack_taken = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_phy_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_stale_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_arch_dst = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_inst_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_regWen = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src1_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_phy_rs1 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_arch_rs1 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src2_valid = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_phy_rs2 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_arch_rs2 = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_rob_idx = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_imm = _reservation_station_23_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src1_value = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_src2_value = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_op1_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_op2_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_alu_sel = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_branch_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_uop_mem_type = _reservation_station_23_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_23_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_23_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_23_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_23_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_23_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_24_clock = clock;
  assign reservation_station_24_reset = reset;
  assign reservation_station_24_io_i_issue_granted = (_issue1_func_code_T_24 | _io_o_issue_packs_1_T_24) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_24_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_24_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_24_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_24_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_24_io_i_write_slot = _reservation_station_24_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_24_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_24_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_24_io_i_uop_valid = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_pc = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_inst = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_func_code = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_target = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_branch_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_select = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_predict_pack_taken = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_phy_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_stale_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_arch_dst = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_inst_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_regWen = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src1_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_phy_rs1 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_arch_rs1 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src2_valid = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_phy_rs2 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_arch_rs2 = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_rob_idx = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_imm = _reservation_station_24_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src1_value = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_src2_value = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_op1_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_op2_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_alu_sel = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_branch_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_uop_mem_type = _reservation_station_24_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_24_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_24_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_24_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_24_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_24_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_25_clock = clock;
  assign reservation_station_25_reset = reset;
  assign reservation_station_25_io_i_issue_granted = (_issue1_func_code_T_25 | _io_o_issue_packs_1_T_25) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_25_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_25_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_25_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_25_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_25_io_i_write_slot = _reservation_station_25_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_25_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_25_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_25_io_i_uop_valid = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_pc = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_inst = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_func_code = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_target = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_branch_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_select = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_predict_pack_taken = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_phy_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_stale_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_arch_dst = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_inst_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_regWen = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src1_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_phy_rs1 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_arch_rs1 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src2_valid = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_phy_rs2 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_arch_rs2 = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_rob_idx = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_imm = _reservation_station_25_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src1_value = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_src2_value = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_op1_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_op2_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_alu_sel = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_branch_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_uop_mem_type = _reservation_station_25_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_25_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_25_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_25_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_25_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_25_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_26_clock = clock;
  assign reservation_station_26_reset = reset;
  assign reservation_station_26_io_i_issue_granted = (_issue1_func_code_T_26 | _io_o_issue_packs_1_T_26) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_26_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_26_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_26_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_26_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_26_io_i_write_slot = _reservation_station_26_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_26_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_26_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_26_io_i_uop_valid = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_pc = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_inst = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_func_code = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_target = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_branch_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_select = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_predict_pack_taken = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_phy_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_stale_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_arch_dst = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_inst_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_regWen = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src1_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_phy_rs1 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_arch_rs1 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src2_valid = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_phy_rs2 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_arch_rs2 = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_rob_idx = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_imm = _reservation_station_26_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src1_value = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_src2_value = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_op1_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_op2_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_alu_sel = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_branch_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_uop_mem_type = _reservation_station_26_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_26_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_26_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_26_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_26_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_26_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_27_clock = clock;
  assign reservation_station_27_reset = reset;
  assign reservation_station_27_io_i_issue_granted = (_issue1_func_code_T_27 | _io_o_issue_packs_1_T_27) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_27_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_27_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_27_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_27_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_27_io_i_write_slot = _reservation_station_27_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_27_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_27_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_27_io_i_uop_valid = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_pc = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_inst = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_func_code = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_target = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_branch_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_select = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_predict_pack_taken = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_phy_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_stale_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_arch_dst = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_inst_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_regWen = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src1_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_phy_rs1 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_arch_rs1 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src2_valid = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_phy_rs2 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_arch_rs2 = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_rob_idx = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_imm = _reservation_station_27_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src1_value = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_src2_value = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_op1_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_op2_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_alu_sel = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_branch_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_uop_mem_type = _reservation_station_27_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_27_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_27_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_27_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_27_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_27_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_28_clock = clock;
  assign reservation_station_28_reset = reset;
  assign reservation_station_28_io_i_issue_granted = (_issue1_func_code_T_28 | _io_o_issue_packs_1_T_28) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_28_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_28_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_28_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_28_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_28_io_i_write_slot = _reservation_station_28_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_28_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_28_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_28_io_i_uop_valid = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_pc = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_inst = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_func_code = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_target = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_branch_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_select = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_predict_pack_taken = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_phy_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_stale_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_arch_dst = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_inst_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_regWen = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src1_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_phy_rs1 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_arch_rs1 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src2_valid = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_phy_rs2 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_arch_rs2 = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_rob_idx = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_imm = _reservation_station_28_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src1_value = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_src2_value = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_op1_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_op2_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_alu_sel = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_branch_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_uop_mem_type = _reservation_station_28_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_28_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_28_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_28_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_28_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_28_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_29_clock = clock;
  assign reservation_station_29_reset = reset;
  assign reservation_station_29_io_i_issue_granted = (_issue1_func_code_T_29 | _io_o_issue_packs_1_T_29) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_29_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_29_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_29_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_29_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_29_io_i_write_slot = _reservation_station_29_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_29_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_29_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_29_io_i_uop_valid = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_pc = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_inst = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_func_code = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_target = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_branch_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_select = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_predict_pack_taken = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_phy_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_stale_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_arch_dst = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_inst_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_regWen = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src1_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_phy_rs1 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_arch_rs1 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src2_valid = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_phy_rs2 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_arch_rs2 = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_rob_idx = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_imm = _reservation_station_29_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src1_value = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_src2_value = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_op1_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_op2_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_alu_sel = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_branch_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_uop_mem_type = _reservation_station_29_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_29_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_29_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_29_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_29_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_29_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_30_clock = clock;
  assign reservation_station_30_reset = reset;
  assign reservation_station_30_io_i_issue_granted = (_issue1_func_code_T_30 | _io_o_issue_packs_1_T_30) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_30_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_30_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_30_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_30_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_30_io_i_write_slot = _reservation_station_30_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_30_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_30_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_30_io_i_uop_valid = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_pc = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_inst = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_func_code = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_target = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_branch_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_select = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_predict_pack_taken = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_phy_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_stale_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_arch_dst = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_inst_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_regWen = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src1_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_phy_rs1 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_arch_rs1 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src2_valid = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_phy_rs2 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_arch_rs2 = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_rob_idx = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_imm = _reservation_station_30_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src1_value = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_src2_value = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_op1_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_op2_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_alu_sel = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_branch_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_uop_mem_type = _reservation_station_30_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_30_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_30_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_30_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_30_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_30_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_31_clock = clock;
  assign reservation_station_31_reset = reset;
  assign reservation_station_31_io_i_issue_granted = (_issue1_func_code_T_31 | _io_o_issue_packs_1_T_31) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_31_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_31_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_31_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_31_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_31_io_i_write_slot = _reservation_station_31_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_31_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_31_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_31_io_i_uop_valid = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_pc = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_inst = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_func_code = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_target = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_branch_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_select = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_predict_pack_taken = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_phy_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_stale_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_arch_dst = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_inst_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_regWen = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src1_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_phy_rs1 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_arch_rs1 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src2_valid = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_phy_rs2 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_arch_rs2 = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_rob_idx = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_imm = _reservation_station_31_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src1_value = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_src2_value = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_op1_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_op2_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_alu_sel = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_branch_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_uop_mem_type = _reservation_station_31_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_31_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_31_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_31_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_31_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_31_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_32_clock = clock;
  assign reservation_station_32_reset = reset;
  assign reservation_station_32_io_i_issue_granted = (_issue1_func_code_T_32 | _io_o_issue_packs_1_T_32) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_32_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_32_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_32_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_32_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_32_io_i_write_slot = _reservation_station_32_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_32_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_32_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_32_io_i_uop_valid = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_pc = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_inst = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_func_code = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_valid = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_target = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_branch_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_select = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_branch_predict_pack_taken = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_phy_dst = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_stale_dst = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_arch_dst = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_inst_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_regWen = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_src1_valid = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_phy_rs1 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_arch_rs1 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_src2_valid = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_phy_rs2 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_arch_rs2 = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_rob_idx = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_imm = _reservation_station_32_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_src1_value = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_src2_value = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_op1_sel = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_op2_sel = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_alu_sel = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_branch_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_uop_mem_type = _reservation_station_32_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_32_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_32_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_32_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_32_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_32_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_33_clock = clock;
  assign reservation_station_33_reset = reset;
  assign reservation_station_33_io_i_issue_granted = (_issue1_func_code_T_33 | _io_o_issue_packs_1_T_33) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_33_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_33_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_33_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_33_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_33_io_i_write_slot = _reservation_station_33_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_33_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_33_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_33_io_i_uop_valid = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_pc = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_inst = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_func_code = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_valid = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_target = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_branch_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_select = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_branch_predict_pack_taken = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_phy_dst = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_stale_dst = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_arch_dst = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_inst_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_regWen = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_src1_valid = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_phy_rs1 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_arch_rs1 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_src2_valid = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_phy_rs2 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_arch_rs2 = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_rob_idx = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_imm = _reservation_station_33_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_src1_value = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_src2_value = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_op1_sel = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_op2_sel = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_alu_sel = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_branch_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_uop_mem_type = _reservation_station_33_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_33_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_33_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_33_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_33_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_33_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_34_clock = clock;
  assign reservation_station_34_reset = reset;
  assign reservation_station_34_io_i_issue_granted = (_issue1_func_code_T_34 | _io_o_issue_packs_1_T_34) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_34_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_34_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_34_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_34_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_34_io_i_write_slot = _reservation_station_34_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_34_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_34_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_34_io_i_uop_valid = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_pc = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_inst = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_func_code = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_valid = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_target = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_branch_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_select = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_branch_predict_pack_taken = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_phy_dst = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_stale_dst = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_arch_dst = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_inst_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_regWen = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_src1_valid = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_phy_rs1 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_arch_rs1 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_src2_valid = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_phy_rs2 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_arch_rs2 = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_rob_idx = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_imm = _reservation_station_34_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_src1_value = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_src2_value = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_op1_sel = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_op2_sel = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_alu_sel = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_branch_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_uop_mem_type = _reservation_station_34_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_34_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_34_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_34_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_34_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_34_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_35_clock = clock;
  assign reservation_station_35_reset = reset;
  assign reservation_station_35_io_i_issue_granted = (_issue1_func_code_T_35 | _io_o_issue_packs_1_T_35) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_35_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_35_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_35_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_35_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_35_io_i_write_slot = _reservation_station_35_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_35_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_35_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_35_io_i_uop_valid = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_pc = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_inst = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_func_code = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_valid = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_target = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_branch_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_select = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_branch_predict_pack_taken = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_phy_dst = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_stale_dst = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_arch_dst = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_inst_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_regWen = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_src1_valid = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_phy_rs1 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_arch_rs1 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_src2_valid = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_phy_rs2 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_arch_rs2 = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_rob_idx = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_imm = _reservation_station_35_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_src1_value = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_src2_value = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_op1_sel = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_op2_sel = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_alu_sel = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_branch_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_uop_mem_type = _reservation_station_35_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_35_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_35_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_35_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_35_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_35_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_36_clock = clock;
  assign reservation_station_36_reset = reset;
  assign reservation_station_36_io_i_issue_granted = (_issue1_func_code_T_36 | _io_o_issue_packs_1_T_36) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_36_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_36_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_36_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_36_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_36_io_i_write_slot = _reservation_station_36_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_36_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_36_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_36_io_i_uop_valid = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_pc = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_inst = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_func_code = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_valid = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_target = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_branch_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_select = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_branch_predict_pack_taken = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_phy_dst = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_stale_dst = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_arch_dst = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_inst_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_regWen = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_src1_valid = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_phy_rs1 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_arch_rs1 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_src2_valid = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_phy_rs2 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_arch_rs2 = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_rob_idx = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_imm = _reservation_station_36_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_src1_value = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_src2_value = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_op1_sel = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_op2_sel = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_alu_sel = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_branch_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_uop_mem_type = _reservation_station_36_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_36_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_36_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_36_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_36_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_36_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_37_clock = clock;
  assign reservation_station_37_reset = reset;
  assign reservation_station_37_io_i_issue_granted = (_issue1_func_code_T_37 | _io_o_issue_packs_1_T_37) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_37_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_37_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_37_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_37_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_37_io_i_write_slot = _reservation_station_37_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_37_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_37_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_37_io_i_uop_valid = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_pc = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_inst = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_func_code = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_valid = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_target = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_branch_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_select = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_branch_predict_pack_taken = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_phy_dst = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_stale_dst = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_arch_dst = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_inst_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_regWen = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_src1_valid = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_phy_rs1 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_arch_rs1 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_src2_valid = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_phy_rs2 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_arch_rs2 = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_rob_idx = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_imm = _reservation_station_37_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_src1_value = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_src2_value = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_op1_sel = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_op2_sel = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_alu_sel = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_branch_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_uop_mem_type = _reservation_station_37_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_37_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_37_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_37_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_37_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_37_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_38_clock = clock;
  assign reservation_station_38_reset = reset;
  assign reservation_station_38_io_i_issue_granted = (_issue1_func_code_T_38 | _io_o_issue_packs_1_T_38) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_38_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_38_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_38_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_38_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_38_io_i_write_slot = _reservation_station_38_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_38_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_38_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_38_io_i_uop_valid = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_pc = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_inst = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_func_code = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_valid = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_target = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_branch_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_select = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_branch_predict_pack_taken = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_phy_dst = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_stale_dst = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_arch_dst = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_inst_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_regWen = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_src1_valid = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_phy_rs1 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_arch_rs1 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_src2_valid = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_phy_rs2 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_arch_rs2 = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_rob_idx = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_imm = _reservation_station_38_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_src1_value = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_src2_value = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_op1_sel = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_op2_sel = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_alu_sel = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_branch_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_uop_mem_type = _reservation_station_38_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_38_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_38_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_38_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_38_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_38_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_39_clock = clock;
  assign reservation_station_39_reset = reset;
  assign reservation_station_39_io_i_issue_granted = (_issue1_func_code_T_39 | _io_o_issue_packs_1_T_39) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_39_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_39_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_39_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_39_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_39_io_i_write_slot = _reservation_station_39_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_39_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_39_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_39_io_i_uop_valid = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_pc = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_inst = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_func_code = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_valid = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_target = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_branch_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_select = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_branch_predict_pack_taken = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_phy_dst = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_stale_dst = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_arch_dst = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_inst_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_regWen = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_src1_valid = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_phy_rs1 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_arch_rs1 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_src2_valid = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_phy_rs2 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_arch_rs2 = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_rob_idx = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_imm = _reservation_station_39_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_src1_value = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_src2_value = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_op1_sel = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_op2_sel = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_alu_sel = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_branch_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_uop_mem_type = _reservation_station_39_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_39_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_39_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_39_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_39_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_39_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_40_clock = clock;
  assign reservation_station_40_reset = reset;
  assign reservation_station_40_io_i_issue_granted = (_issue1_func_code_T_40 | _io_o_issue_packs_1_T_40) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_40_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_40_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_40_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_40_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_40_io_i_write_slot = _reservation_station_40_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_40_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_40_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_40_io_i_uop_valid = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_pc = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_inst = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_func_code = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_valid = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_target = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_branch_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_select = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_branch_predict_pack_taken = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_phy_dst = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_stale_dst = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_arch_dst = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_inst_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_regWen = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_src1_valid = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_phy_rs1 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_arch_rs1 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_src2_valid = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_phy_rs2 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_arch_rs2 = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_rob_idx = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_imm = _reservation_station_40_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_src1_value = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_src2_value = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_op1_sel = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_op2_sel = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_alu_sel = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_branch_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_uop_mem_type = _reservation_station_40_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_40_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_40_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_40_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_40_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_40_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_41_clock = clock;
  assign reservation_station_41_reset = reset;
  assign reservation_station_41_io_i_issue_granted = (_issue1_func_code_T_41 | _io_o_issue_packs_1_T_41) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_41_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_41_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_41_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_41_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_41_io_i_write_slot = _reservation_station_41_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_41_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_41_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_41_io_i_uop_valid = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_pc = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_inst = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_func_code = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_valid = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_target = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_branch_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_select = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_branch_predict_pack_taken = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_phy_dst = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_stale_dst = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_arch_dst = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_inst_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_regWen = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_src1_valid = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_phy_rs1 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_arch_rs1 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_src2_valid = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_phy_rs2 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_arch_rs2 = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_rob_idx = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_imm = _reservation_station_41_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_src1_value = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_src2_value = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_op1_sel = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_op2_sel = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_alu_sel = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_branch_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_uop_mem_type = _reservation_station_41_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_41_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_41_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_41_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_41_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_41_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_42_clock = clock;
  assign reservation_station_42_reset = reset;
  assign reservation_station_42_io_i_issue_granted = (_issue1_func_code_T_42 | _io_o_issue_packs_1_T_42) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_42_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_42_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_42_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_42_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_42_io_i_write_slot = _reservation_station_42_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_42_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_42_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_42_io_i_uop_valid = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_pc = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_inst = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_func_code = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_valid = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_target = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_branch_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_select = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_branch_predict_pack_taken = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_phy_dst = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_stale_dst = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_arch_dst = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_inst_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_regWen = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_src1_valid = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_phy_rs1 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_arch_rs1 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_src2_valid = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_phy_rs2 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_arch_rs2 = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_rob_idx = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_imm = _reservation_station_42_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_src1_value = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_src2_value = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_op1_sel = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_op2_sel = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_alu_sel = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_branch_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_uop_mem_type = _reservation_station_42_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_42_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_42_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_42_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_42_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_42_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_43_clock = clock;
  assign reservation_station_43_reset = reset;
  assign reservation_station_43_io_i_issue_granted = (_issue1_func_code_T_43 | _io_o_issue_packs_1_T_43) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_43_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_43_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_43_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_43_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_43_io_i_write_slot = _reservation_station_43_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_43_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_43_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_43_io_i_uop_valid = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_pc = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_inst = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_func_code = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_valid = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_target = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_branch_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_select = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_branch_predict_pack_taken = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_phy_dst = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_stale_dst = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_arch_dst = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_inst_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_regWen = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_src1_valid = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_phy_rs1 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_arch_rs1 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_src2_valid = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_phy_rs2 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_arch_rs2 = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_rob_idx = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_imm = _reservation_station_43_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_src1_value = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_src2_value = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_op1_sel = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_op2_sel = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_alu_sel = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_branch_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_uop_mem_type = _reservation_station_43_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_43_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_43_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_43_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_43_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_43_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_44_clock = clock;
  assign reservation_station_44_reset = reset;
  assign reservation_station_44_io_i_issue_granted = (_issue1_func_code_T_44 | _io_o_issue_packs_1_T_44) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_44_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_44_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_44_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_44_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_44_io_i_write_slot = _reservation_station_44_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_44_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_44_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_44_io_i_uop_valid = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_pc = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_inst = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_func_code = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_valid = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_target = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_branch_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_select = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_branch_predict_pack_taken = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_phy_dst = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_stale_dst = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_arch_dst = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_inst_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_regWen = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_src1_valid = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_phy_rs1 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_arch_rs1 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_src2_valid = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_phy_rs2 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_arch_rs2 = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_rob_idx = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_imm = _reservation_station_44_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_src1_value = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_src2_value = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_op1_sel = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_op2_sel = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_alu_sel = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_branch_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_uop_mem_type = _reservation_station_44_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_44_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_44_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_44_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_44_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_44_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_45_clock = clock;
  assign reservation_station_45_reset = reset;
  assign reservation_station_45_io_i_issue_granted = (_issue1_func_code_T_45 | _io_o_issue_packs_1_T_45) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_45_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_45_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_45_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_45_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_45_io_i_write_slot = _reservation_station_45_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_45_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_45_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_45_io_i_uop_valid = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_pc = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_inst = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_func_code = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_valid = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_target = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_branch_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_select = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_branch_predict_pack_taken = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_phy_dst = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_stale_dst = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_arch_dst = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_inst_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_regWen = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_src1_valid = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_phy_rs1 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_arch_rs1 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_src2_valid = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_phy_rs2 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_arch_rs2 = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_rob_idx = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_imm = _reservation_station_45_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_src1_value = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_src2_value = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_op1_sel = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_op2_sel = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_alu_sel = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_branch_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_uop_mem_type = _reservation_station_45_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_45_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_45_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_45_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_45_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_45_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_46_clock = clock;
  assign reservation_station_46_reset = reset;
  assign reservation_station_46_io_i_issue_granted = (_issue1_func_code_T_46 | _io_o_issue_packs_1_T_46) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_46_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_46_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_46_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_46_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_46_io_i_write_slot = _reservation_station_46_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_46_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_46_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_46_io_i_uop_valid = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_pc = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_inst = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_func_code = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_valid = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_target = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_branch_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_select = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_branch_predict_pack_taken = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_phy_dst = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_stale_dst = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_arch_dst = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_inst_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_regWen = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_src1_valid = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_phy_rs1 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_arch_rs1 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_src2_valid = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_phy_rs2 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_arch_rs2 = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_rob_idx = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_imm = _reservation_station_46_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_src1_value = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_src2_value = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_op1_sel = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_op2_sel = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_alu_sel = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_branch_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_uop_mem_type = _reservation_station_46_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_46_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_46_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_46_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_46_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_46_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_47_clock = clock;
  assign reservation_station_47_reset = reset;
  assign reservation_station_47_io_i_issue_granted = (_issue1_func_code_T_47 | _io_o_issue_packs_1_T_47) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_47_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_47_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_47_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_47_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_47_io_i_write_slot = _reservation_station_47_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_47_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_47_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_47_io_i_uop_valid = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_pc = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_inst = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_func_code = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_valid = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_target = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_branch_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_select = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_branch_predict_pack_taken = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_phy_dst = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_stale_dst = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_arch_dst = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_inst_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_regWen = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_src1_valid = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_phy_rs1 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_arch_rs1 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_src2_valid = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_phy_rs2 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_arch_rs2 = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_rob_idx = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_imm = _reservation_station_47_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_src1_value = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_src2_value = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_op1_sel = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_op2_sel = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_alu_sel = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_branch_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_uop_mem_type = _reservation_station_47_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_47_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_47_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_47_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_47_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_47_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_48_clock = clock;
  assign reservation_station_48_reset = reset;
  assign reservation_station_48_io_i_issue_granted = (_issue1_func_code_T_48 | _io_o_issue_packs_1_T_48) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_48_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_48_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_48_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_48_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_48_io_i_write_slot = _reservation_station_48_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_48_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_48_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_48_io_i_uop_valid = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_pc = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_inst = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_func_code = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_valid = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_target = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_branch_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_select = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_branch_predict_pack_taken = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_phy_dst = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_stale_dst = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_arch_dst = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_inst_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_regWen = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_src1_valid = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_phy_rs1 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_arch_rs1 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_src2_valid = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_phy_rs2 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_arch_rs2 = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_rob_idx = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_imm = _reservation_station_48_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_src1_value = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_src2_value = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_op1_sel = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_op2_sel = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_alu_sel = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_branch_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_uop_mem_type = _reservation_station_48_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_48_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_48_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_48_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_48_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_48_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_49_clock = clock;
  assign reservation_station_49_reset = reset;
  assign reservation_station_49_io_i_issue_granted = (_issue1_func_code_T_49 | _io_o_issue_packs_1_T_49) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_49_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_49_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_49_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_49_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_49_io_i_write_slot = _reservation_station_49_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_49_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_49_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_49_io_i_uop_valid = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_pc = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_inst = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_func_code = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_valid = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_target = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_branch_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_select = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_branch_predict_pack_taken = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_phy_dst = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_stale_dst = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_arch_dst = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_inst_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_regWen = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_src1_valid = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_phy_rs1 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_arch_rs1 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_src2_valid = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_phy_rs2 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_arch_rs2 = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_rob_idx = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_imm = _reservation_station_49_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_src1_value = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_src2_value = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_op1_sel = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_op2_sel = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_alu_sel = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_branch_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_uop_mem_type = _reservation_station_49_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_49_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_49_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_49_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_49_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_49_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_50_clock = clock;
  assign reservation_station_50_reset = reset;
  assign reservation_station_50_io_i_issue_granted = (_issue1_func_code_T_50 | _io_o_issue_packs_1_T_50) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_50_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_50_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_50_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_50_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_50_io_i_write_slot = _reservation_station_50_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_50_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_50_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_50_io_i_uop_valid = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_pc = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_inst = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_func_code = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_valid = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_target = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_branch_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_select = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_branch_predict_pack_taken = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_phy_dst = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_stale_dst = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_arch_dst = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_inst_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_regWen = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_src1_valid = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_phy_rs1 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_arch_rs1 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_src2_valid = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_phy_rs2 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_arch_rs2 = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_rob_idx = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_imm = _reservation_station_50_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_src1_value = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_src2_value = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_op1_sel = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_op2_sel = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_alu_sel = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_branch_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_uop_mem_type = _reservation_station_50_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_50_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_50_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_50_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_50_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_50_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_51_clock = clock;
  assign reservation_station_51_reset = reset;
  assign reservation_station_51_io_i_issue_granted = (_issue1_func_code_T_51 | _io_o_issue_packs_1_T_51) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_51_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_51_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_51_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_51_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_51_io_i_write_slot = _reservation_station_51_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_51_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_51_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_51_io_i_uop_valid = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_pc = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_inst = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_func_code = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_valid = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_target = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_branch_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_select = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_branch_predict_pack_taken = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_phy_dst = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_stale_dst = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_arch_dst = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_inst_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_regWen = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_src1_valid = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_phy_rs1 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_arch_rs1 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_src2_valid = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_phy_rs2 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_arch_rs2 = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_rob_idx = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_imm = _reservation_station_51_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_src1_value = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_src2_value = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_op1_sel = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_op2_sel = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_alu_sel = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_branch_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_uop_mem_type = _reservation_station_51_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_51_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_51_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_51_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_51_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_51_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_52_clock = clock;
  assign reservation_station_52_reset = reset;
  assign reservation_station_52_io_i_issue_granted = (_issue1_func_code_T_52 | _io_o_issue_packs_1_T_52) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_52_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_52_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_52_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_52_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_52_io_i_write_slot = _reservation_station_52_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_52_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_52_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_52_io_i_uop_valid = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_pc = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_inst = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_func_code = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_valid = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_target = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_branch_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_select = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_branch_predict_pack_taken = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_phy_dst = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_stale_dst = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_arch_dst = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_inst_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_regWen = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_src1_valid = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_phy_rs1 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_arch_rs1 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_src2_valid = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_phy_rs2 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_arch_rs2 = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_rob_idx = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_imm = _reservation_station_52_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_src1_value = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_src2_value = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_op1_sel = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_op2_sel = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_alu_sel = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_branch_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_uop_mem_type = _reservation_station_52_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_52_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_52_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_52_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_52_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_52_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_53_clock = clock;
  assign reservation_station_53_reset = reset;
  assign reservation_station_53_io_i_issue_granted = (_issue1_func_code_T_53 | _io_o_issue_packs_1_T_53) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_53_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_53_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_53_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_53_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_53_io_i_write_slot = _reservation_station_53_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_53_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_53_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_53_io_i_uop_valid = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_pc = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_inst = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_func_code = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_valid = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_target = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_branch_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_select = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_branch_predict_pack_taken = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_phy_dst = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_stale_dst = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_arch_dst = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_inst_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_regWen = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_src1_valid = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_phy_rs1 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_arch_rs1 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_src2_valid = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_phy_rs2 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_arch_rs2 = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_rob_idx = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_imm = _reservation_station_53_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_src1_value = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_src2_value = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_op1_sel = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_op2_sel = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_alu_sel = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_branch_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_uop_mem_type = _reservation_station_53_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_53_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_53_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_53_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_53_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_53_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_54_clock = clock;
  assign reservation_station_54_reset = reset;
  assign reservation_station_54_io_i_issue_granted = (_issue1_func_code_T_54 | _io_o_issue_packs_1_T_54) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_54_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_54_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_54_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_54_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_54_io_i_write_slot = _reservation_station_54_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_54_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_54_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_54_io_i_uop_valid = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_pc = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_inst = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_func_code = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_valid = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_target = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_branch_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_select = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_branch_predict_pack_taken = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_phy_dst = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_stale_dst = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_arch_dst = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_inst_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_regWen = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_src1_valid = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_phy_rs1 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_arch_rs1 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_src2_valid = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_phy_rs2 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_arch_rs2 = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_rob_idx = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_imm = _reservation_station_54_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_src1_value = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_src2_value = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_op1_sel = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_op2_sel = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_alu_sel = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_branch_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_uop_mem_type = _reservation_station_54_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_54_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_54_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_54_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_54_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_54_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_55_clock = clock;
  assign reservation_station_55_reset = reset;
  assign reservation_station_55_io_i_issue_granted = (_issue1_func_code_T_55 | _io_o_issue_packs_1_T_55) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_55_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_55_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_55_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_55_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_55_io_i_write_slot = _reservation_station_55_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_55_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_55_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_55_io_i_uop_valid = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_pc = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_inst = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_func_code = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_valid = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_target = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_branch_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_select = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_branch_predict_pack_taken = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_phy_dst = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_stale_dst = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_arch_dst = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_inst_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_regWen = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_src1_valid = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_phy_rs1 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_arch_rs1 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_src2_valid = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_phy_rs2 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_arch_rs2 = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_rob_idx = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_imm = _reservation_station_55_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_src1_value = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_src2_value = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_op1_sel = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_op2_sel = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_alu_sel = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_branch_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_uop_mem_type = _reservation_station_55_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_55_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_55_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_55_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_55_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_55_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_56_clock = clock;
  assign reservation_station_56_reset = reset;
  assign reservation_station_56_io_i_issue_granted = (_issue1_func_code_T_56 | _io_o_issue_packs_1_T_56) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_56_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_56_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_56_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_56_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_56_io_i_write_slot = _reservation_station_56_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_56_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_56_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_56_io_i_uop_valid = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_pc = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_inst = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_func_code = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_valid = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_target = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_branch_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_select = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_branch_predict_pack_taken = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_phy_dst = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_stale_dst = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_arch_dst = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_inst_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_regWen = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_src1_valid = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_phy_rs1 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_arch_rs1 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_src2_valid = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_phy_rs2 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_arch_rs2 = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_rob_idx = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_imm = _reservation_station_56_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_src1_value = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_src2_value = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_op1_sel = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_op2_sel = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_alu_sel = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_branch_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_uop_mem_type = _reservation_station_56_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_56_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_56_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_56_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_56_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_56_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_57_clock = clock;
  assign reservation_station_57_reset = reset;
  assign reservation_station_57_io_i_issue_granted = (_issue1_func_code_T_57 | _io_o_issue_packs_1_T_57) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_57_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_57_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_57_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_57_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_57_io_i_write_slot = _reservation_station_57_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_57_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_57_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_57_io_i_uop_valid = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_pc = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_inst = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_func_code = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_valid = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_target = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_branch_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_select = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_branch_predict_pack_taken = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_phy_dst = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_stale_dst = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_arch_dst = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_inst_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_regWen = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_src1_valid = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_phy_rs1 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_arch_rs1 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_src2_valid = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_phy_rs2 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_arch_rs2 = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_rob_idx = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_imm = _reservation_station_57_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_src1_value = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_src2_value = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_op1_sel = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_op2_sel = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_alu_sel = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_branch_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_uop_mem_type = _reservation_station_57_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_57_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_57_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_57_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_57_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_57_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_58_clock = clock;
  assign reservation_station_58_reset = reset;
  assign reservation_station_58_io_i_issue_granted = (_issue1_func_code_T_58 | _io_o_issue_packs_1_T_58) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_58_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_58_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_58_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_58_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_58_io_i_write_slot = _reservation_station_58_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_58_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_58_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_58_io_i_uop_valid = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_pc = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_inst = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_func_code = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_valid = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_target = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_branch_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_select = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_branch_predict_pack_taken = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_phy_dst = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_stale_dst = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_arch_dst = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_inst_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_regWen = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_src1_valid = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_phy_rs1 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_arch_rs1 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_src2_valid = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_phy_rs2 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_arch_rs2 = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_rob_idx = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_imm = _reservation_station_58_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_src1_value = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_src2_value = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_op1_sel = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_op2_sel = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_alu_sel = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_branch_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_uop_mem_type = _reservation_station_58_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_58_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_58_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_58_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_58_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_58_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_59_clock = clock;
  assign reservation_station_59_reset = reset;
  assign reservation_station_59_io_i_issue_granted = (_issue1_func_code_T_59 | _io_o_issue_packs_1_T_59) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_59_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_59_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_59_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_59_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_59_io_i_write_slot = _reservation_station_59_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_59_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_59_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_59_io_i_uop_valid = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_pc = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_inst = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_func_code = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_valid = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_target = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_branch_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_select = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_branch_predict_pack_taken = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_phy_dst = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_stale_dst = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_arch_dst = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_inst_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_regWen = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_src1_valid = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_phy_rs1 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_arch_rs1 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_src2_valid = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_phy_rs2 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_arch_rs2 = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_rob_idx = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_imm = _reservation_station_59_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_src1_value = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_src2_value = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_op1_sel = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_op2_sel = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_alu_sel = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_branch_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_uop_mem_type = _reservation_station_59_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_59_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_59_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_59_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_59_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_59_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_60_clock = clock;
  assign reservation_station_60_reset = reset;
  assign reservation_station_60_io_i_issue_granted = (_issue1_func_code_T_60 | _io_o_issue_packs_1_T_60) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_60_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_60_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_60_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_60_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_60_io_i_write_slot = _reservation_station_60_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_60_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_60_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_60_io_i_uop_valid = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_pc = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_inst = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_func_code = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_valid = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_target = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_branch_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_select = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_branch_predict_pack_taken = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_phy_dst = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_stale_dst = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_arch_dst = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_inst_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_regWen = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_src1_valid = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_phy_rs1 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_arch_rs1 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_src2_valid = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_phy_rs2 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_arch_rs2 = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_rob_idx = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_imm = _reservation_station_60_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_src1_value = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_src2_value = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_op1_sel = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_op2_sel = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_alu_sel = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_branch_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_uop_mem_type = _reservation_station_60_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_60_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_60_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_60_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_60_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_60_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_61_clock = clock;
  assign reservation_station_61_reset = reset;
  assign reservation_station_61_io_i_issue_granted = (_issue1_func_code_T_61 | _io_o_issue_packs_1_T_61) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_61_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_61_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_61_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_61_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_61_io_i_write_slot = _reservation_station_61_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_61_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_61_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_61_io_i_uop_valid = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_pc = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_inst = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_func_code = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_valid = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_target = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_branch_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_select = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_branch_predict_pack_taken = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_phy_dst = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_stale_dst = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_arch_dst = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_inst_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_regWen = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_src1_valid = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_phy_rs1 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_arch_rs1 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_src2_valid = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_phy_rs2 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_arch_rs2 = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_rob_idx = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_imm = _reservation_station_61_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_src1_value = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_src2_value = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_op1_sel = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_op2_sel = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_alu_sel = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_branch_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_uop_mem_type = _reservation_station_61_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_61_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_61_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_61_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_61_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_61_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_62_clock = clock;
  assign reservation_station_62_reset = reset;
  assign reservation_station_62_io_i_issue_granted = (_issue1_func_code_T_62 | _io_o_issue_packs_1_T_62) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_62_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_62_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_62_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_62_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_62_io_i_write_slot = _reservation_station_62_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_62_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_62_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_62_io_i_uop_valid = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_pc = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_inst = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_func_code = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_valid = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_target = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_branch_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_select = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_branch_predict_pack_taken = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_phy_dst = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_stale_dst = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_arch_dst = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_inst_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_regWen = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_src1_valid = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_phy_rs1 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_arch_rs1 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_src2_valid = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_phy_rs2 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_arch_rs2 = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_rob_idx = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_imm = _reservation_station_62_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_src1_value = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_src2_value = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_op1_sel = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_op2_sel = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_alu_sel = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_branch_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_uop_mem_type = _reservation_station_62_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_62_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_62_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_62_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_62_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_62_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
  assign reservation_station_63_clock = clock;
  assign reservation_station_63_reset = reset;
  assign reservation_station_63_io_i_issue_granted = (_issue1_func_code_T_63 | _io_o_issue_packs_1_T_63) & ~(
    io_i_exception | io_i_rollback_valid); // @[reservation_station.scala 112:94]
  assign reservation_station_63_io_i_branch_resolve_pack_valid = io_i_branch_resolve_pack_valid; // @[reservation_station.scala 113:54]
  assign reservation_station_63_io_i_branch_resolve_pack_mispred = io_i_branch_resolve_pack_mispred; // @[reservation_station.scala 113:54]
  assign reservation_station_63_io_i_branch_resolve_pack_rob_idx = io_i_branch_resolve_pack_rob_idx; // @[reservation_station.scala 113:54]
  assign reservation_station_63_io_i_exception = io_i_exception; // @[reservation_station.scala 114:44]
  assign reservation_station_63_io_i_write_slot = _reservation_station_63_io_i_write_slot_T_2 ?
    io_i_dispatch_packs_0_valid : _reservation_station_63_io_i_write_slot_T_5 & io_i_dispatch_packs_1_valid; // @[Mux.scala 101:16]
  assign reservation_station_63_io_i_wakeup_port = io_i_wakeup_port; // @[reservation_station.scala 115:46]
  assign reservation_station_63_io_i_uop_valid = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_valid
     : io_i_dispatch_packs_1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_pc = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_pc :
    io_i_dispatch_packs_1_pc; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_inst = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_inst
     : io_i_dispatch_packs_1_inst; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_func_code = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_func_code : io_i_dispatch_packs_1_func_code; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_valid = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_valid : io_i_dispatch_packs_1_branch_predict_pack_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_target = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_target : io_i_dispatch_packs_1_branch_predict_pack_target; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_branch_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_branch_type : io_i_dispatch_packs_1_branch_predict_pack_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_select = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_select : io_i_dispatch_packs_1_branch_predict_pack_select; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_branch_predict_pack_taken = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_predict_pack_taken : io_i_dispatch_packs_1_branch_predict_pack_taken; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_phy_dst = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_dst : io_i_dispatch_packs_1_phy_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_stale_dst = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_stale_dst : io_i_dispatch_packs_1_stale_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_arch_dst = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_dst : io_i_dispatch_packs_1_arch_dst; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_inst_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_inst_type : io_i_dispatch_packs_1_inst_type; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_regWen = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_regWen : io_i_dispatch_packs_1_regWen; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_src1_valid = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_valid : io_i_dispatch_packs_1_src1_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_phy_rs1 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs1 : io_i_dispatch_packs_1_phy_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_arch_rs1 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs1 : io_i_dispatch_packs_1_arch_rs1; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_src2_valid = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_valid : io_i_dispatch_packs_1_src2_valid; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_phy_rs2 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_phy_rs2 : io_i_dispatch_packs_1_phy_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_arch_rs2 = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_arch_rs2 : io_i_dispatch_packs_1_arch_rs2; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_rob_idx = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_rob_idx : io_i_dispatch_packs_1_rob_idx; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_imm = _reservation_station_63_io_i_write_slot_T ? io_i_dispatch_packs_0_imm :
    io_i_dispatch_packs_1_imm; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_src1_value = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src1_value : io_i_dispatch_packs_1_src1_value; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_src2_value = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_src2_value : io_i_dispatch_packs_1_src2_value; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_op1_sel = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op1_sel : io_i_dispatch_packs_1_op1_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_op2_sel = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_op2_sel : io_i_dispatch_packs_1_op2_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_alu_sel = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_alu_sel : io_i_dispatch_packs_1_alu_sel; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_branch_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_branch_type : io_i_dispatch_packs_1_branch_type; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_uop_mem_type = _reservation_station_63_io_i_write_slot_T ?
    io_i_dispatch_packs_0_mem_type : io_i_dispatch_packs_1_mem_type; // @[reservation_station.scala 123:44]
  assign reservation_station_63_io_i_exe_dst1 = io_i_ex_res_packs_0_valid & io_i_ex_res_packs_0_uop_func_code != 7'h20
     ? io_i_ex_res_packs_0_uop_phy_dst : 7'h0; // @[reservation_station.scala 126:49]
  assign reservation_station_63_io_i_exe_dst2 = io_i_ex_res_packs_1_valid & io_i_ex_res_packs_1_uop_func_code != 7'h20
     ? io_i_ex_res_packs_1_uop_phy_dst : 7'h0; // @[reservation_station.scala 127:49]
  assign reservation_station_63_io_i_exe_value1 = io_i_ex_res_packs_0_uop_dst_value; // @[reservation_station.scala 129:45]
  assign reservation_station_63_io_i_exe_value2 = io_i_ex_res_packs_1_uop_dst_value; // @[reservation_station.scala 130:45]
  assign reservation_station_63_io_i_ROB_first_entry = io_i_ROB_first_entry; // @[reservation_station.scala 132:50]
endmodule

module Wallace_Tree(
  input  [130:0] io_i_partial_products_0,
  input  [130:0] io_i_partial_products_1,
  input  [130:0] io_i_partial_products_2,
  input  [130:0] io_i_partial_products_3,
  input  [130:0] io_i_partial_products_4,
  input  [130:0] io_i_partial_products_5,
  input  [130:0] io_i_partial_products_6,
  input  [130:0] io_i_partial_products_7,
  input  [130:0] io_i_partial_products_8,
  input  [130:0] io_i_partial_products_9,
  input  [130:0] io_i_partial_products_10,
  input  [130:0] io_i_partial_products_11,
  input  [130:0] io_i_partial_products_12,
  input  [130:0] io_i_partial_products_13,
  input  [130:0] io_i_partial_products_14,
  input  [130:0] io_i_partial_products_15,
  input  [130:0] io_i_partial_products_16,
  input  [130:0] io_i_partial_products_17,
  input  [130:0] io_i_partial_products_18,
  input  [130:0] io_i_partial_products_19,
  input  [130:0] io_i_partial_products_20,
  input  [130:0] io_i_partial_products_21,
  output [130:0] io_o_s,
  output [130:0] io_o_c
);
  wire [18:0] wallace_tree_cells_0_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_0_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_0_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_0_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_0_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_1_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_1_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_1_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_1_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_1_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_2_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_2_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_2_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_2_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_2_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_3_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_3_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_3_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_3_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_3_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_4_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_4_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_4_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_4_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_4_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_5_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_5_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_5_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_5_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_5_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_6_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_6_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_6_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_6_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_6_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_7_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_7_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_7_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_7_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_7_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_8_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_8_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_8_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_8_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_8_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_9_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_9_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_9_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_9_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_9_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_10_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_10_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_10_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_10_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_10_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_11_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_11_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_11_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_11_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_11_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_12_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_12_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_12_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_12_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_12_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_13_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_13_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_13_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_13_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_13_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_14_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_14_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_14_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_14_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_14_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_15_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_15_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_15_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_15_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_15_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_16_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_16_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_16_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_16_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_16_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_17_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_17_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_17_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_17_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_17_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_18_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_18_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_18_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_18_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_18_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_19_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_19_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_19_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_19_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_19_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_20_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_20_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_20_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_20_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_20_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_21_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_21_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_21_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_21_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_21_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_22_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_22_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_22_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_22_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_22_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_23_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_23_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_23_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_23_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_23_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_24_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_24_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_24_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_24_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_24_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_25_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_25_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_25_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_25_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_25_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_26_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_26_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_26_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_26_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_26_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_27_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_27_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_27_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_27_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_27_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_28_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_28_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_28_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_28_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_28_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_29_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_29_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_29_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_29_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_29_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_30_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_30_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_30_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_30_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_30_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_31_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_31_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_31_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_31_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_31_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_32_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_32_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_32_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_32_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_32_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_33_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_33_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_33_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_33_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_33_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_34_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_34_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_34_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_34_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_34_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_35_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_35_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_35_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_35_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_35_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_36_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_36_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_36_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_36_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_36_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_37_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_37_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_37_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_37_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_37_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_38_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_38_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_38_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_38_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_38_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_39_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_39_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_39_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_39_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_39_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_40_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_40_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_40_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_40_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_40_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_41_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_41_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_41_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_41_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_41_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_42_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_42_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_42_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_42_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_42_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_43_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_43_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_43_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_43_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_43_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_44_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_44_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_44_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_44_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_44_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_45_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_45_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_45_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_45_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_45_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_46_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_46_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_46_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_46_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_46_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_47_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_47_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_47_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_47_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_47_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_48_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_48_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_48_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_48_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_48_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_49_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_49_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_49_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_49_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_49_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_50_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_50_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_50_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_50_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_50_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_51_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_51_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_51_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_51_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_51_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_52_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_52_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_52_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_52_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_52_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_53_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_53_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_53_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_53_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_53_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_54_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_54_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_54_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_54_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_54_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_55_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_55_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_55_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_55_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_55_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_56_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_56_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_56_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_56_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_56_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_57_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_57_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_57_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_57_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_57_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_58_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_58_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_58_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_58_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_58_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_59_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_59_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_59_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_59_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_59_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_60_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_60_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_60_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_60_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_60_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_61_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_61_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_61_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_61_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_61_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_62_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_62_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_62_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_62_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_62_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_63_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_63_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_63_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_63_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_63_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_64_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_64_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_64_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_64_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_64_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_65_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_65_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_65_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_65_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_65_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_66_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_66_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_66_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_66_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_66_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_67_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_67_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_67_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_67_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_67_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_68_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_68_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_68_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_68_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_68_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_69_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_69_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_69_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_69_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_69_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_70_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_70_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_70_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_70_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_70_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_71_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_71_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_71_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_71_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_71_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_72_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_72_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_72_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_72_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_72_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_73_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_73_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_73_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_73_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_73_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_74_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_74_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_74_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_74_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_74_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_75_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_75_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_75_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_75_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_75_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_76_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_76_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_76_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_76_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_76_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_77_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_77_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_77_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_77_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_77_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_78_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_78_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_78_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_78_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_78_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_79_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_79_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_79_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_79_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_79_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_80_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_80_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_80_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_80_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_80_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_81_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_81_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_81_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_81_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_81_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_82_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_82_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_82_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_82_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_82_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_83_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_83_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_83_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_83_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_83_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_84_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_84_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_84_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_84_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_84_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_85_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_85_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_85_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_85_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_85_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_86_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_86_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_86_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_86_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_86_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_87_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_87_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_87_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_87_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_87_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_88_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_88_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_88_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_88_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_88_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_89_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_89_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_89_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_89_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_89_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_90_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_90_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_90_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_90_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_90_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_91_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_91_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_91_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_91_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_91_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_92_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_92_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_92_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_92_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_92_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_93_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_93_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_93_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_93_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_93_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_94_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_94_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_94_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_94_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_94_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_95_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_95_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_95_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_95_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_95_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_96_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_96_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_96_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_96_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_96_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_97_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_97_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_97_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_97_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_97_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_98_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_98_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_98_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_98_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_98_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_99_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_99_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_99_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_99_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_99_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_100_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_100_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_100_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_100_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_100_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_101_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_101_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_101_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_101_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_101_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_102_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_102_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_102_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_102_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_102_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_103_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_103_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_103_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_103_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_103_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_104_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_104_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_104_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_104_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_104_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_105_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_105_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_105_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_105_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_105_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_106_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_106_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_106_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_106_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_106_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_107_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_107_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_107_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_107_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_107_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_108_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_108_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_108_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_108_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_108_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_109_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_109_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_109_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_109_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_109_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_110_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_110_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_110_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_110_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_110_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_111_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_111_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_111_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_111_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_111_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_112_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_112_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_112_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_112_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_112_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_113_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_113_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_113_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_113_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_113_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_114_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_114_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_114_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_114_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_114_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_115_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_115_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_115_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_115_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_115_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_116_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_116_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_116_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_116_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_116_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_117_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_117_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_117_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_117_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_117_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_118_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_118_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_118_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_118_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_118_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_119_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_119_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_119_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_119_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_119_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_120_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_120_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_120_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_120_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_120_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_121_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_121_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_121_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_121_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_121_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_122_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_122_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_122_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_122_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_122_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_123_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_123_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_123_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_123_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_123_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_124_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_124_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_124_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_124_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_124_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_125_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_125_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_125_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_125_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_125_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_126_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_126_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_126_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_126_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_126_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_127_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_127_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_127_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_127_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_127_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_128_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_128_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_128_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_128_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_128_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_129_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_129_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_129_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_129_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_129_io_o_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_130_io_i_inter_c; // @[wallace_tree.scala 137:50]
  wire [21:0] wallace_tree_cells_130_io_i_s; // @[wallace_tree.scala 137:50]
  wire [18:0] wallace_tree_cells_130_io_o_inter_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_130_io_o_c; // @[wallace_tree.scala 137:50]
  wire  wallace_tree_cells_130_io_o_s; // @[wallace_tree.scala 137:50]
  wire  inversed_pp_0_0 = io_i_partial_products_0[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_0 = io_i_partial_products_0[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_0 = io_i_partial_products_0[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_0 = io_i_partial_products_0[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_0 = io_i_partial_products_0[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_0 = io_i_partial_products_0[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_0 = io_i_partial_products_0[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_0 = io_i_partial_products_0[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_0 = io_i_partial_products_0[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_0 = io_i_partial_products_0[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_0 = io_i_partial_products_0[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_0 = io_i_partial_products_0[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_0 = io_i_partial_products_0[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_0 = io_i_partial_products_0[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_0 = io_i_partial_products_0[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_0 = io_i_partial_products_0[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_0 = io_i_partial_products_0[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_0 = io_i_partial_products_0[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_0 = io_i_partial_products_0[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_0 = io_i_partial_products_0[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_0 = io_i_partial_products_0[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_0 = io_i_partial_products_0[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_0 = io_i_partial_products_0[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_0 = io_i_partial_products_0[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_0 = io_i_partial_products_0[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_0 = io_i_partial_products_0[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_0 = io_i_partial_products_0[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_0 = io_i_partial_products_0[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_0 = io_i_partial_products_0[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_0 = io_i_partial_products_0[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_0 = io_i_partial_products_0[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_0 = io_i_partial_products_0[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_0 = io_i_partial_products_0[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_0 = io_i_partial_products_0[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_0 = io_i_partial_products_0[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_0 = io_i_partial_products_0[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_0 = io_i_partial_products_0[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_0 = io_i_partial_products_0[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_0 = io_i_partial_products_0[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_0 = io_i_partial_products_0[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_0 = io_i_partial_products_0[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_0 = io_i_partial_products_0[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_0 = io_i_partial_products_0[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_0 = io_i_partial_products_0[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_0 = io_i_partial_products_0[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_0 = io_i_partial_products_0[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_0 = io_i_partial_products_0[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_0 = io_i_partial_products_0[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_0 = io_i_partial_products_0[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_0 = io_i_partial_products_0[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_0 = io_i_partial_products_0[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_0 = io_i_partial_products_0[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_0 = io_i_partial_products_0[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_0 = io_i_partial_products_0[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_0 = io_i_partial_products_0[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_0 = io_i_partial_products_0[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_0 = io_i_partial_products_0[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_0 = io_i_partial_products_0[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_0 = io_i_partial_products_0[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_0 = io_i_partial_products_0[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_0 = io_i_partial_products_0[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_0 = io_i_partial_products_0[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_0 = io_i_partial_products_0[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_0 = io_i_partial_products_0[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_0 = io_i_partial_products_0[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_0 = io_i_partial_products_0[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_0 = io_i_partial_products_0[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_0 = io_i_partial_products_0[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_0 = io_i_partial_products_0[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_0 = io_i_partial_products_0[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_0 = io_i_partial_products_0[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_0 = io_i_partial_products_0[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_0 = io_i_partial_products_0[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_0 = io_i_partial_products_0[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_0 = io_i_partial_products_0[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_0 = io_i_partial_products_0[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_0 = io_i_partial_products_0[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_0 = io_i_partial_products_0[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_0 = io_i_partial_products_0[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_0 = io_i_partial_products_0[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_0 = io_i_partial_products_0[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_0 = io_i_partial_products_0[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_0 = io_i_partial_products_0[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_0 = io_i_partial_products_0[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_0 = io_i_partial_products_0[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_0 = io_i_partial_products_0[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_0 = io_i_partial_products_0[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_0 = io_i_partial_products_0[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_0 = io_i_partial_products_0[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_0 = io_i_partial_products_0[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_0 = io_i_partial_products_0[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_0 = io_i_partial_products_0[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_0 = io_i_partial_products_0[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_0 = io_i_partial_products_0[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_0 = io_i_partial_products_0[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_0 = io_i_partial_products_0[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_0 = io_i_partial_products_0[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_0 = io_i_partial_products_0[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_0 = io_i_partial_products_0[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_0 = io_i_partial_products_0[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_0 = io_i_partial_products_0[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_0 = io_i_partial_products_0[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_0 = io_i_partial_products_0[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_0 = io_i_partial_products_0[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_0 = io_i_partial_products_0[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_0 = io_i_partial_products_0[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_0 = io_i_partial_products_0[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_0 = io_i_partial_products_0[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_0 = io_i_partial_products_0[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_0 = io_i_partial_products_0[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_0 = io_i_partial_products_0[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_0 = io_i_partial_products_0[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_0 = io_i_partial_products_0[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_0 = io_i_partial_products_0[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_0 = io_i_partial_products_0[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_0 = io_i_partial_products_0[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_0 = io_i_partial_products_0[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_0 = io_i_partial_products_0[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_0 = io_i_partial_products_0[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_0 = io_i_partial_products_0[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_0 = io_i_partial_products_0[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_0 = io_i_partial_products_0[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_0 = io_i_partial_products_0[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_0 = io_i_partial_products_0[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_0 = io_i_partial_products_0[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_0 = io_i_partial_products_0[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_0 = io_i_partial_products_0[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_0 = io_i_partial_products_0[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_0 = io_i_partial_products_0[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_0 = io_i_partial_products_0[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_0 = io_i_partial_products_0[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_1 = io_i_partial_products_1[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_1 = io_i_partial_products_1[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_1 = io_i_partial_products_1[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_1 = io_i_partial_products_1[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_1 = io_i_partial_products_1[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_1 = io_i_partial_products_1[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_1 = io_i_partial_products_1[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_1 = io_i_partial_products_1[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_1 = io_i_partial_products_1[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_1 = io_i_partial_products_1[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_1 = io_i_partial_products_1[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_1 = io_i_partial_products_1[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_1 = io_i_partial_products_1[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_1 = io_i_partial_products_1[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_1 = io_i_partial_products_1[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_1 = io_i_partial_products_1[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_1 = io_i_partial_products_1[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_1 = io_i_partial_products_1[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_1 = io_i_partial_products_1[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_1 = io_i_partial_products_1[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_1 = io_i_partial_products_1[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_1 = io_i_partial_products_1[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_1 = io_i_partial_products_1[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_1 = io_i_partial_products_1[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_1 = io_i_partial_products_1[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_1 = io_i_partial_products_1[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_1 = io_i_partial_products_1[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_1 = io_i_partial_products_1[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_1 = io_i_partial_products_1[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_1 = io_i_partial_products_1[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_1 = io_i_partial_products_1[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_1 = io_i_partial_products_1[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_1 = io_i_partial_products_1[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_1 = io_i_partial_products_1[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_1 = io_i_partial_products_1[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_1 = io_i_partial_products_1[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_1 = io_i_partial_products_1[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_1 = io_i_partial_products_1[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_1 = io_i_partial_products_1[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_1 = io_i_partial_products_1[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_1 = io_i_partial_products_1[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_1 = io_i_partial_products_1[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_1 = io_i_partial_products_1[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_1 = io_i_partial_products_1[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_1 = io_i_partial_products_1[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_1 = io_i_partial_products_1[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_1 = io_i_partial_products_1[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_1 = io_i_partial_products_1[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_1 = io_i_partial_products_1[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_1 = io_i_partial_products_1[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_1 = io_i_partial_products_1[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_1 = io_i_partial_products_1[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_1 = io_i_partial_products_1[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_1 = io_i_partial_products_1[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_1 = io_i_partial_products_1[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_1 = io_i_partial_products_1[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_1 = io_i_partial_products_1[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_1 = io_i_partial_products_1[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_1 = io_i_partial_products_1[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_1 = io_i_partial_products_1[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_1 = io_i_partial_products_1[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_1 = io_i_partial_products_1[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_1 = io_i_partial_products_1[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_1 = io_i_partial_products_1[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_1 = io_i_partial_products_1[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_1 = io_i_partial_products_1[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_1 = io_i_partial_products_1[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_1 = io_i_partial_products_1[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_1 = io_i_partial_products_1[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_1 = io_i_partial_products_1[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_1 = io_i_partial_products_1[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_1 = io_i_partial_products_1[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_1 = io_i_partial_products_1[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_1 = io_i_partial_products_1[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_1 = io_i_partial_products_1[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_1 = io_i_partial_products_1[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_1 = io_i_partial_products_1[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_1 = io_i_partial_products_1[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_1 = io_i_partial_products_1[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_1 = io_i_partial_products_1[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_1 = io_i_partial_products_1[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_1 = io_i_partial_products_1[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_1 = io_i_partial_products_1[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_1 = io_i_partial_products_1[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_1 = io_i_partial_products_1[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_1 = io_i_partial_products_1[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_1 = io_i_partial_products_1[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_1 = io_i_partial_products_1[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_1 = io_i_partial_products_1[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_1 = io_i_partial_products_1[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_1 = io_i_partial_products_1[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_1 = io_i_partial_products_1[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_1 = io_i_partial_products_1[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_1 = io_i_partial_products_1[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_1 = io_i_partial_products_1[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_1 = io_i_partial_products_1[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_1 = io_i_partial_products_1[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_1 = io_i_partial_products_1[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_1 = io_i_partial_products_1[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_1 = io_i_partial_products_1[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_1 = io_i_partial_products_1[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_1 = io_i_partial_products_1[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_1 = io_i_partial_products_1[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_1 = io_i_partial_products_1[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_1 = io_i_partial_products_1[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_1 = io_i_partial_products_1[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_1 = io_i_partial_products_1[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_1 = io_i_partial_products_1[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_1 = io_i_partial_products_1[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_1 = io_i_partial_products_1[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_1 = io_i_partial_products_1[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_1 = io_i_partial_products_1[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_1 = io_i_partial_products_1[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_1 = io_i_partial_products_1[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_1 = io_i_partial_products_1[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_1 = io_i_partial_products_1[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_1 = io_i_partial_products_1[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_1 = io_i_partial_products_1[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_1 = io_i_partial_products_1[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_1 = io_i_partial_products_1[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_1 = io_i_partial_products_1[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_1 = io_i_partial_products_1[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_1 = io_i_partial_products_1[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_1 = io_i_partial_products_1[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_1 = io_i_partial_products_1[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_1 = io_i_partial_products_1[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_1 = io_i_partial_products_1[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_1 = io_i_partial_products_1[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_1 = io_i_partial_products_1[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_1 = io_i_partial_products_1[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_1 = io_i_partial_products_1[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_2 = io_i_partial_products_2[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_2 = io_i_partial_products_2[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_2 = io_i_partial_products_2[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_2 = io_i_partial_products_2[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_2 = io_i_partial_products_2[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_2 = io_i_partial_products_2[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_2 = io_i_partial_products_2[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_2 = io_i_partial_products_2[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_2 = io_i_partial_products_2[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_2 = io_i_partial_products_2[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_2 = io_i_partial_products_2[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_2 = io_i_partial_products_2[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_2 = io_i_partial_products_2[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_2 = io_i_partial_products_2[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_2 = io_i_partial_products_2[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_2 = io_i_partial_products_2[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_2 = io_i_partial_products_2[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_2 = io_i_partial_products_2[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_2 = io_i_partial_products_2[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_2 = io_i_partial_products_2[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_2 = io_i_partial_products_2[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_2 = io_i_partial_products_2[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_2 = io_i_partial_products_2[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_2 = io_i_partial_products_2[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_2 = io_i_partial_products_2[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_2 = io_i_partial_products_2[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_2 = io_i_partial_products_2[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_2 = io_i_partial_products_2[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_2 = io_i_partial_products_2[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_2 = io_i_partial_products_2[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_2 = io_i_partial_products_2[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_2 = io_i_partial_products_2[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_2 = io_i_partial_products_2[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_2 = io_i_partial_products_2[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_2 = io_i_partial_products_2[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_2 = io_i_partial_products_2[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_2 = io_i_partial_products_2[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_2 = io_i_partial_products_2[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_2 = io_i_partial_products_2[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_2 = io_i_partial_products_2[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_2 = io_i_partial_products_2[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_2 = io_i_partial_products_2[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_2 = io_i_partial_products_2[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_2 = io_i_partial_products_2[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_2 = io_i_partial_products_2[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_2 = io_i_partial_products_2[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_2 = io_i_partial_products_2[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_2 = io_i_partial_products_2[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_2 = io_i_partial_products_2[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_2 = io_i_partial_products_2[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_2 = io_i_partial_products_2[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_2 = io_i_partial_products_2[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_2 = io_i_partial_products_2[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_2 = io_i_partial_products_2[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_2 = io_i_partial_products_2[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_2 = io_i_partial_products_2[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_2 = io_i_partial_products_2[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_2 = io_i_partial_products_2[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_2 = io_i_partial_products_2[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_2 = io_i_partial_products_2[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_2 = io_i_partial_products_2[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_2 = io_i_partial_products_2[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_2 = io_i_partial_products_2[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_2 = io_i_partial_products_2[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_2 = io_i_partial_products_2[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_2 = io_i_partial_products_2[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_2 = io_i_partial_products_2[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_2 = io_i_partial_products_2[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_2 = io_i_partial_products_2[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_2 = io_i_partial_products_2[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_2 = io_i_partial_products_2[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_2 = io_i_partial_products_2[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_2 = io_i_partial_products_2[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_2 = io_i_partial_products_2[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_2 = io_i_partial_products_2[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_2 = io_i_partial_products_2[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_2 = io_i_partial_products_2[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_2 = io_i_partial_products_2[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_2 = io_i_partial_products_2[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_2 = io_i_partial_products_2[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_2 = io_i_partial_products_2[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_2 = io_i_partial_products_2[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_2 = io_i_partial_products_2[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_2 = io_i_partial_products_2[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_2 = io_i_partial_products_2[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_2 = io_i_partial_products_2[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_2 = io_i_partial_products_2[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_2 = io_i_partial_products_2[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_2 = io_i_partial_products_2[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_2 = io_i_partial_products_2[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_2 = io_i_partial_products_2[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_2 = io_i_partial_products_2[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_2 = io_i_partial_products_2[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_2 = io_i_partial_products_2[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_2 = io_i_partial_products_2[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_2 = io_i_partial_products_2[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_2 = io_i_partial_products_2[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_2 = io_i_partial_products_2[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_2 = io_i_partial_products_2[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_2 = io_i_partial_products_2[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_2 = io_i_partial_products_2[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_2 = io_i_partial_products_2[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_2 = io_i_partial_products_2[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_2 = io_i_partial_products_2[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_2 = io_i_partial_products_2[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_2 = io_i_partial_products_2[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_2 = io_i_partial_products_2[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_2 = io_i_partial_products_2[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_2 = io_i_partial_products_2[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_2 = io_i_partial_products_2[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_2 = io_i_partial_products_2[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_2 = io_i_partial_products_2[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_2 = io_i_partial_products_2[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_2 = io_i_partial_products_2[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_2 = io_i_partial_products_2[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_2 = io_i_partial_products_2[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_2 = io_i_partial_products_2[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_2 = io_i_partial_products_2[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_2 = io_i_partial_products_2[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_2 = io_i_partial_products_2[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_2 = io_i_partial_products_2[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_2 = io_i_partial_products_2[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_2 = io_i_partial_products_2[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_2 = io_i_partial_products_2[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_2 = io_i_partial_products_2[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_2 = io_i_partial_products_2[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_2 = io_i_partial_products_2[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_2 = io_i_partial_products_2[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_2 = io_i_partial_products_2[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_2 = io_i_partial_products_2[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_2 = io_i_partial_products_2[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_3 = io_i_partial_products_3[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_3 = io_i_partial_products_3[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_3 = io_i_partial_products_3[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_3 = io_i_partial_products_3[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_3 = io_i_partial_products_3[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_3 = io_i_partial_products_3[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_3 = io_i_partial_products_3[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_3 = io_i_partial_products_3[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_3 = io_i_partial_products_3[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_3 = io_i_partial_products_3[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_3 = io_i_partial_products_3[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_3 = io_i_partial_products_3[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_3 = io_i_partial_products_3[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_3 = io_i_partial_products_3[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_3 = io_i_partial_products_3[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_3 = io_i_partial_products_3[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_3 = io_i_partial_products_3[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_3 = io_i_partial_products_3[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_3 = io_i_partial_products_3[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_3 = io_i_partial_products_3[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_3 = io_i_partial_products_3[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_3 = io_i_partial_products_3[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_3 = io_i_partial_products_3[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_3 = io_i_partial_products_3[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_3 = io_i_partial_products_3[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_3 = io_i_partial_products_3[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_3 = io_i_partial_products_3[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_3 = io_i_partial_products_3[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_3 = io_i_partial_products_3[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_3 = io_i_partial_products_3[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_3 = io_i_partial_products_3[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_3 = io_i_partial_products_3[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_3 = io_i_partial_products_3[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_3 = io_i_partial_products_3[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_3 = io_i_partial_products_3[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_3 = io_i_partial_products_3[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_3 = io_i_partial_products_3[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_3 = io_i_partial_products_3[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_3 = io_i_partial_products_3[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_3 = io_i_partial_products_3[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_3 = io_i_partial_products_3[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_3 = io_i_partial_products_3[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_3 = io_i_partial_products_3[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_3 = io_i_partial_products_3[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_3 = io_i_partial_products_3[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_3 = io_i_partial_products_3[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_3 = io_i_partial_products_3[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_3 = io_i_partial_products_3[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_3 = io_i_partial_products_3[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_3 = io_i_partial_products_3[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_3 = io_i_partial_products_3[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_3 = io_i_partial_products_3[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_3 = io_i_partial_products_3[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_3 = io_i_partial_products_3[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_3 = io_i_partial_products_3[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_3 = io_i_partial_products_3[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_3 = io_i_partial_products_3[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_3 = io_i_partial_products_3[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_3 = io_i_partial_products_3[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_3 = io_i_partial_products_3[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_3 = io_i_partial_products_3[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_3 = io_i_partial_products_3[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_3 = io_i_partial_products_3[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_3 = io_i_partial_products_3[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_3 = io_i_partial_products_3[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_3 = io_i_partial_products_3[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_3 = io_i_partial_products_3[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_3 = io_i_partial_products_3[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_3 = io_i_partial_products_3[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_3 = io_i_partial_products_3[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_3 = io_i_partial_products_3[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_3 = io_i_partial_products_3[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_3 = io_i_partial_products_3[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_3 = io_i_partial_products_3[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_3 = io_i_partial_products_3[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_3 = io_i_partial_products_3[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_3 = io_i_partial_products_3[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_3 = io_i_partial_products_3[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_3 = io_i_partial_products_3[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_3 = io_i_partial_products_3[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_3 = io_i_partial_products_3[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_3 = io_i_partial_products_3[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_3 = io_i_partial_products_3[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_3 = io_i_partial_products_3[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_3 = io_i_partial_products_3[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_3 = io_i_partial_products_3[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_3 = io_i_partial_products_3[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_3 = io_i_partial_products_3[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_3 = io_i_partial_products_3[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_3 = io_i_partial_products_3[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_3 = io_i_partial_products_3[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_3 = io_i_partial_products_3[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_3 = io_i_partial_products_3[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_3 = io_i_partial_products_3[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_3 = io_i_partial_products_3[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_3 = io_i_partial_products_3[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_3 = io_i_partial_products_3[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_3 = io_i_partial_products_3[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_3 = io_i_partial_products_3[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_3 = io_i_partial_products_3[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_3 = io_i_partial_products_3[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_3 = io_i_partial_products_3[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_3 = io_i_partial_products_3[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_3 = io_i_partial_products_3[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_3 = io_i_partial_products_3[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_3 = io_i_partial_products_3[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_3 = io_i_partial_products_3[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_3 = io_i_partial_products_3[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_3 = io_i_partial_products_3[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_3 = io_i_partial_products_3[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_3 = io_i_partial_products_3[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_3 = io_i_partial_products_3[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_3 = io_i_partial_products_3[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_3 = io_i_partial_products_3[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_3 = io_i_partial_products_3[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_3 = io_i_partial_products_3[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_3 = io_i_partial_products_3[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_3 = io_i_partial_products_3[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_3 = io_i_partial_products_3[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_3 = io_i_partial_products_3[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_3 = io_i_partial_products_3[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_3 = io_i_partial_products_3[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_3 = io_i_partial_products_3[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_3 = io_i_partial_products_3[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_3 = io_i_partial_products_3[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_3 = io_i_partial_products_3[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_3 = io_i_partial_products_3[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_3 = io_i_partial_products_3[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_3 = io_i_partial_products_3[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_3 = io_i_partial_products_3[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_3 = io_i_partial_products_3[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_4 = io_i_partial_products_4[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_4 = io_i_partial_products_4[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_4 = io_i_partial_products_4[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_4 = io_i_partial_products_4[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_4 = io_i_partial_products_4[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_4 = io_i_partial_products_4[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_4 = io_i_partial_products_4[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_4 = io_i_partial_products_4[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_4 = io_i_partial_products_4[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_4 = io_i_partial_products_4[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_4 = io_i_partial_products_4[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_4 = io_i_partial_products_4[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_4 = io_i_partial_products_4[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_4 = io_i_partial_products_4[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_4 = io_i_partial_products_4[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_4 = io_i_partial_products_4[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_4 = io_i_partial_products_4[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_4 = io_i_partial_products_4[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_4 = io_i_partial_products_4[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_4 = io_i_partial_products_4[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_4 = io_i_partial_products_4[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_4 = io_i_partial_products_4[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_4 = io_i_partial_products_4[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_4 = io_i_partial_products_4[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_4 = io_i_partial_products_4[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_4 = io_i_partial_products_4[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_4 = io_i_partial_products_4[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_4 = io_i_partial_products_4[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_4 = io_i_partial_products_4[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_4 = io_i_partial_products_4[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_4 = io_i_partial_products_4[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_4 = io_i_partial_products_4[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_4 = io_i_partial_products_4[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_4 = io_i_partial_products_4[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_4 = io_i_partial_products_4[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_4 = io_i_partial_products_4[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_4 = io_i_partial_products_4[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_4 = io_i_partial_products_4[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_4 = io_i_partial_products_4[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_4 = io_i_partial_products_4[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_4 = io_i_partial_products_4[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_4 = io_i_partial_products_4[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_4 = io_i_partial_products_4[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_4 = io_i_partial_products_4[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_4 = io_i_partial_products_4[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_4 = io_i_partial_products_4[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_4 = io_i_partial_products_4[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_4 = io_i_partial_products_4[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_4 = io_i_partial_products_4[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_4 = io_i_partial_products_4[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_4 = io_i_partial_products_4[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_4 = io_i_partial_products_4[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_4 = io_i_partial_products_4[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_4 = io_i_partial_products_4[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_4 = io_i_partial_products_4[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_4 = io_i_partial_products_4[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_4 = io_i_partial_products_4[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_4 = io_i_partial_products_4[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_4 = io_i_partial_products_4[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_4 = io_i_partial_products_4[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_4 = io_i_partial_products_4[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_4 = io_i_partial_products_4[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_4 = io_i_partial_products_4[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_4 = io_i_partial_products_4[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_4 = io_i_partial_products_4[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_4 = io_i_partial_products_4[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_4 = io_i_partial_products_4[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_4 = io_i_partial_products_4[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_4 = io_i_partial_products_4[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_4 = io_i_partial_products_4[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_4 = io_i_partial_products_4[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_4 = io_i_partial_products_4[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_4 = io_i_partial_products_4[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_4 = io_i_partial_products_4[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_4 = io_i_partial_products_4[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_4 = io_i_partial_products_4[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_4 = io_i_partial_products_4[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_4 = io_i_partial_products_4[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_4 = io_i_partial_products_4[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_4 = io_i_partial_products_4[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_4 = io_i_partial_products_4[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_4 = io_i_partial_products_4[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_4 = io_i_partial_products_4[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_4 = io_i_partial_products_4[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_4 = io_i_partial_products_4[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_4 = io_i_partial_products_4[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_4 = io_i_partial_products_4[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_4 = io_i_partial_products_4[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_4 = io_i_partial_products_4[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_4 = io_i_partial_products_4[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_4 = io_i_partial_products_4[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_4 = io_i_partial_products_4[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_4 = io_i_partial_products_4[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_4 = io_i_partial_products_4[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_4 = io_i_partial_products_4[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_4 = io_i_partial_products_4[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_4 = io_i_partial_products_4[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_4 = io_i_partial_products_4[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_4 = io_i_partial_products_4[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_4 = io_i_partial_products_4[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_4 = io_i_partial_products_4[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_4 = io_i_partial_products_4[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_4 = io_i_partial_products_4[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_4 = io_i_partial_products_4[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_4 = io_i_partial_products_4[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_4 = io_i_partial_products_4[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_4 = io_i_partial_products_4[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_4 = io_i_partial_products_4[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_4 = io_i_partial_products_4[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_4 = io_i_partial_products_4[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_4 = io_i_partial_products_4[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_4 = io_i_partial_products_4[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_4 = io_i_partial_products_4[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_4 = io_i_partial_products_4[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_4 = io_i_partial_products_4[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_4 = io_i_partial_products_4[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_4 = io_i_partial_products_4[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_4 = io_i_partial_products_4[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_4 = io_i_partial_products_4[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_4 = io_i_partial_products_4[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_4 = io_i_partial_products_4[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_4 = io_i_partial_products_4[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_4 = io_i_partial_products_4[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_4 = io_i_partial_products_4[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_4 = io_i_partial_products_4[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_4 = io_i_partial_products_4[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_4 = io_i_partial_products_4[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_4 = io_i_partial_products_4[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_4 = io_i_partial_products_4[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_4 = io_i_partial_products_4[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_4 = io_i_partial_products_4[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_5 = io_i_partial_products_5[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_5 = io_i_partial_products_5[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_5 = io_i_partial_products_5[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_5 = io_i_partial_products_5[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_5 = io_i_partial_products_5[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_5 = io_i_partial_products_5[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_5 = io_i_partial_products_5[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_5 = io_i_partial_products_5[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_5 = io_i_partial_products_5[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_5 = io_i_partial_products_5[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_5 = io_i_partial_products_5[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_5 = io_i_partial_products_5[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_5 = io_i_partial_products_5[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_5 = io_i_partial_products_5[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_5 = io_i_partial_products_5[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_5 = io_i_partial_products_5[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_5 = io_i_partial_products_5[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_5 = io_i_partial_products_5[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_5 = io_i_partial_products_5[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_5 = io_i_partial_products_5[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_5 = io_i_partial_products_5[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_5 = io_i_partial_products_5[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_5 = io_i_partial_products_5[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_5 = io_i_partial_products_5[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_5 = io_i_partial_products_5[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_5 = io_i_partial_products_5[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_5 = io_i_partial_products_5[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_5 = io_i_partial_products_5[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_5 = io_i_partial_products_5[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_5 = io_i_partial_products_5[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_5 = io_i_partial_products_5[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_5 = io_i_partial_products_5[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_5 = io_i_partial_products_5[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_5 = io_i_partial_products_5[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_5 = io_i_partial_products_5[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_5 = io_i_partial_products_5[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_5 = io_i_partial_products_5[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_5 = io_i_partial_products_5[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_5 = io_i_partial_products_5[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_5 = io_i_partial_products_5[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_5 = io_i_partial_products_5[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_5 = io_i_partial_products_5[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_5 = io_i_partial_products_5[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_5 = io_i_partial_products_5[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_5 = io_i_partial_products_5[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_5 = io_i_partial_products_5[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_5 = io_i_partial_products_5[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_5 = io_i_partial_products_5[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_5 = io_i_partial_products_5[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_5 = io_i_partial_products_5[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_5 = io_i_partial_products_5[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_5 = io_i_partial_products_5[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_5 = io_i_partial_products_5[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_5 = io_i_partial_products_5[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_5 = io_i_partial_products_5[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_5 = io_i_partial_products_5[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_5 = io_i_partial_products_5[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_5 = io_i_partial_products_5[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_5 = io_i_partial_products_5[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_5 = io_i_partial_products_5[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_5 = io_i_partial_products_5[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_5 = io_i_partial_products_5[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_5 = io_i_partial_products_5[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_5 = io_i_partial_products_5[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_5 = io_i_partial_products_5[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_5 = io_i_partial_products_5[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_5 = io_i_partial_products_5[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_5 = io_i_partial_products_5[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_5 = io_i_partial_products_5[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_5 = io_i_partial_products_5[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_5 = io_i_partial_products_5[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_5 = io_i_partial_products_5[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_5 = io_i_partial_products_5[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_5 = io_i_partial_products_5[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_5 = io_i_partial_products_5[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_5 = io_i_partial_products_5[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_5 = io_i_partial_products_5[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_5 = io_i_partial_products_5[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_5 = io_i_partial_products_5[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_5 = io_i_partial_products_5[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_5 = io_i_partial_products_5[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_5 = io_i_partial_products_5[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_5 = io_i_partial_products_5[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_5 = io_i_partial_products_5[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_5 = io_i_partial_products_5[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_5 = io_i_partial_products_5[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_5 = io_i_partial_products_5[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_5 = io_i_partial_products_5[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_5 = io_i_partial_products_5[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_5 = io_i_partial_products_5[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_5 = io_i_partial_products_5[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_5 = io_i_partial_products_5[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_5 = io_i_partial_products_5[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_5 = io_i_partial_products_5[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_5 = io_i_partial_products_5[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_5 = io_i_partial_products_5[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_5 = io_i_partial_products_5[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_5 = io_i_partial_products_5[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_5 = io_i_partial_products_5[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_5 = io_i_partial_products_5[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_5 = io_i_partial_products_5[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_5 = io_i_partial_products_5[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_5 = io_i_partial_products_5[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_5 = io_i_partial_products_5[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_5 = io_i_partial_products_5[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_5 = io_i_partial_products_5[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_5 = io_i_partial_products_5[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_5 = io_i_partial_products_5[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_5 = io_i_partial_products_5[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_5 = io_i_partial_products_5[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_5 = io_i_partial_products_5[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_5 = io_i_partial_products_5[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_5 = io_i_partial_products_5[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_5 = io_i_partial_products_5[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_5 = io_i_partial_products_5[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_5 = io_i_partial_products_5[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_5 = io_i_partial_products_5[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_5 = io_i_partial_products_5[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_5 = io_i_partial_products_5[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_5 = io_i_partial_products_5[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_5 = io_i_partial_products_5[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_5 = io_i_partial_products_5[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_5 = io_i_partial_products_5[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_5 = io_i_partial_products_5[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_5 = io_i_partial_products_5[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_5 = io_i_partial_products_5[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_5 = io_i_partial_products_5[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_5 = io_i_partial_products_5[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_5 = io_i_partial_products_5[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_5 = io_i_partial_products_5[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_5 = io_i_partial_products_5[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_6 = io_i_partial_products_6[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_6 = io_i_partial_products_6[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_6 = io_i_partial_products_6[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_6 = io_i_partial_products_6[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_6 = io_i_partial_products_6[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_6 = io_i_partial_products_6[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_6 = io_i_partial_products_6[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_6 = io_i_partial_products_6[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_6 = io_i_partial_products_6[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_6 = io_i_partial_products_6[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_6 = io_i_partial_products_6[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_6 = io_i_partial_products_6[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_6 = io_i_partial_products_6[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_6 = io_i_partial_products_6[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_6 = io_i_partial_products_6[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_6 = io_i_partial_products_6[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_6 = io_i_partial_products_6[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_6 = io_i_partial_products_6[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_6 = io_i_partial_products_6[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_6 = io_i_partial_products_6[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_6 = io_i_partial_products_6[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_6 = io_i_partial_products_6[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_6 = io_i_partial_products_6[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_6 = io_i_partial_products_6[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_6 = io_i_partial_products_6[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_6 = io_i_partial_products_6[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_6 = io_i_partial_products_6[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_6 = io_i_partial_products_6[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_6 = io_i_partial_products_6[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_6 = io_i_partial_products_6[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_6 = io_i_partial_products_6[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_6 = io_i_partial_products_6[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_6 = io_i_partial_products_6[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_6 = io_i_partial_products_6[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_6 = io_i_partial_products_6[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_6 = io_i_partial_products_6[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_6 = io_i_partial_products_6[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_6 = io_i_partial_products_6[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_6 = io_i_partial_products_6[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_6 = io_i_partial_products_6[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_6 = io_i_partial_products_6[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_6 = io_i_partial_products_6[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_6 = io_i_partial_products_6[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_6 = io_i_partial_products_6[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_6 = io_i_partial_products_6[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_6 = io_i_partial_products_6[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_6 = io_i_partial_products_6[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_6 = io_i_partial_products_6[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_6 = io_i_partial_products_6[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_6 = io_i_partial_products_6[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_6 = io_i_partial_products_6[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_6 = io_i_partial_products_6[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_6 = io_i_partial_products_6[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_6 = io_i_partial_products_6[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_6 = io_i_partial_products_6[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_6 = io_i_partial_products_6[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_6 = io_i_partial_products_6[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_6 = io_i_partial_products_6[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_6 = io_i_partial_products_6[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_6 = io_i_partial_products_6[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_6 = io_i_partial_products_6[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_6 = io_i_partial_products_6[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_6 = io_i_partial_products_6[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_6 = io_i_partial_products_6[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_6 = io_i_partial_products_6[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_6 = io_i_partial_products_6[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_6 = io_i_partial_products_6[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_6 = io_i_partial_products_6[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_6 = io_i_partial_products_6[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_6 = io_i_partial_products_6[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_6 = io_i_partial_products_6[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_6 = io_i_partial_products_6[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_6 = io_i_partial_products_6[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_6 = io_i_partial_products_6[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_6 = io_i_partial_products_6[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_6 = io_i_partial_products_6[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_6 = io_i_partial_products_6[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_6 = io_i_partial_products_6[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_6 = io_i_partial_products_6[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_6 = io_i_partial_products_6[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_6 = io_i_partial_products_6[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_6 = io_i_partial_products_6[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_6 = io_i_partial_products_6[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_6 = io_i_partial_products_6[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_6 = io_i_partial_products_6[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_6 = io_i_partial_products_6[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_6 = io_i_partial_products_6[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_6 = io_i_partial_products_6[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_6 = io_i_partial_products_6[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_6 = io_i_partial_products_6[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_6 = io_i_partial_products_6[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_6 = io_i_partial_products_6[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_6 = io_i_partial_products_6[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_6 = io_i_partial_products_6[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_6 = io_i_partial_products_6[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_6 = io_i_partial_products_6[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_6 = io_i_partial_products_6[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_6 = io_i_partial_products_6[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_6 = io_i_partial_products_6[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_6 = io_i_partial_products_6[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_6 = io_i_partial_products_6[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_6 = io_i_partial_products_6[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_6 = io_i_partial_products_6[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_6 = io_i_partial_products_6[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_6 = io_i_partial_products_6[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_6 = io_i_partial_products_6[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_6 = io_i_partial_products_6[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_6 = io_i_partial_products_6[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_6 = io_i_partial_products_6[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_6 = io_i_partial_products_6[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_6 = io_i_partial_products_6[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_6 = io_i_partial_products_6[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_6 = io_i_partial_products_6[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_6 = io_i_partial_products_6[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_6 = io_i_partial_products_6[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_6 = io_i_partial_products_6[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_6 = io_i_partial_products_6[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_6 = io_i_partial_products_6[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_6 = io_i_partial_products_6[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_6 = io_i_partial_products_6[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_6 = io_i_partial_products_6[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_6 = io_i_partial_products_6[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_6 = io_i_partial_products_6[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_6 = io_i_partial_products_6[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_6 = io_i_partial_products_6[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_6 = io_i_partial_products_6[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_6 = io_i_partial_products_6[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_6 = io_i_partial_products_6[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_6 = io_i_partial_products_6[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_6 = io_i_partial_products_6[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_6 = io_i_partial_products_6[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_7 = io_i_partial_products_7[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_7 = io_i_partial_products_7[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_7 = io_i_partial_products_7[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_7 = io_i_partial_products_7[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_7 = io_i_partial_products_7[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_7 = io_i_partial_products_7[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_7 = io_i_partial_products_7[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_7 = io_i_partial_products_7[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_7 = io_i_partial_products_7[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_7 = io_i_partial_products_7[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_7 = io_i_partial_products_7[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_7 = io_i_partial_products_7[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_7 = io_i_partial_products_7[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_7 = io_i_partial_products_7[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_7 = io_i_partial_products_7[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_7 = io_i_partial_products_7[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_7 = io_i_partial_products_7[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_7 = io_i_partial_products_7[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_7 = io_i_partial_products_7[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_7 = io_i_partial_products_7[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_7 = io_i_partial_products_7[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_7 = io_i_partial_products_7[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_7 = io_i_partial_products_7[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_7 = io_i_partial_products_7[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_7 = io_i_partial_products_7[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_7 = io_i_partial_products_7[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_7 = io_i_partial_products_7[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_7 = io_i_partial_products_7[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_7 = io_i_partial_products_7[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_7 = io_i_partial_products_7[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_7 = io_i_partial_products_7[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_7 = io_i_partial_products_7[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_7 = io_i_partial_products_7[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_7 = io_i_partial_products_7[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_7 = io_i_partial_products_7[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_7 = io_i_partial_products_7[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_7 = io_i_partial_products_7[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_7 = io_i_partial_products_7[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_7 = io_i_partial_products_7[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_7 = io_i_partial_products_7[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_7 = io_i_partial_products_7[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_7 = io_i_partial_products_7[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_7 = io_i_partial_products_7[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_7 = io_i_partial_products_7[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_7 = io_i_partial_products_7[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_7 = io_i_partial_products_7[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_7 = io_i_partial_products_7[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_7 = io_i_partial_products_7[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_7 = io_i_partial_products_7[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_7 = io_i_partial_products_7[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_7 = io_i_partial_products_7[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_7 = io_i_partial_products_7[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_7 = io_i_partial_products_7[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_7 = io_i_partial_products_7[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_7 = io_i_partial_products_7[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_7 = io_i_partial_products_7[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_7 = io_i_partial_products_7[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_7 = io_i_partial_products_7[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_7 = io_i_partial_products_7[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_7 = io_i_partial_products_7[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_7 = io_i_partial_products_7[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_7 = io_i_partial_products_7[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_7 = io_i_partial_products_7[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_7 = io_i_partial_products_7[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_7 = io_i_partial_products_7[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_7 = io_i_partial_products_7[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_7 = io_i_partial_products_7[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_7 = io_i_partial_products_7[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_7 = io_i_partial_products_7[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_7 = io_i_partial_products_7[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_7 = io_i_partial_products_7[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_7 = io_i_partial_products_7[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_7 = io_i_partial_products_7[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_7 = io_i_partial_products_7[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_7 = io_i_partial_products_7[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_7 = io_i_partial_products_7[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_7 = io_i_partial_products_7[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_7 = io_i_partial_products_7[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_7 = io_i_partial_products_7[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_7 = io_i_partial_products_7[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_7 = io_i_partial_products_7[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_7 = io_i_partial_products_7[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_7 = io_i_partial_products_7[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_7 = io_i_partial_products_7[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_7 = io_i_partial_products_7[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_7 = io_i_partial_products_7[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_7 = io_i_partial_products_7[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_7 = io_i_partial_products_7[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_7 = io_i_partial_products_7[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_7 = io_i_partial_products_7[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_7 = io_i_partial_products_7[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_7 = io_i_partial_products_7[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_7 = io_i_partial_products_7[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_7 = io_i_partial_products_7[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_7 = io_i_partial_products_7[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_7 = io_i_partial_products_7[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_7 = io_i_partial_products_7[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_7 = io_i_partial_products_7[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_7 = io_i_partial_products_7[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_7 = io_i_partial_products_7[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_7 = io_i_partial_products_7[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_7 = io_i_partial_products_7[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_7 = io_i_partial_products_7[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_7 = io_i_partial_products_7[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_7 = io_i_partial_products_7[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_7 = io_i_partial_products_7[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_7 = io_i_partial_products_7[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_7 = io_i_partial_products_7[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_7 = io_i_partial_products_7[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_7 = io_i_partial_products_7[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_7 = io_i_partial_products_7[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_7 = io_i_partial_products_7[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_7 = io_i_partial_products_7[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_7 = io_i_partial_products_7[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_7 = io_i_partial_products_7[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_7 = io_i_partial_products_7[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_7 = io_i_partial_products_7[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_7 = io_i_partial_products_7[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_7 = io_i_partial_products_7[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_7 = io_i_partial_products_7[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_7 = io_i_partial_products_7[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_7 = io_i_partial_products_7[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_7 = io_i_partial_products_7[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_7 = io_i_partial_products_7[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_7 = io_i_partial_products_7[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_7 = io_i_partial_products_7[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_7 = io_i_partial_products_7[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_7 = io_i_partial_products_7[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_7 = io_i_partial_products_7[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_7 = io_i_partial_products_7[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_7 = io_i_partial_products_7[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_8 = io_i_partial_products_8[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_8 = io_i_partial_products_8[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_8 = io_i_partial_products_8[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_8 = io_i_partial_products_8[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_8 = io_i_partial_products_8[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_8 = io_i_partial_products_8[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_8 = io_i_partial_products_8[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_8 = io_i_partial_products_8[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_8 = io_i_partial_products_8[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_8 = io_i_partial_products_8[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_8 = io_i_partial_products_8[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_8 = io_i_partial_products_8[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_8 = io_i_partial_products_8[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_8 = io_i_partial_products_8[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_8 = io_i_partial_products_8[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_8 = io_i_partial_products_8[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_8 = io_i_partial_products_8[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_8 = io_i_partial_products_8[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_8 = io_i_partial_products_8[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_8 = io_i_partial_products_8[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_8 = io_i_partial_products_8[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_8 = io_i_partial_products_8[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_8 = io_i_partial_products_8[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_8 = io_i_partial_products_8[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_8 = io_i_partial_products_8[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_8 = io_i_partial_products_8[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_8 = io_i_partial_products_8[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_8 = io_i_partial_products_8[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_8 = io_i_partial_products_8[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_8 = io_i_partial_products_8[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_8 = io_i_partial_products_8[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_8 = io_i_partial_products_8[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_8 = io_i_partial_products_8[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_8 = io_i_partial_products_8[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_8 = io_i_partial_products_8[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_8 = io_i_partial_products_8[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_8 = io_i_partial_products_8[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_8 = io_i_partial_products_8[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_8 = io_i_partial_products_8[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_8 = io_i_partial_products_8[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_8 = io_i_partial_products_8[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_8 = io_i_partial_products_8[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_8 = io_i_partial_products_8[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_8 = io_i_partial_products_8[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_8 = io_i_partial_products_8[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_8 = io_i_partial_products_8[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_8 = io_i_partial_products_8[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_8 = io_i_partial_products_8[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_8 = io_i_partial_products_8[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_8 = io_i_partial_products_8[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_8 = io_i_partial_products_8[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_8 = io_i_partial_products_8[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_8 = io_i_partial_products_8[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_8 = io_i_partial_products_8[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_8 = io_i_partial_products_8[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_8 = io_i_partial_products_8[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_8 = io_i_partial_products_8[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_8 = io_i_partial_products_8[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_8 = io_i_partial_products_8[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_8 = io_i_partial_products_8[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_8 = io_i_partial_products_8[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_8 = io_i_partial_products_8[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_8 = io_i_partial_products_8[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_8 = io_i_partial_products_8[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_8 = io_i_partial_products_8[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_8 = io_i_partial_products_8[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_8 = io_i_partial_products_8[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_8 = io_i_partial_products_8[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_8 = io_i_partial_products_8[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_8 = io_i_partial_products_8[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_8 = io_i_partial_products_8[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_8 = io_i_partial_products_8[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_8 = io_i_partial_products_8[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_8 = io_i_partial_products_8[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_8 = io_i_partial_products_8[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_8 = io_i_partial_products_8[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_8 = io_i_partial_products_8[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_8 = io_i_partial_products_8[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_8 = io_i_partial_products_8[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_8 = io_i_partial_products_8[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_8 = io_i_partial_products_8[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_8 = io_i_partial_products_8[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_8 = io_i_partial_products_8[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_8 = io_i_partial_products_8[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_8 = io_i_partial_products_8[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_8 = io_i_partial_products_8[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_8 = io_i_partial_products_8[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_8 = io_i_partial_products_8[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_8 = io_i_partial_products_8[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_8 = io_i_partial_products_8[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_8 = io_i_partial_products_8[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_8 = io_i_partial_products_8[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_8 = io_i_partial_products_8[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_8 = io_i_partial_products_8[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_8 = io_i_partial_products_8[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_8 = io_i_partial_products_8[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_8 = io_i_partial_products_8[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_8 = io_i_partial_products_8[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_8 = io_i_partial_products_8[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_8 = io_i_partial_products_8[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_8 = io_i_partial_products_8[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_8 = io_i_partial_products_8[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_8 = io_i_partial_products_8[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_8 = io_i_partial_products_8[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_8 = io_i_partial_products_8[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_8 = io_i_partial_products_8[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_8 = io_i_partial_products_8[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_8 = io_i_partial_products_8[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_8 = io_i_partial_products_8[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_8 = io_i_partial_products_8[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_8 = io_i_partial_products_8[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_8 = io_i_partial_products_8[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_8 = io_i_partial_products_8[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_8 = io_i_partial_products_8[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_8 = io_i_partial_products_8[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_8 = io_i_partial_products_8[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_8 = io_i_partial_products_8[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_8 = io_i_partial_products_8[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_8 = io_i_partial_products_8[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_8 = io_i_partial_products_8[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_8 = io_i_partial_products_8[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_8 = io_i_partial_products_8[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_8 = io_i_partial_products_8[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_8 = io_i_partial_products_8[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_8 = io_i_partial_products_8[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_8 = io_i_partial_products_8[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_8 = io_i_partial_products_8[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_8 = io_i_partial_products_8[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_8 = io_i_partial_products_8[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_8 = io_i_partial_products_8[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_8 = io_i_partial_products_8[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_9 = io_i_partial_products_9[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_9 = io_i_partial_products_9[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_9 = io_i_partial_products_9[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_9 = io_i_partial_products_9[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_9 = io_i_partial_products_9[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_9 = io_i_partial_products_9[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_9 = io_i_partial_products_9[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_9 = io_i_partial_products_9[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_9 = io_i_partial_products_9[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_9 = io_i_partial_products_9[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_9 = io_i_partial_products_9[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_9 = io_i_partial_products_9[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_9 = io_i_partial_products_9[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_9 = io_i_partial_products_9[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_9 = io_i_partial_products_9[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_9 = io_i_partial_products_9[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_9 = io_i_partial_products_9[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_9 = io_i_partial_products_9[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_9 = io_i_partial_products_9[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_9 = io_i_partial_products_9[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_9 = io_i_partial_products_9[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_9 = io_i_partial_products_9[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_9 = io_i_partial_products_9[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_9 = io_i_partial_products_9[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_9 = io_i_partial_products_9[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_9 = io_i_partial_products_9[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_9 = io_i_partial_products_9[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_9 = io_i_partial_products_9[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_9 = io_i_partial_products_9[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_9 = io_i_partial_products_9[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_9 = io_i_partial_products_9[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_9 = io_i_partial_products_9[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_9 = io_i_partial_products_9[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_9 = io_i_partial_products_9[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_9 = io_i_partial_products_9[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_9 = io_i_partial_products_9[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_9 = io_i_partial_products_9[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_9 = io_i_partial_products_9[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_9 = io_i_partial_products_9[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_9 = io_i_partial_products_9[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_9 = io_i_partial_products_9[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_9 = io_i_partial_products_9[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_9 = io_i_partial_products_9[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_9 = io_i_partial_products_9[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_9 = io_i_partial_products_9[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_9 = io_i_partial_products_9[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_9 = io_i_partial_products_9[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_9 = io_i_partial_products_9[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_9 = io_i_partial_products_9[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_9 = io_i_partial_products_9[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_9 = io_i_partial_products_9[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_9 = io_i_partial_products_9[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_9 = io_i_partial_products_9[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_9 = io_i_partial_products_9[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_9 = io_i_partial_products_9[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_9 = io_i_partial_products_9[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_9 = io_i_partial_products_9[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_9 = io_i_partial_products_9[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_9 = io_i_partial_products_9[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_9 = io_i_partial_products_9[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_9 = io_i_partial_products_9[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_9 = io_i_partial_products_9[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_9 = io_i_partial_products_9[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_9 = io_i_partial_products_9[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_9 = io_i_partial_products_9[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_9 = io_i_partial_products_9[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_9 = io_i_partial_products_9[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_9 = io_i_partial_products_9[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_9 = io_i_partial_products_9[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_9 = io_i_partial_products_9[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_9 = io_i_partial_products_9[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_9 = io_i_partial_products_9[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_9 = io_i_partial_products_9[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_9 = io_i_partial_products_9[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_9 = io_i_partial_products_9[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_9 = io_i_partial_products_9[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_9 = io_i_partial_products_9[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_9 = io_i_partial_products_9[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_9 = io_i_partial_products_9[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_9 = io_i_partial_products_9[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_9 = io_i_partial_products_9[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_9 = io_i_partial_products_9[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_9 = io_i_partial_products_9[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_9 = io_i_partial_products_9[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_9 = io_i_partial_products_9[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_9 = io_i_partial_products_9[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_9 = io_i_partial_products_9[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_9 = io_i_partial_products_9[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_9 = io_i_partial_products_9[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_9 = io_i_partial_products_9[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_9 = io_i_partial_products_9[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_9 = io_i_partial_products_9[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_9 = io_i_partial_products_9[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_9 = io_i_partial_products_9[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_9 = io_i_partial_products_9[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_9 = io_i_partial_products_9[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_9 = io_i_partial_products_9[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_9 = io_i_partial_products_9[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_9 = io_i_partial_products_9[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_9 = io_i_partial_products_9[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_9 = io_i_partial_products_9[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_9 = io_i_partial_products_9[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_9 = io_i_partial_products_9[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_9 = io_i_partial_products_9[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_9 = io_i_partial_products_9[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_9 = io_i_partial_products_9[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_9 = io_i_partial_products_9[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_9 = io_i_partial_products_9[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_9 = io_i_partial_products_9[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_9 = io_i_partial_products_9[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_9 = io_i_partial_products_9[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_9 = io_i_partial_products_9[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_9 = io_i_partial_products_9[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_9 = io_i_partial_products_9[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_9 = io_i_partial_products_9[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_9 = io_i_partial_products_9[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_9 = io_i_partial_products_9[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_9 = io_i_partial_products_9[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_9 = io_i_partial_products_9[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_9 = io_i_partial_products_9[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_9 = io_i_partial_products_9[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_9 = io_i_partial_products_9[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_9 = io_i_partial_products_9[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_9 = io_i_partial_products_9[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_9 = io_i_partial_products_9[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_9 = io_i_partial_products_9[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_9 = io_i_partial_products_9[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_9 = io_i_partial_products_9[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_9 = io_i_partial_products_9[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_9 = io_i_partial_products_9[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_9 = io_i_partial_products_9[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_10 = io_i_partial_products_10[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_10 = io_i_partial_products_10[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_10 = io_i_partial_products_10[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_10 = io_i_partial_products_10[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_10 = io_i_partial_products_10[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_10 = io_i_partial_products_10[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_10 = io_i_partial_products_10[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_10 = io_i_partial_products_10[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_10 = io_i_partial_products_10[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_10 = io_i_partial_products_10[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_10 = io_i_partial_products_10[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_10 = io_i_partial_products_10[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_10 = io_i_partial_products_10[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_10 = io_i_partial_products_10[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_10 = io_i_partial_products_10[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_10 = io_i_partial_products_10[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_10 = io_i_partial_products_10[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_10 = io_i_partial_products_10[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_10 = io_i_partial_products_10[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_10 = io_i_partial_products_10[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_10 = io_i_partial_products_10[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_10 = io_i_partial_products_10[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_10 = io_i_partial_products_10[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_10 = io_i_partial_products_10[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_10 = io_i_partial_products_10[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_10 = io_i_partial_products_10[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_10 = io_i_partial_products_10[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_10 = io_i_partial_products_10[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_10 = io_i_partial_products_10[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_10 = io_i_partial_products_10[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_10 = io_i_partial_products_10[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_10 = io_i_partial_products_10[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_10 = io_i_partial_products_10[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_10 = io_i_partial_products_10[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_10 = io_i_partial_products_10[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_10 = io_i_partial_products_10[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_10 = io_i_partial_products_10[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_10 = io_i_partial_products_10[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_10 = io_i_partial_products_10[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_10 = io_i_partial_products_10[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_10 = io_i_partial_products_10[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_10 = io_i_partial_products_10[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_10 = io_i_partial_products_10[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_10 = io_i_partial_products_10[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_10 = io_i_partial_products_10[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_10 = io_i_partial_products_10[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_10 = io_i_partial_products_10[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_10 = io_i_partial_products_10[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_10 = io_i_partial_products_10[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_10 = io_i_partial_products_10[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_10 = io_i_partial_products_10[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_10 = io_i_partial_products_10[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_10 = io_i_partial_products_10[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_10 = io_i_partial_products_10[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_10 = io_i_partial_products_10[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_10 = io_i_partial_products_10[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_10 = io_i_partial_products_10[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_10 = io_i_partial_products_10[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_10 = io_i_partial_products_10[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_10 = io_i_partial_products_10[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_10 = io_i_partial_products_10[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_10 = io_i_partial_products_10[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_10 = io_i_partial_products_10[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_10 = io_i_partial_products_10[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_10 = io_i_partial_products_10[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_10 = io_i_partial_products_10[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_10 = io_i_partial_products_10[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_10 = io_i_partial_products_10[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_10 = io_i_partial_products_10[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_10 = io_i_partial_products_10[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_10 = io_i_partial_products_10[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_10 = io_i_partial_products_10[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_10 = io_i_partial_products_10[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_10 = io_i_partial_products_10[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_10 = io_i_partial_products_10[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_10 = io_i_partial_products_10[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_10 = io_i_partial_products_10[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_10 = io_i_partial_products_10[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_10 = io_i_partial_products_10[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_10 = io_i_partial_products_10[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_10 = io_i_partial_products_10[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_10 = io_i_partial_products_10[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_10 = io_i_partial_products_10[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_10 = io_i_partial_products_10[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_10 = io_i_partial_products_10[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_10 = io_i_partial_products_10[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_10 = io_i_partial_products_10[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_10 = io_i_partial_products_10[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_10 = io_i_partial_products_10[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_10 = io_i_partial_products_10[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_10 = io_i_partial_products_10[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_10 = io_i_partial_products_10[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_10 = io_i_partial_products_10[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_10 = io_i_partial_products_10[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_10 = io_i_partial_products_10[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_10 = io_i_partial_products_10[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_10 = io_i_partial_products_10[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_10 = io_i_partial_products_10[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_10 = io_i_partial_products_10[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_10 = io_i_partial_products_10[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_10 = io_i_partial_products_10[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_10 = io_i_partial_products_10[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_10 = io_i_partial_products_10[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_10 = io_i_partial_products_10[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_10 = io_i_partial_products_10[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_10 = io_i_partial_products_10[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_10 = io_i_partial_products_10[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_10 = io_i_partial_products_10[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_10 = io_i_partial_products_10[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_10 = io_i_partial_products_10[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_10 = io_i_partial_products_10[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_10 = io_i_partial_products_10[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_10 = io_i_partial_products_10[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_10 = io_i_partial_products_10[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_10 = io_i_partial_products_10[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_10 = io_i_partial_products_10[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_10 = io_i_partial_products_10[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_10 = io_i_partial_products_10[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_10 = io_i_partial_products_10[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_10 = io_i_partial_products_10[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_10 = io_i_partial_products_10[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_10 = io_i_partial_products_10[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_10 = io_i_partial_products_10[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_10 = io_i_partial_products_10[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_10 = io_i_partial_products_10[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_10 = io_i_partial_products_10[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_10 = io_i_partial_products_10[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_10 = io_i_partial_products_10[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_10 = io_i_partial_products_10[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_10 = io_i_partial_products_10[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_10 = io_i_partial_products_10[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_11 = io_i_partial_products_11[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_11 = io_i_partial_products_11[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_11 = io_i_partial_products_11[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_11 = io_i_partial_products_11[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_11 = io_i_partial_products_11[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_11 = io_i_partial_products_11[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_11 = io_i_partial_products_11[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_11 = io_i_partial_products_11[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_11 = io_i_partial_products_11[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_11 = io_i_partial_products_11[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_11 = io_i_partial_products_11[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_11 = io_i_partial_products_11[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_11 = io_i_partial_products_11[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_11 = io_i_partial_products_11[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_11 = io_i_partial_products_11[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_11 = io_i_partial_products_11[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_11 = io_i_partial_products_11[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_11 = io_i_partial_products_11[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_11 = io_i_partial_products_11[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_11 = io_i_partial_products_11[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_11 = io_i_partial_products_11[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_11 = io_i_partial_products_11[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_11 = io_i_partial_products_11[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_11 = io_i_partial_products_11[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_11 = io_i_partial_products_11[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_11 = io_i_partial_products_11[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_11 = io_i_partial_products_11[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_11 = io_i_partial_products_11[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_11 = io_i_partial_products_11[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_11 = io_i_partial_products_11[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_11 = io_i_partial_products_11[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_11 = io_i_partial_products_11[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_11 = io_i_partial_products_11[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_11 = io_i_partial_products_11[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_11 = io_i_partial_products_11[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_11 = io_i_partial_products_11[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_11 = io_i_partial_products_11[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_11 = io_i_partial_products_11[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_11 = io_i_partial_products_11[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_11 = io_i_partial_products_11[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_11 = io_i_partial_products_11[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_11 = io_i_partial_products_11[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_11 = io_i_partial_products_11[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_11 = io_i_partial_products_11[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_11 = io_i_partial_products_11[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_11 = io_i_partial_products_11[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_11 = io_i_partial_products_11[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_11 = io_i_partial_products_11[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_11 = io_i_partial_products_11[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_11 = io_i_partial_products_11[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_11 = io_i_partial_products_11[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_11 = io_i_partial_products_11[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_11 = io_i_partial_products_11[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_11 = io_i_partial_products_11[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_11 = io_i_partial_products_11[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_11 = io_i_partial_products_11[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_11 = io_i_partial_products_11[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_11 = io_i_partial_products_11[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_11 = io_i_partial_products_11[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_11 = io_i_partial_products_11[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_11 = io_i_partial_products_11[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_11 = io_i_partial_products_11[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_11 = io_i_partial_products_11[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_11 = io_i_partial_products_11[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_11 = io_i_partial_products_11[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_11 = io_i_partial_products_11[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_11 = io_i_partial_products_11[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_11 = io_i_partial_products_11[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_11 = io_i_partial_products_11[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_11 = io_i_partial_products_11[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_11 = io_i_partial_products_11[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_11 = io_i_partial_products_11[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_11 = io_i_partial_products_11[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_11 = io_i_partial_products_11[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_11 = io_i_partial_products_11[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_11 = io_i_partial_products_11[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_11 = io_i_partial_products_11[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_11 = io_i_partial_products_11[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_11 = io_i_partial_products_11[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_11 = io_i_partial_products_11[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_11 = io_i_partial_products_11[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_11 = io_i_partial_products_11[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_11 = io_i_partial_products_11[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_11 = io_i_partial_products_11[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_11 = io_i_partial_products_11[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_11 = io_i_partial_products_11[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_11 = io_i_partial_products_11[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_11 = io_i_partial_products_11[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_11 = io_i_partial_products_11[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_11 = io_i_partial_products_11[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_11 = io_i_partial_products_11[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_11 = io_i_partial_products_11[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_11 = io_i_partial_products_11[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_11 = io_i_partial_products_11[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_11 = io_i_partial_products_11[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_11 = io_i_partial_products_11[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_11 = io_i_partial_products_11[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_11 = io_i_partial_products_11[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_11 = io_i_partial_products_11[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_11 = io_i_partial_products_11[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_11 = io_i_partial_products_11[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_11 = io_i_partial_products_11[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_11 = io_i_partial_products_11[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_11 = io_i_partial_products_11[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_11 = io_i_partial_products_11[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_11 = io_i_partial_products_11[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_11 = io_i_partial_products_11[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_11 = io_i_partial_products_11[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_11 = io_i_partial_products_11[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_11 = io_i_partial_products_11[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_11 = io_i_partial_products_11[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_11 = io_i_partial_products_11[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_11 = io_i_partial_products_11[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_11 = io_i_partial_products_11[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_11 = io_i_partial_products_11[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_11 = io_i_partial_products_11[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_11 = io_i_partial_products_11[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_11 = io_i_partial_products_11[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_11 = io_i_partial_products_11[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_11 = io_i_partial_products_11[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_11 = io_i_partial_products_11[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_11 = io_i_partial_products_11[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_11 = io_i_partial_products_11[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_11 = io_i_partial_products_11[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_11 = io_i_partial_products_11[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_11 = io_i_partial_products_11[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_11 = io_i_partial_products_11[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_11 = io_i_partial_products_11[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_11 = io_i_partial_products_11[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_11 = io_i_partial_products_11[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_11 = io_i_partial_products_11[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_12 = io_i_partial_products_12[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_12 = io_i_partial_products_12[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_12 = io_i_partial_products_12[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_12 = io_i_partial_products_12[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_12 = io_i_partial_products_12[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_12 = io_i_partial_products_12[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_12 = io_i_partial_products_12[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_12 = io_i_partial_products_12[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_12 = io_i_partial_products_12[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_12 = io_i_partial_products_12[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_12 = io_i_partial_products_12[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_12 = io_i_partial_products_12[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_12 = io_i_partial_products_12[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_12 = io_i_partial_products_12[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_12 = io_i_partial_products_12[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_12 = io_i_partial_products_12[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_12 = io_i_partial_products_12[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_12 = io_i_partial_products_12[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_12 = io_i_partial_products_12[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_12 = io_i_partial_products_12[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_12 = io_i_partial_products_12[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_12 = io_i_partial_products_12[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_12 = io_i_partial_products_12[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_12 = io_i_partial_products_12[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_12 = io_i_partial_products_12[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_12 = io_i_partial_products_12[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_12 = io_i_partial_products_12[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_12 = io_i_partial_products_12[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_12 = io_i_partial_products_12[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_12 = io_i_partial_products_12[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_12 = io_i_partial_products_12[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_12 = io_i_partial_products_12[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_12 = io_i_partial_products_12[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_12 = io_i_partial_products_12[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_12 = io_i_partial_products_12[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_12 = io_i_partial_products_12[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_12 = io_i_partial_products_12[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_12 = io_i_partial_products_12[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_12 = io_i_partial_products_12[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_12 = io_i_partial_products_12[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_12 = io_i_partial_products_12[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_12 = io_i_partial_products_12[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_12 = io_i_partial_products_12[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_12 = io_i_partial_products_12[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_12 = io_i_partial_products_12[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_12 = io_i_partial_products_12[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_12 = io_i_partial_products_12[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_12 = io_i_partial_products_12[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_12 = io_i_partial_products_12[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_12 = io_i_partial_products_12[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_12 = io_i_partial_products_12[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_12 = io_i_partial_products_12[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_12 = io_i_partial_products_12[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_12 = io_i_partial_products_12[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_12 = io_i_partial_products_12[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_12 = io_i_partial_products_12[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_12 = io_i_partial_products_12[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_12 = io_i_partial_products_12[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_12 = io_i_partial_products_12[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_12 = io_i_partial_products_12[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_12 = io_i_partial_products_12[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_12 = io_i_partial_products_12[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_12 = io_i_partial_products_12[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_12 = io_i_partial_products_12[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_12 = io_i_partial_products_12[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_12 = io_i_partial_products_12[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_12 = io_i_partial_products_12[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_12 = io_i_partial_products_12[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_12 = io_i_partial_products_12[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_12 = io_i_partial_products_12[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_12 = io_i_partial_products_12[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_12 = io_i_partial_products_12[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_12 = io_i_partial_products_12[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_12 = io_i_partial_products_12[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_12 = io_i_partial_products_12[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_12 = io_i_partial_products_12[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_12 = io_i_partial_products_12[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_12 = io_i_partial_products_12[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_12 = io_i_partial_products_12[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_12 = io_i_partial_products_12[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_12 = io_i_partial_products_12[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_12 = io_i_partial_products_12[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_12 = io_i_partial_products_12[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_12 = io_i_partial_products_12[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_12 = io_i_partial_products_12[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_12 = io_i_partial_products_12[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_12 = io_i_partial_products_12[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_12 = io_i_partial_products_12[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_12 = io_i_partial_products_12[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_12 = io_i_partial_products_12[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_12 = io_i_partial_products_12[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_12 = io_i_partial_products_12[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_12 = io_i_partial_products_12[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_12 = io_i_partial_products_12[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_12 = io_i_partial_products_12[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_12 = io_i_partial_products_12[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_12 = io_i_partial_products_12[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_12 = io_i_partial_products_12[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_12 = io_i_partial_products_12[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_12 = io_i_partial_products_12[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_12 = io_i_partial_products_12[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_12 = io_i_partial_products_12[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_12 = io_i_partial_products_12[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_12 = io_i_partial_products_12[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_12 = io_i_partial_products_12[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_12 = io_i_partial_products_12[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_12 = io_i_partial_products_12[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_12 = io_i_partial_products_12[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_12 = io_i_partial_products_12[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_12 = io_i_partial_products_12[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_12 = io_i_partial_products_12[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_12 = io_i_partial_products_12[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_12 = io_i_partial_products_12[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_12 = io_i_partial_products_12[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_12 = io_i_partial_products_12[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_12 = io_i_partial_products_12[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_12 = io_i_partial_products_12[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_12 = io_i_partial_products_12[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_12 = io_i_partial_products_12[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_12 = io_i_partial_products_12[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_12 = io_i_partial_products_12[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_12 = io_i_partial_products_12[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_12 = io_i_partial_products_12[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_12 = io_i_partial_products_12[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_12 = io_i_partial_products_12[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_12 = io_i_partial_products_12[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_12 = io_i_partial_products_12[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_12 = io_i_partial_products_12[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_12 = io_i_partial_products_12[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_12 = io_i_partial_products_12[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_12 = io_i_partial_products_12[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_13 = io_i_partial_products_13[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_13 = io_i_partial_products_13[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_13 = io_i_partial_products_13[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_13 = io_i_partial_products_13[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_13 = io_i_partial_products_13[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_13 = io_i_partial_products_13[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_13 = io_i_partial_products_13[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_13 = io_i_partial_products_13[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_13 = io_i_partial_products_13[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_13 = io_i_partial_products_13[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_13 = io_i_partial_products_13[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_13 = io_i_partial_products_13[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_13 = io_i_partial_products_13[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_13 = io_i_partial_products_13[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_13 = io_i_partial_products_13[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_13 = io_i_partial_products_13[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_13 = io_i_partial_products_13[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_13 = io_i_partial_products_13[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_13 = io_i_partial_products_13[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_13 = io_i_partial_products_13[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_13 = io_i_partial_products_13[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_13 = io_i_partial_products_13[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_13 = io_i_partial_products_13[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_13 = io_i_partial_products_13[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_13 = io_i_partial_products_13[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_13 = io_i_partial_products_13[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_13 = io_i_partial_products_13[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_13 = io_i_partial_products_13[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_13 = io_i_partial_products_13[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_13 = io_i_partial_products_13[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_13 = io_i_partial_products_13[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_13 = io_i_partial_products_13[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_13 = io_i_partial_products_13[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_13 = io_i_partial_products_13[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_13 = io_i_partial_products_13[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_13 = io_i_partial_products_13[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_13 = io_i_partial_products_13[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_13 = io_i_partial_products_13[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_13 = io_i_partial_products_13[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_13 = io_i_partial_products_13[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_13 = io_i_partial_products_13[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_13 = io_i_partial_products_13[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_13 = io_i_partial_products_13[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_13 = io_i_partial_products_13[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_13 = io_i_partial_products_13[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_13 = io_i_partial_products_13[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_13 = io_i_partial_products_13[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_13 = io_i_partial_products_13[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_13 = io_i_partial_products_13[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_13 = io_i_partial_products_13[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_13 = io_i_partial_products_13[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_13 = io_i_partial_products_13[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_13 = io_i_partial_products_13[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_13 = io_i_partial_products_13[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_13 = io_i_partial_products_13[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_13 = io_i_partial_products_13[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_13 = io_i_partial_products_13[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_13 = io_i_partial_products_13[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_13 = io_i_partial_products_13[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_13 = io_i_partial_products_13[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_13 = io_i_partial_products_13[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_13 = io_i_partial_products_13[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_13 = io_i_partial_products_13[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_13 = io_i_partial_products_13[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_13 = io_i_partial_products_13[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_13 = io_i_partial_products_13[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_13 = io_i_partial_products_13[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_13 = io_i_partial_products_13[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_13 = io_i_partial_products_13[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_13 = io_i_partial_products_13[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_13 = io_i_partial_products_13[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_13 = io_i_partial_products_13[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_13 = io_i_partial_products_13[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_13 = io_i_partial_products_13[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_13 = io_i_partial_products_13[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_13 = io_i_partial_products_13[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_13 = io_i_partial_products_13[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_13 = io_i_partial_products_13[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_13 = io_i_partial_products_13[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_13 = io_i_partial_products_13[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_13 = io_i_partial_products_13[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_13 = io_i_partial_products_13[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_13 = io_i_partial_products_13[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_13 = io_i_partial_products_13[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_13 = io_i_partial_products_13[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_13 = io_i_partial_products_13[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_13 = io_i_partial_products_13[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_13 = io_i_partial_products_13[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_13 = io_i_partial_products_13[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_13 = io_i_partial_products_13[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_13 = io_i_partial_products_13[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_13 = io_i_partial_products_13[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_13 = io_i_partial_products_13[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_13 = io_i_partial_products_13[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_13 = io_i_partial_products_13[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_13 = io_i_partial_products_13[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_13 = io_i_partial_products_13[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_13 = io_i_partial_products_13[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_13 = io_i_partial_products_13[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_13 = io_i_partial_products_13[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_13 = io_i_partial_products_13[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_13 = io_i_partial_products_13[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_13 = io_i_partial_products_13[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_13 = io_i_partial_products_13[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_13 = io_i_partial_products_13[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_13 = io_i_partial_products_13[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_13 = io_i_partial_products_13[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_13 = io_i_partial_products_13[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_13 = io_i_partial_products_13[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_13 = io_i_partial_products_13[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_13 = io_i_partial_products_13[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_13 = io_i_partial_products_13[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_13 = io_i_partial_products_13[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_13 = io_i_partial_products_13[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_13 = io_i_partial_products_13[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_13 = io_i_partial_products_13[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_13 = io_i_partial_products_13[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_13 = io_i_partial_products_13[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_13 = io_i_partial_products_13[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_13 = io_i_partial_products_13[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_13 = io_i_partial_products_13[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_13 = io_i_partial_products_13[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_13 = io_i_partial_products_13[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_13 = io_i_partial_products_13[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_13 = io_i_partial_products_13[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_13 = io_i_partial_products_13[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_13 = io_i_partial_products_13[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_13 = io_i_partial_products_13[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_13 = io_i_partial_products_13[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_13 = io_i_partial_products_13[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_13 = io_i_partial_products_13[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_14 = io_i_partial_products_14[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_14 = io_i_partial_products_14[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_14 = io_i_partial_products_14[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_14 = io_i_partial_products_14[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_14 = io_i_partial_products_14[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_14 = io_i_partial_products_14[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_14 = io_i_partial_products_14[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_14 = io_i_partial_products_14[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_14 = io_i_partial_products_14[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_14 = io_i_partial_products_14[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_14 = io_i_partial_products_14[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_14 = io_i_partial_products_14[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_14 = io_i_partial_products_14[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_14 = io_i_partial_products_14[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_14 = io_i_partial_products_14[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_14 = io_i_partial_products_14[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_14 = io_i_partial_products_14[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_14 = io_i_partial_products_14[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_14 = io_i_partial_products_14[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_14 = io_i_partial_products_14[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_14 = io_i_partial_products_14[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_14 = io_i_partial_products_14[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_14 = io_i_partial_products_14[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_14 = io_i_partial_products_14[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_14 = io_i_partial_products_14[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_14 = io_i_partial_products_14[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_14 = io_i_partial_products_14[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_14 = io_i_partial_products_14[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_14 = io_i_partial_products_14[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_14 = io_i_partial_products_14[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_14 = io_i_partial_products_14[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_14 = io_i_partial_products_14[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_14 = io_i_partial_products_14[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_14 = io_i_partial_products_14[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_14 = io_i_partial_products_14[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_14 = io_i_partial_products_14[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_14 = io_i_partial_products_14[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_14 = io_i_partial_products_14[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_14 = io_i_partial_products_14[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_14 = io_i_partial_products_14[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_14 = io_i_partial_products_14[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_14 = io_i_partial_products_14[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_14 = io_i_partial_products_14[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_14 = io_i_partial_products_14[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_14 = io_i_partial_products_14[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_14 = io_i_partial_products_14[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_14 = io_i_partial_products_14[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_14 = io_i_partial_products_14[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_14 = io_i_partial_products_14[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_14 = io_i_partial_products_14[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_14 = io_i_partial_products_14[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_14 = io_i_partial_products_14[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_14 = io_i_partial_products_14[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_14 = io_i_partial_products_14[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_14 = io_i_partial_products_14[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_14 = io_i_partial_products_14[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_14 = io_i_partial_products_14[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_14 = io_i_partial_products_14[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_14 = io_i_partial_products_14[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_14 = io_i_partial_products_14[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_14 = io_i_partial_products_14[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_14 = io_i_partial_products_14[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_14 = io_i_partial_products_14[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_14 = io_i_partial_products_14[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_14 = io_i_partial_products_14[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_14 = io_i_partial_products_14[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_14 = io_i_partial_products_14[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_14 = io_i_partial_products_14[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_14 = io_i_partial_products_14[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_14 = io_i_partial_products_14[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_14 = io_i_partial_products_14[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_14 = io_i_partial_products_14[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_14 = io_i_partial_products_14[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_14 = io_i_partial_products_14[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_14 = io_i_partial_products_14[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_14 = io_i_partial_products_14[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_14 = io_i_partial_products_14[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_14 = io_i_partial_products_14[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_14 = io_i_partial_products_14[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_14 = io_i_partial_products_14[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_14 = io_i_partial_products_14[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_14 = io_i_partial_products_14[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_14 = io_i_partial_products_14[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_14 = io_i_partial_products_14[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_14 = io_i_partial_products_14[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_14 = io_i_partial_products_14[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_14 = io_i_partial_products_14[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_14 = io_i_partial_products_14[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_14 = io_i_partial_products_14[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_14 = io_i_partial_products_14[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_14 = io_i_partial_products_14[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_14 = io_i_partial_products_14[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_14 = io_i_partial_products_14[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_14 = io_i_partial_products_14[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_14 = io_i_partial_products_14[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_14 = io_i_partial_products_14[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_14 = io_i_partial_products_14[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_14 = io_i_partial_products_14[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_14 = io_i_partial_products_14[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_14 = io_i_partial_products_14[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_14 = io_i_partial_products_14[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_14 = io_i_partial_products_14[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_14 = io_i_partial_products_14[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_14 = io_i_partial_products_14[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_14 = io_i_partial_products_14[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_14 = io_i_partial_products_14[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_14 = io_i_partial_products_14[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_14 = io_i_partial_products_14[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_14 = io_i_partial_products_14[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_14 = io_i_partial_products_14[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_14 = io_i_partial_products_14[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_14 = io_i_partial_products_14[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_14 = io_i_partial_products_14[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_14 = io_i_partial_products_14[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_14 = io_i_partial_products_14[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_14 = io_i_partial_products_14[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_14 = io_i_partial_products_14[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_14 = io_i_partial_products_14[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_14 = io_i_partial_products_14[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_14 = io_i_partial_products_14[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_14 = io_i_partial_products_14[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_14 = io_i_partial_products_14[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_14 = io_i_partial_products_14[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_14 = io_i_partial_products_14[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_14 = io_i_partial_products_14[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_14 = io_i_partial_products_14[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_14 = io_i_partial_products_14[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_14 = io_i_partial_products_14[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_14 = io_i_partial_products_14[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_14 = io_i_partial_products_14[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_14 = io_i_partial_products_14[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_15 = io_i_partial_products_15[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_15 = io_i_partial_products_15[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_15 = io_i_partial_products_15[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_15 = io_i_partial_products_15[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_15 = io_i_partial_products_15[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_15 = io_i_partial_products_15[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_15 = io_i_partial_products_15[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_15 = io_i_partial_products_15[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_15 = io_i_partial_products_15[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_15 = io_i_partial_products_15[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_15 = io_i_partial_products_15[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_15 = io_i_partial_products_15[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_15 = io_i_partial_products_15[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_15 = io_i_partial_products_15[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_15 = io_i_partial_products_15[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_15 = io_i_partial_products_15[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_15 = io_i_partial_products_15[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_15 = io_i_partial_products_15[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_15 = io_i_partial_products_15[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_15 = io_i_partial_products_15[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_15 = io_i_partial_products_15[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_15 = io_i_partial_products_15[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_15 = io_i_partial_products_15[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_15 = io_i_partial_products_15[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_15 = io_i_partial_products_15[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_15 = io_i_partial_products_15[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_15 = io_i_partial_products_15[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_15 = io_i_partial_products_15[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_15 = io_i_partial_products_15[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_15 = io_i_partial_products_15[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_15 = io_i_partial_products_15[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_15 = io_i_partial_products_15[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_15 = io_i_partial_products_15[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_15 = io_i_partial_products_15[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_15 = io_i_partial_products_15[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_15 = io_i_partial_products_15[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_15 = io_i_partial_products_15[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_15 = io_i_partial_products_15[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_15 = io_i_partial_products_15[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_15 = io_i_partial_products_15[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_15 = io_i_partial_products_15[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_15 = io_i_partial_products_15[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_15 = io_i_partial_products_15[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_15 = io_i_partial_products_15[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_15 = io_i_partial_products_15[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_15 = io_i_partial_products_15[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_15 = io_i_partial_products_15[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_15 = io_i_partial_products_15[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_15 = io_i_partial_products_15[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_15 = io_i_partial_products_15[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_15 = io_i_partial_products_15[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_15 = io_i_partial_products_15[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_15 = io_i_partial_products_15[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_15 = io_i_partial_products_15[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_15 = io_i_partial_products_15[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_15 = io_i_partial_products_15[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_15 = io_i_partial_products_15[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_15 = io_i_partial_products_15[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_15 = io_i_partial_products_15[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_15 = io_i_partial_products_15[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_15 = io_i_partial_products_15[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_15 = io_i_partial_products_15[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_15 = io_i_partial_products_15[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_15 = io_i_partial_products_15[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_15 = io_i_partial_products_15[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_15 = io_i_partial_products_15[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_15 = io_i_partial_products_15[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_15 = io_i_partial_products_15[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_15 = io_i_partial_products_15[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_15 = io_i_partial_products_15[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_15 = io_i_partial_products_15[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_15 = io_i_partial_products_15[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_15 = io_i_partial_products_15[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_15 = io_i_partial_products_15[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_15 = io_i_partial_products_15[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_15 = io_i_partial_products_15[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_15 = io_i_partial_products_15[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_15 = io_i_partial_products_15[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_15 = io_i_partial_products_15[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_15 = io_i_partial_products_15[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_15 = io_i_partial_products_15[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_15 = io_i_partial_products_15[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_15 = io_i_partial_products_15[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_15 = io_i_partial_products_15[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_15 = io_i_partial_products_15[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_15 = io_i_partial_products_15[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_15 = io_i_partial_products_15[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_15 = io_i_partial_products_15[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_15 = io_i_partial_products_15[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_15 = io_i_partial_products_15[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_15 = io_i_partial_products_15[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_15 = io_i_partial_products_15[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_15 = io_i_partial_products_15[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_15 = io_i_partial_products_15[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_15 = io_i_partial_products_15[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_15 = io_i_partial_products_15[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_15 = io_i_partial_products_15[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_15 = io_i_partial_products_15[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_15 = io_i_partial_products_15[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_15 = io_i_partial_products_15[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_15 = io_i_partial_products_15[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_15 = io_i_partial_products_15[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_15 = io_i_partial_products_15[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_15 = io_i_partial_products_15[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_15 = io_i_partial_products_15[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_15 = io_i_partial_products_15[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_15 = io_i_partial_products_15[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_15 = io_i_partial_products_15[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_15 = io_i_partial_products_15[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_15 = io_i_partial_products_15[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_15 = io_i_partial_products_15[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_15 = io_i_partial_products_15[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_15 = io_i_partial_products_15[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_15 = io_i_partial_products_15[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_15 = io_i_partial_products_15[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_15 = io_i_partial_products_15[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_15 = io_i_partial_products_15[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_15 = io_i_partial_products_15[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_15 = io_i_partial_products_15[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_15 = io_i_partial_products_15[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_15 = io_i_partial_products_15[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_15 = io_i_partial_products_15[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_15 = io_i_partial_products_15[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_15 = io_i_partial_products_15[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_15 = io_i_partial_products_15[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_15 = io_i_partial_products_15[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_15 = io_i_partial_products_15[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_15 = io_i_partial_products_15[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_15 = io_i_partial_products_15[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_15 = io_i_partial_products_15[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_15 = io_i_partial_products_15[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_16 = io_i_partial_products_16[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_16 = io_i_partial_products_16[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_16 = io_i_partial_products_16[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_16 = io_i_partial_products_16[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_16 = io_i_partial_products_16[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_16 = io_i_partial_products_16[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_16 = io_i_partial_products_16[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_16 = io_i_partial_products_16[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_16 = io_i_partial_products_16[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_16 = io_i_partial_products_16[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_16 = io_i_partial_products_16[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_16 = io_i_partial_products_16[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_16 = io_i_partial_products_16[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_16 = io_i_partial_products_16[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_16 = io_i_partial_products_16[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_16 = io_i_partial_products_16[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_16 = io_i_partial_products_16[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_16 = io_i_partial_products_16[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_16 = io_i_partial_products_16[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_16 = io_i_partial_products_16[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_16 = io_i_partial_products_16[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_16 = io_i_partial_products_16[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_16 = io_i_partial_products_16[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_16 = io_i_partial_products_16[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_16 = io_i_partial_products_16[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_16 = io_i_partial_products_16[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_16 = io_i_partial_products_16[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_16 = io_i_partial_products_16[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_16 = io_i_partial_products_16[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_16 = io_i_partial_products_16[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_16 = io_i_partial_products_16[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_16 = io_i_partial_products_16[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_16 = io_i_partial_products_16[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_16 = io_i_partial_products_16[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_16 = io_i_partial_products_16[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_16 = io_i_partial_products_16[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_16 = io_i_partial_products_16[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_16 = io_i_partial_products_16[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_16 = io_i_partial_products_16[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_16 = io_i_partial_products_16[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_16 = io_i_partial_products_16[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_16 = io_i_partial_products_16[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_16 = io_i_partial_products_16[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_16 = io_i_partial_products_16[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_16 = io_i_partial_products_16[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_16 = io_i_partial_products_16[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_16 = io_i_partial_products_16[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_16 = io_i_partial_products_16[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_16 = io_i_partial_products_16[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_16 = io_i_partial_products_16[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_16 = io_i_partial_products_16[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_16 = io_i_partial_products_16[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_16 = io_i_partial_products_16[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_16 = io_i_partial_products_16[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_16 = io_i_partial_products_16[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_16 = io_i_partial_products_16[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_16 = io_i_partial_products_16[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_16 = io_i_partial_products_16[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_16 = io_i_partial_products_16[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_16 = io_i_partial_products_16[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_16 = io_i_partial_products_16[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_16 = io_i_partial_products_16[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_16 = io_i_partial_products_16[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_16 = io_i_partial_products_16[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_16 = io_i_partial_products_16[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_16 = io_i_partial_products_16[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_16 = io_i_partial_products_16[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_16 = io_i_partial_products_16[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_16 = io_i_partial_products_16[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_16 = io_i_partial_products_16[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_16 = io_i_partial_products_16[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_16 = io_i_partial_products_16[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_16 = io_i_partial_products_16[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_16 = io_i_partial_products_16[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_16 = io_i_partial_products_16[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_16 = io_i_partial_products_16[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_16 = io_i_partial_products_16[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_16 = io_i_partial_products_16[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_16 = io_i_partial_products_16[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_16 = io_i_partial_products_16[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_16 = io_i_partial_products_16[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_16 = io_i_partial_products_16[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_16 = io_i_partial_products_16[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_16 = io_i_partial_products_16[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_16 = io_i_partial_products_16[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_16 = io_i_partial_products_16[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_16 = io_i_partial_products_16[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_16 = io_i_partial_products_16[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_16 = io_i_partial_products_16[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_16 = io_i_partial_products_16[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_16 = io_i_partial_products_16[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_16 = io_i_partial_products_16[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_16 = io_i_partial_products_16[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_16 = io_i_partial_products_16[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_16 = io_i_partial_products_16[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_16 = io_i_partial_products_16[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_16 = io_i_partial_products_16[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_16 = io_i_partial_products_16[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_16 = io_i_partial_products_16[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_16 = io_i_partial_products_16[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_16 = io_i_partial_products_16[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_16 = io_i_partial_products_16[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_16 = io_i_partial_products_16[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_16 = io_i_partial_products_16[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_16 = io_i_partial_products_16[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_16 = io_i_partial_products_16[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_16 = io_i_partial_products_16[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_16 = io_i_partial_products_16[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_16 = io_i_partial_products_16[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_16 = io_i_partial_products_16[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_16 = io_i_partial_products_16[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_16 = io_i_partial_products_16[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_16 = io_i_partial_products_16[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_16 = io_i_partial_products_16[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_16 = io_i_partial_products_16[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_16 = io_i_partial_products_16[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_16 = io_i_partial_products_16[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_16 = io_i_partial_products_16[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_16 = io_i_partial_products_16[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_16 = io_i_partial_products_16[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_16 = io_i_partial_products_16[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_16 = io_i_partial_products_16[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_16 = io_i_partial_products_16[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_16 = io_i_partial_products_16[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_16 = io_i_partial_products_16[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_16 = io_i_partial_products_16[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_16 = io_i_partial_products_16[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_16 = io_i_partial_products_16[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_16 = io_i_partial_products_16[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_16 = io_i_partial_products_16[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_16 = io_i_partial_products_16[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_17 = io_i_partial_products_17[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_17 = io_i_partial_products_17[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_17 = io_i_partial_products_17[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_17 = io_i_partial_products_17[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_17 = io_i_partial_products_17[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_17 = io_i_partial_products_17[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_17 = io_i_partial_products_17[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_17 = io_i_partial_products_17[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_17 = io_i_partial_products_17[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_17 = io_i_partial_products_17[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_17 = io_i_partial_products_17[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_17 = io_i_partial_products_17[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_17 = io_i_partial_products_17[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_17 = io_i_partial_products_17[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_17 = io_i_partial_products_17[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_17 = io_i_partial_products_17[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_17 = io_i_partial_products_17[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_17 = io_i_partial_products_17[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_17 = io_i_partial_products_17[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_17 = io_i_partial_products_17[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_17 = io_i_partial_products_17[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_17 = io_i_partial_products_17[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_17 = io_i_partial_products_17[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_17 = io_i_partial_products_17[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_17 = io_i_partial_products_17[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_17 = io_i_partial_products_17[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_17 = io_i_partial_products_17[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_17 = io_i_partial_products_17[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_17 = io_i_partial_products_17[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_17 = io_i_partial_products_17[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_17 = io_i_partial_products_17[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_17 = io_i_partial_products_17[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_17 = io_i_partial_products_17[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_17 = io_i_partial_products_17[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_17 = io_i_partial_products_17[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_17 = io_i_partial_products_17[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_17 = io_i_partial_products_17[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_17 = io_i_partial_products_17[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_17 = io_i_partial_products_17[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_17 = io_i_partial_products_17[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_17 = io_i_partial_products_17[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_17 = io_i_partial_products_17[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_17 = io_i_partial_products_17[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_17 = io_i_partial_products_17[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_17 = io_i_partial_products_17[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_17 = io_i_partial_products_17[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_17 = io_i_partial_products_17[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_17 = io_i_partial_products_17[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_17 = io_i_partial_products_17[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_17 = io_i_partial_products_17[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_17 = io_i_partial_products_17[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_17 = io_i_partial_products_17[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_17 = io_i_partial_products_17[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_17 = io_i_partial_products_17[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_17 = io_i_partial_products_17[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_17 = io_i_partial_products_17[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_17 = io_i_partial_products_17[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_17 = io_i_partial_products_17[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_17 = io_i_partial_products_17[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_17 = io_i_partial_products_17[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_17 = io_i_partial_products_17[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_17 = io_i_partial_products_17[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_17 = io_i_partial_products_17[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_17 = io_i_partial_products_17[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_17 = io_i_partial_products_17[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_17 = io_i_partial_products_17[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_17 = io_i_partial_products_17[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_17 = io_i_partial_products_17[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_17 = io_i_partial_products_17[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_17 = io_i_partial_products_17[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_17 = io_i_partial_products_17[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_17 = io_i_partial_products_17[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_17 = io_i_partial_products_17[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_17 = io_i_partial_products_17[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_17 = io_i_partial_products_17[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_17 = io_i_partial_products_17[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_17 = io_i_partial_products_17[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_17 = io_i_partial_products_17[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_17 = io_i_partial_products_17[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_17 = io_i_partial_products_17[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_17 = io_i_partial_products_17[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_17 = io_i_partial_products_17[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_17 = io_i_partial_products_17[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_17 = io_i_partial_products_17[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_17 = io_i_partial_products_17[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_17 = io_i_partial_products_17[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_17 = io_i_partial_products_17[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_17 = io_i_partial_products_17[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_17 = io_i_partial_products_17[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_17 = io_i_partial_products_17[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_17 = io_i_partial_products_17[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_17 = io_i_partial_products_17[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_17 = io_i_partial_products_17[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_17 = io_i_partial_products_17[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_17 = io_i_partial_products_17[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_17 = io_i_partial_products_17[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_17 = io_i_partial_products_17[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_17 = io_i_partial_products_17[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_17 = io_i_partial_products_17[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_17 = io_i_partial_products_17[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_17 = io_i_partial_products_17[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_17 = io_i_partial_products_17[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_17 = io_i_partial_products_17[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_17 = io_i_partial_products_17[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_17 = io_i_partial_products_17[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_17 = io_i_partial_products_17[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_17 = io_i_partial_products_17[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_17 = io_i_partial_products_17[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_17 = io_i_partial_products_17[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_17 = io_i_partial_products_17[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_17 = io_i_partial_products_17[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_17 = io_i_partial_products_17[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_17 = io_i_partial_products_17[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_17 = io_i_partial_products_17[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_17 = io_i_partial_products_17[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_17 = io_i_partial_products_17[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_17 = io_i_partial_products_17[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_17 = io_i_partial_products_17[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_17 = io_i_partial_products_17[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_17 = io_i_partial_products_17[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_17 = io_i_partial_products_17[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_17 = io_i_partial_products_17[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_17 = io_i_partial_products_17[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_17 = io_i_partial_products_17[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_17 = io_i_partial_products_17[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_17 = io_i_partial_products_17[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_17 = io_i_partial_products_17[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_17 = io_i_partial_products_17[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_17 = io_i_partial_products_17[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_17 = io_i_partial_products_17[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_17 = io_i_partial_products_17[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_18 = io_i_partial_products_18[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_18 = io_i_partial_products_18[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_18 = io_i_partial_products_18[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_18 = io_i_partial_products_18[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_18 = io_i_partial_products_18[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_18 = io_i_partial_products_18[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_18 = io_i_partial_products_18[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_18 = io_i_partial_products_18[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_18 = io_i_partial_products_18[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_18 = io_i_partial_products_18[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_18 = io_i_partial_products_18[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_18 = io_i_partial_products_18[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_18 = io_i_partial_products_18[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_18 = io_i_partial_products_18[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_18 = io_i_partial_products_18[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_18 = io_i_partial_products_18[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_18 = io_i_partial_products_18[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_18 = io_i_partial_products_18[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_18 = io_i_partial_products_18[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_18 = io_i_partial_products_18[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_18 = io_i_partial_products_18[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_18 = io_i_partial_products_18[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_18 = io_i_partial_products_18[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_18 = io_i_partial_products_18[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_18 = io_i_partial_products_18[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_18 = io_i_partial_products_18[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_18 = io_i_partial_products_18[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_18 = io_i_partial_products_18[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_18 = io_i_partial_products_18[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_18 = io_i_partial_products_18[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_18 = io_i_partial_products_18[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_18 = io_i_partial_products_18[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_18 = io_i_partial_products_18[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_18 = io_i_partial_products_18[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_18 = io_i_partial_products_18[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_18 = io_i_partial_products_18[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_18 = io_i_partial_products_18[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_18 = io_i_partial_products_18[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_18 = io_i_partial_products_18[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_18 = io_i_partial_products_18[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_18 = io_i_partial_products_18[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_18 = io_i_partial_products_18[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_18 = io_i_partial_products_18[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_18 = io_i_partial_products_18[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_18 = io_i_partial_products_18[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_18 = io_i_partial_products_18[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_18 = io_i_partial_products_18[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_18 = io_i_partial_products_18[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_18 = io_i_partial_products_18[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_18 = io_i_partial_products_18[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_18 = io_i_partial_products_18[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_18 = io_i_partial_products_18[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_18 = io_i_partial_products_18[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_18 = io_i_partial_products_18[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_18 = io_i_partial_products_18[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_18 = io_i_partial_products_18[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_18 = io_i_partial_products_18[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_18 = io_i_partial_products_18[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_18 = io_i_partial_products_18[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_18 = io_i_partial_products_18[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_18 = io_i_partial_products_18[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_18 = io_i_partial_products_18[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_18 = io_i_partial_products_18[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_18 = io_i_partial_products_18[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_18 = io_i_partial_products_18[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_18 = io_i_partial_products_18[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_18 = io_i_partial_products_18[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_18 = io_i_partial_products_18[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_18 = io_i_partial_products_18[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_18 = io_i_partial_products_18[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_18 = io_i_partial_products_18[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_18 = io_i_partial_products_18[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_18 = io_i_partial_products_18[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_18 = io_i_partial_products_18[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_18 = io_i_partial_products_18[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_18 = io_i_partial_products_18[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_18 = io_i_partial_products_18[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_18 = io_i_partial_products_18[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_18 = io_i_partial_products_18[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_18 = io_i_partial_products_18[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_18 = io_i_partial_products_18[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_18 = io_i_partial_products_18[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_18 = io_i_partial_products_18[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_18 = io_i_partial_products_18[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_18 = io_i_partial_products_18[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_18 = io_i_partial_products_18[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_18 = io_i_partial_products_18[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_18 = io_i_partial_products_18[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_18 = io_i_partial_products_18[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_18 = io_i_partial_products_18[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_18 = io_i_partial_products_18[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_18 = io_i_partial_products_18[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_18 = io_i_partial_products_18[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_18 = io_i_partial_products_18[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_18 = io_i_partial_products_18[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_18 = io_i_partial_products_18[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_18 = io_i_partial_products_18[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_18 = io_i_partial_products_18[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_18 = io_i_partial_products_18[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_18 = io_i_partial_products_18[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_18 = io_i_partial_products_18[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_18 = io_i_partial_products_18[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_18 = io_i_partial_products_18[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_18 = io_i_partial_products_18[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_18 = io_i_partial_products_18[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_18 = io_i_partial_products_18[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_18 = io_i_partial_products_18[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_18 = io_i_partial_products_18[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_18 = io_i_partial_products_18[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_18 = io_i_partial_products_18[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_18 = io_i_partial_products_18[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_18 = io_i_partial_products_18[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_18 = io_i_partial_products_18[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_18 = io_i_partial_products_18[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_18 = io_i_partial_products_18[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_18 = io_i_partial_products_18[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_18 = io_i_partial_products_18[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_18 = io_i_partial_products_18[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_18 = io_i_partial_products_18[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_18 = io_i_partial_products_18[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_18 = io_i_partial_products_18[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_18 = io_i_partial_products_18[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_18 = io_i_partial_products_18[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_18 = io_i_partial_products_18[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_18 = io_i_partial_products_18[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_18 = io_i_partial_products_18[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_18 = io_i_partial_products_18[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_18 = io_i_partial_products_18[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_18 = io_i_partial_products_18[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_18 = io_i_partial_products_18[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_18 = io_i_partial_products_18[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_19 = io_i_partial_products_19[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_19 = io_i_partial_products_19[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_19 = io_i_partial_products_19[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_19 = io_i_partial_products_19[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_19 = io_i_partial_products_19[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_19 = io_i_partial_products_19[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_19 = io_i_partial_products_19[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_19 = io_i_partial_products_19[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_19 = io_i_partial_products_19[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_19 = io_i_partial_products_19[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_19 = io_i_partial_products_19[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_19 = io_i_partial_products_19[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_19 = io_i_partial_products_19[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_19 = io_i_partial_products_19[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_19 = io_i_partial_products_19[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_19 = io_i_partial_products_19[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_19 = io_i_partial_products_19[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_19 = io_i_partial_products_19[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_19 = io_i_partial_products_19[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_19 = io_i_partial_products_19[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_19 = io_i_partial_products_19[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_19 = io_i_partial_products_19[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_19 = io_i_partial_products_19[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_19 = io_i_partial_products_19[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_19 = io_i_partial_products_19[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_19 = io_i_partial_products_19[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_19 = io_i_partial_products_19[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_19 = io_i_partial_products_19[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_19 = io_i_partial_products_19[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_19 = io_i_partial_products_19[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_19 = io_i_partial_products_19[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_19 = io_i_partial_products_19[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_19 = io_i_partial_products_19[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_19 = io_i_partial_products_19[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_19 = io_i_partial_products_19[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_19 = io_i_partial_products_19[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_19 = io_i_partial_products_19[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_19 = io_i_partial_products_19[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_19 = io_i_partial_products_19[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_19 = io_i_partial_products_19[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_19 = io_i_partial_products_19[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_19 = io_i_partial_products_19[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_19 = io_i_partial_products_19[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_19 = io_i_partial_products_19[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_19 = io_i_partial_products_19[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_19 = io_i_partial_products_19[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_19 = io_i_partial_products_19[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_19 = io_i_partial_products_19[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_19 = io_i_partial_products_19[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_19 = io_i_partial_products_19[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_19 = io_i_partial_products_19[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_19 = io_i_partial_products_19[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_19 = io_i_partial_products_19[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_19 = io_i_partial_products_19[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_19 = io_i_partial_products_19[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_19 = io_i_partial_products_19[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_19 = io_i_partial_products_19[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_19 = io_i_partial_products_19[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_19 = io_i_partial_products_19[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_19 = io_i_partial_products_19[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_19 = io_i_partial_products_19[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_19 = io_i_partial_products_19[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_19 = io_i_partial_products_19[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_19 = io_i_partial_products_19[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_19 = io_i_partial_products_19[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_19 = io_i_partial_products_19[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_19 = io_i_partial_products_19[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_19 = io_i_partial_products_19[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_19 = io_i_partial_products_19[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_19 = io_i_partial_products_19[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_19 = io_i_partial_products_19[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_19 = io_i_partial_products_19[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_19 = io_i_partial_products_19[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_19 = io_i_partial_products_19[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_19 = io_i_partial_products_19[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_19 = io_i_partial_products_19[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_19 = io_i_partial_products_19[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_19 = io_i_partial_products_19[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_19 = io_i_partial_products_19[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_19 = io_i_partial_products_19[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_19 = io_i_partial_products_19[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_19 = io_i_partial_products_19[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_19 = io_i_partial_products_19[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_19 = io_i_partial_products_19[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_19 = io_i_partial_products_19[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_19 = io_i_partial_products_19[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_19 = io_i_partial_products_19[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_19 = io_i_partial_products_19[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_19 = io_i_partial_products_19[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_19 = io_i_partial_products_19[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_19 = io_i_partial_products_19[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_19 = io_i_partial_products_19[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_19 = io_i_partial_products_19[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_19 = io_i_partial_products_19[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_19 = io_i_partial_products_19[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_19 = io_i_partial_products_19[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_19 = io_i_partial_products_19[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_19 = io_i_partial_products_19[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_19 = io_i_partial_products_19[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_19 = io_i_partial_products_19[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_19 = io_i_partial_products_19[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_19 = io_i_partial_products_19[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_19 = io_i_partial_products_19[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_19 = io_i_partial_products_19[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_19 = io_i_partial_products_19[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_19 = io_i_partial_products_19[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_19 = io_i_partial_products_19[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_19 = io_i_partial_products_19[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_19 = io_i_partial_products_19[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_19 = io_i_partial_products_19[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_19 = io_i_partial_products_19[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_19 = io_i_partial_products_19[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_19 = io_i_partial_products_19[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_19 = io_i_partial_products_19[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_19 = io_i_partial_products_19[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_19 = io_i_partial_products_19[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_19 = io_i_partial_products_19[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_19 = io_i_partial_products_19[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_19 = io_i_partial_products_19[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_19 = io_i_partial_products_19[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_19 = io_i_partial_products_19[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_19 = io_i_partial_products_19[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_19 = io_i_partial_products_19[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_19 = io_i_partial_products_19[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_19 = io_i_partial_products_19[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_19 = io_i_partial_products_19[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_19 = io_i_partial_products_19[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_19 = io_i_partial_products_19[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_19 = io_i_partial_products_19[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_19 = io_i_partial_products_19[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_19 = io_i_partial_products_19[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_20 = io_i_partial_products_20[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_20 = io_i_partial_products_20[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_20 = io_i_partial_products_20[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_20 = io_i_partial_products_20[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_20 = io_i_partial_products_20[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_20 = io_i_partial_products_20[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_20 = io_i_partial_products_20[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_20 = io_i_partial_products_20[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_20 = io_i_partial_products_20[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_20 = io_i_partial_products_20[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_20 = io_i_partial_products_20[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_20 = io_i_partial_products_20[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_20 = io_i_partial_products_20[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_20 = io_i_partial_products_20[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_20 = io_i_partial_products_20[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_20 = io_i_partial_products_20[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_20 = io_i_partial_products_20[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_20 = io_i_partial_products_20[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_20 = io_i_partial_products_20[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_20 = io_i_partial_products_20[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_20 = io_i_partial_products_20[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_20 = io_i_partial_products_20[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_20 = io_i_partial_products_20[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_20 = io_i_partial_products_20[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_20 = io_i_partial_products_20[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_20 = io_i_partial_products_20[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_20 = io_i_partial_products_20[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_20 = io_i_partial_products_20[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_20 = io_i_partial_products_20[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_20 = io_i_partial_products_20[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_20 = io_i_partial_products_20[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_20 = io_i_partial_products_20[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_20 = io_i_partial_products_20[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_20 = io_i_partial_products_20[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_20 = io_i_partial_products_20[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_20 = io_i_partial_products_20[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_20 = io_i_partial_products_20[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_20 = io_i_partial_products_20[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_20 = io_i_partial_products_20[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_20 = io_i_partial_products_20[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_20 = io_i_partial_products_20[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_20 = io_i_partial_products_20[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_20 = io_i_partial_products_20[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_20 = io_i_partial_products_20[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_20 = io_i_partial_products_20[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_20 = io_i_partial_products_20[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_20 = io_i_partial_products_20[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_20 = io_i_partial_products_20[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_20 = io_i_partial_products_20[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_20 = io_i_partial_products_20[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_20 = io_i_partial_products_20[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_20 = io_i_partial_products_20[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_20 = io_i_partial_products_20[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_20 = io_i_partial_products_20[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_20 = io_i_partial_products_20[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_20 = io_i_partial_products_20[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_20 = io_i_partial_products_20[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_20 = io_i_partial_products_20[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_20 = io_i_partial_products_20[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_20 = io_i_partial_products_20[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_20 = io_i_partial_products_20[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_20 = io_i_partial_products_20[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_20 = io_i_partial_products_20[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_20 = io_i_partial_products_20[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_20 = io_i_partial_products_20[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_20 = io_i_partial_products_20[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_20 = io_i_partial_products_20[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_20 = io_i_partial_products_20[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_20 = io_i_partial_products_20[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_20 = io_i_partial_products_20[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_20 = io_i_partial_products_20[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_20 = io_i_partial_products_20[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_20 = io_i_partial_products_20[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_20 = io_i_partial_products_20[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_20 = io_i_partial_products_20[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_20 = io_i_partial_products_20[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_20 = io_i_partial_products_20[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_20 = io_i_partial_products_20[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_20 = io_i_partial_products_20[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_20 = io_i_partial_products_20[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_20 = io_i_partial_products_20[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_20 = io_i_partial_products_20[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_20 = io_i_partial_products_20[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_20 = io_i_partial_products_20[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_20 = io_i_partial_products_20[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_20 = io_i_partial_products_20[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_20 = io_i_partial_products_20[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_20 = io_i_partial_products_20[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_20 = io_i_partial_products_20[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_20 = io_i_partial_products_20[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_20 = io_i_partial_products_20[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_20 = io_i_partial_products_20[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_20 = io_i_partial_products_20[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_20 = io_i_partial_products_20[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_20 = io_i_partial_products_20[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_20 = io_i_partial_products_20[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_20 = io_i_partial_products_20[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_20 = io_i_partial_products_20[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_20 = io_i_partial_products_20[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_20 = io_i_partial_products_20[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_20 = io_i_partial_products_20[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_20 = io_i_partial_products_20[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_20 = io_i_partial_products_20[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_20 = io_i_partial_products_20[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_20 = io_i_partial_products_20[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_20 = io_i_partial_products_20[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_20 = io_i_partial_products_20[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_20 = io_i_partial_products_20[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_20 = io_i_partial_products_20[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_20 = io_i_partial_products_20[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_20 = io_i_partial_products_20[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_20 = io_i_partial_products_20[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_20 = io_i_partial_products_20[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_20 = io_i_partial_products_20[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_20 = io_i_partial_products_20[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_20 = io_i_partial_products_20[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_20 = io_i_partial_products_20[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_20 = io_i_partial_products_20[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_20 = io_i_partial_products_20[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_20 = io_i_partial_products_20[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_20 = io_i_partial_products_20[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_20 = io_i_partial_products_20[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_20 = io_i_partial_products_20[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_20 = io_i_partial_products_20[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_20 = io_i_partial_products_20[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_20 = io_i_partial_products_20[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_20 = io_i_partial_products_20[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_20 = io_i_partial_products_20[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_20 = io_i_partial_products_20[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_20 = io_i_partial_products_20[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_20 = io_i_partial_products_20[130]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_0_21 = io_i_partial_products_21[0]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_1_21 = io_i_partial_products_21[1]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_2_21 = io_i_partial_products_21[2]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_3_21 = io_i_partial_products_21[3]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_4_21 = io_i_partial_products_21[4]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_5_21 = io_i_partial_products_21[5]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_6_21 = io_i_partial_products_21[6]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_7_21 = io_i_partial_products_21[7]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_8_21 = io_i_partial_products_21[8]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_9_21 = io_i_partial_products_21[9]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_10_21 = io_i_partial_products_21[10]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_11_21 = io_i_partial_products_21[11]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_12_21 = io_i_partial_products_21[12]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_13_21 = io_i_partial_products_21[13]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_14_21 = io_i_partial_products_21[14]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_15_21 = io_i_partial_products_21[15]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_16_21 = io_i_partial_products_21[16]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_17_21 = io_i_partial_products_21[17]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_18_21 = io_i_partial_products_21[18]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_19_21 = io_i_partial_products_21[19]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_20_21 = io_i_partial_products_21[20]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_21_21 = io_i_partial_products_21[21]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_22_21 = io_i_partial_products_21[22]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_23_21 = io_i_partial_products_21[23]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_24_21 = io_i_partial_products_21[24]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_25_21 = io_i_partial_products_21[25]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_26_21 = io_i_partial_products_21[26]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_27_21 = io_i_partial_products_21[27]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_28_21 = io_i_partial_products_21[28]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_29_21 = io_i_partial_products_21[29]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_30_21 = io_i_partial_products_21[30]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_31_21 = io_i_partial_products_21[31]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_32_21 = io_i_partial_products_21[32]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_33_21 = io_i_partial_products_21[33]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_34_21 = io_i_partial_products_21[34]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_35_21 = io_i_partial_products_21[35]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_36_21 = io_i_partial_products_21[36]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_37_21 = io_i_partial_products_21[37]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_38_21 = io_i_partial_products_21[38]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_39_21 = io_i_partial_products_21[39]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_40_21 = io_i_partial_products_21[40]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_41_21 = io_i_partial_products_21[41]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_42_21 = io_i_partial_products_21[42]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_43_21 = io_i_partial_products_21[43]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_44_21 = io_i_partial_products_21[44]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_45_21 = io_i_partial_products_21[45]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_46_21 = io_i_partial_products_21[46]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_47_21 = io_i_partial_products_21[47]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_48_21 = io_i_partial_products_21[48]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_49_21 = io_i_partial_products_21[49]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_50_21 = io_i_partial_products_21[50]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_51_21 = io_i_partial_products_21[51]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_52_21 = io_i_partial_products_21[52]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_53_21 = io_i_partial_products_21[53]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_54_21 = io_i_partial_products_21[54]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_55_21 = io_i_partial_products_21[55]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_56_21 = io_i_partial_products_21[56]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_57_21 = io_i_partial_products_21[57]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_58_21 = io_i_partial_products_21[58]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_59_21 = io_i_partial_products_21[59]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_60_21 = io_i_partial_products_21[60]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_61_21 = io_i_partial_products_21[61]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_62_21 = io_i_partial_products_21[62]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_63_21 = io_i_partial_products_21[63]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_64_21 = io_i_partial_products_21[64]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_65_21 = io_i_partial_products_21[65]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_66_21 = io_i_partial_products_21[66]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_67_21 = io_i_partial_products_21[67]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_68_21 = io_i_partial_products_21[68]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_69_21 = io_i_partial_products_21[69]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_70_21 = io_i_partial_products_21[70]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_71_21 = io_i_partial_products_21[71]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_72_21 = io_i_partial_products_21[72]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_73_21 = io_i_partial_products_21[73]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_74_21 = io_i_partial_products_21[74]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_75_21 = io_i_partial_products_21[75]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_76_21 = io_i_partial_products_21[76]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_77_21 = io_i_partial_products_21[77]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_78_21 = io_i_partial_products_21[78]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_79_21 = io_i_partial_products_21[79]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_80_21 = io_i_partial_products_21[80]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_81_21 = io_i_partial_products_21[81]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_82_21 = io_i_partial_products_21[82]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_83_21 = io_i_partial_products_21[83]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_84_21 = io_i_partial_products_21[84]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_85_21 = io_i_partial_products_21[85]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_86_21 = io_i_partial_products_21[86]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_87_21 = io_i_partial_products_21[87]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_88_21 = io_i_partial_products_21[88]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_89_21 = io_i_partial_products_21[89]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_90_21 = io_i_partial_products_21[90]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_91_21 = io_i_partial_products_21[91]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_92_21 = io_i_partial_products_21[92]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_93_21 = io_i_partial_products_21[93]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_94_21 = io_i_partial_products_21[94]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_95_21 = io_i_partial_products_21[95]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_96_21 = io_i_partial_products_21[96]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_97_21 = io_i_partial_products_21[97]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_98_21 = io_i_partial_products_21[98]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_99_21 = io_i_partial_products_21[99]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_100_21 = io_i_partial_products_21[100]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_101_21 = io_i_partial_products_21[101]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_102_21 = io_i_partial_products_21[102]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_103_21 = io_i_partial_products_21[103]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_104_21 = io_i_partial_products_21[104]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_105_21 = io_i_partial_products_21[105]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_106_21 = io_i_partial_products_21[106]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_107_21 = io_i_partial_products_21[107]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_108_21 = io_i_partial_products_21[108]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_109_21 = io_i_partial_products_21[109]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_110_21 = io_i_partial_products_21[110]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_111_21 = io_i_partial_products_21[111]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_112_21 = io_i_partial_products_21[112]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_113_21 = io_i_partial_products_21[113]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_114_21 = io_i_partial_products_21[114]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_115_21 = io_i_partial_products_21[115]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_116_21 = io_i_partial_products_21[116]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_117_21 = io_i_partial_products_21[117]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_118_21 = io_i_partial_products_21[118]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_119_21 = io_i_partial_products_21[119]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_120_21 = io_i_partial_products_21[120]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_121_21 = io_i_partial_products_21[121]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_122_21 = io_i_partial_products_21[122]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_123_21 = io_i_partial_products_21[123]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_124_21 = io_i_partial_products_21[124]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_125_21 = io_i_partial_products_21[125]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_126_21 = io_i_partial_products_21[126]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_127_21 = io_i_partial_products_21[127]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_128_21 = io_i_partial_products_21[128]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_129_21 = io_i_partial_products_21[129]; // @[wallace_tree.scala 142:58]
  wire  inversed_pp_130_21 = io_i_partial_products_21[130]; // @[wallace_tree.scala 142:58]
  wire [4:0] wallace_tree_cells_0_io_i_s_lo_lo = {inversed_pp_0_4,inversed_pp_0_3,inversed_pp_0_2,inversed_pp_0_1,
    inversed_pp_0_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_0_io_i_s_lo = {inversed_pp_0_10,inversed_pp_0_9,inversed_pp_0_8,inversed_pp_0_7,
    inversed_pp_0_6,inversed_pp_0_5,wallace_tree_cells_0_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_0_io_i_s_hi_lo = {inversed_pp_0_15,inversed_pp_0_14,inversed_pp_0_13,inversed_pp_0_12,
    inversed_pp_0_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_0_io_i_s_hi = {inversed_pp_0_21,inversed_pp_0_20,inversed_pp_0_19,inversed_pp_0_18,
    inversed_pp_0_17,inversed_pp_0_16,wallace_tree_cells_0_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_1_io_i_s_lo_lo = {inversed_pp_1_4,inversed_pp_1_3,inversed_pp_1_2,inversed_pp_1_1,
    inversed_pp_1_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_1_io_i_s_lo = {inversed_pp_1_10,inversed_pp_1_9,inversed_pp_1_8,inversed_pp_1_7,
    inversed_pp_1_6,inversed_pp_1_5,wallace_tree_cells_1_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_1_io_i_s_hi_lo = {inversed_pp_1_15,inversed_pp_1_14,inversed_pp_1_13,inversed_pp_1_12,
    inversed_pp_1_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_1_io_i_s_hi = {inversed_pp_1_21,inversed_pp_1_20,inversed_pp_1_19,inversed_pp_1_18,
    inversed_pp_1_17,inversed_pp_1_16,wallace_tree_cells_1_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_2_io_i_s_lo_lo = {inversed_pp_2_4,inversed_pp_2_3,inversed_pp_2_2,inversed_pp_2_1,
    inversed_pp_2_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_2_io_i_s_lo = {inversed_pp_2_10,inversed_pp_2_9,inversed_pp_2_8,inversed_pp_2_7,
    inversed_pp_2_6,inversed_pp_2_5,wallace_tree_cells_2_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_2_io_i_s_hi_lo = {inversed_pp_2_15,inversed_pp_2_14,inversed_pp_2_13,inversed_pp_2_12,
    inversed_pp_2_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_2_io_i_s_hi = {inversed_pp_2_21,inversed_pp_2_20,inversed_pp_2_19,inversed_pp_2_18,
    inversed_pp_2_17,inversed_pp_2_16,wallace_tree_cells_2_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_3_io_i_s_lo_lo = {inversed_pp_3_4,inversed_pp_3_3,inversed_pp_3_2,inversed_pp_3_1,
    inversed_pp_3_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_3_io_i_s_lo = {inversed_pp_3_10,inversed_pp_3_9,inversed_pp_3_8,inversed_pp_3_7,
    inversed_pp_3_6,inversed_pp_3_5,wallace_tree_cells_3_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_3_io_i_s_hi_lo = {inversed_pp_3_15,inversed_pp_3_14,inversed_pp_3_13,inversed_pp_3_12,
    inversed_pp_3_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_3_io_i_s_hi = {inversed_pp_3_21,inversed_pp_3_20,inversed_pp_3_19,inversed_pp_3_18,
    inversed_pp_3_17,inversed_pp_3_16,wallace_tree_cells_3_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_4_io_i_s_lo_lo = {inversed_pp_4_4,inversed_pp_4_3,inversed_pp_4_2,inversed_pp_4_1,
    inversed_pp_4_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_4_io_i_s_lo = {inversed_pp_4_10,inversed_pp_4_9,inversed_pp_4_8,inversed_pp_4_7,
    inversed_pp_4_6,inversed_pp_4_5,wallace_tree_cells_4_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_4_io_i_s_hi_lo = {inversed_pp_4_15,inversed_pp_4_14,inversed_pp_4_13,inversed_pp_4_12,
    inversed_pp_4_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_4_io_i_s_hi = {inversed_pp_4_21,inversed_pp_4_20,inversed_pp_4_19,inversed_pp_4_18,
    inversed_pp_4_17,inversed_pp_4_16,wallace_tree_cells_4_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_5_io_i_s_lo_lo = {inversed_pp_5_4,inversed_pp_5_3,inversed_pp_5_2,inversed_pp_5_1,
    inversed_pp_5_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_5_io_i_s_lo = {inversed_pp_5_10,inversed_pp_5_9,inversed_pp_5_8,inversed_pp_5_7,
    inversed_pp_5_6,inversed_pp_5_5,wallace_tree_cells_5_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_5_io_i_s_hi_lo = {inversed_pp_5_15,inversed_pp_5_14,inversed_pp_5_13,inversed_pp_5_12,
    inversed_pp_5_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_5_io_i_s_hi = {inversed_pp_5_21,inversed_pp_5_20,inversed_pp_5_19,inversed_pp_5_18,
    inversed_pp_5_17,inversed_pp_5_16,wallace_tree_cells_5_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_6_io_i_s_lo_lo = {inversed_pp_6_4,inversed_pp_6_3,inversed_pp_6_2,inversed_pp_6_1,
    inversed_pp_6_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_6_io_i_s_lo = {inversed_pp_6_10,inversed_pp_6_9,inversed_pp_6_8,inversed_pp_6_7,
    inversed_pp_6_6,inversed_pp_6_5,wallace_tree_cells_6_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_6_io_i_s_hi_lo = {inversed_pp_6_15,inversed_pp_6_14,inversed_pp_6_13,inversed_pp_6_12,
    inversed_pp_6_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_6_io_i_s_hi = {inversed_pp_6_21,inversed_pp_6_20,inversed_pp_6_19,inversed_pp_6_18,
    inversed_pp_6_17,inversed_pp_6_16,wallace_tree_cells_6_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_7_io_i_s_lo_lo = {inversed_pp_7_4,inversed_pp_7_3,inversed_pp_7_2,inversed_pp_7_1,
    inversed_pp_7_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_7_io_i_s_lo = {inversed_pp_7_10,inversed_pp_7_9,inversed_pp_7_8,inversed_pp_7_7,
    inversed_pp_7_6,inversed_pp_7_5,wallace_tree_cells_7_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_7_io_i_s_hi_lo = {inversed_pp_7_15,inversed_pp_7_14,inversed_pp_7_13,inversed_pp_7_12,
    inversed_pp_7_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_7_io_i_s_hi = {inversed_pp_7_21,inversed_pp_7_20,inversed_pp_7_19,inversed_pp_7_18,
    inversed_pp_7_17,inversed_pp_7_16,wallace_tree_cells_7_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_8_io_i_s_lo_lo = {inversed_pp_8_4,inversed_pp_8_3,inversed_pp_8_2,inversed_pp_8_1,
    inversed_pp_8_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_8_io_i_s_lo = {inversed_pp_8_10,inversed_pp_8_9,inversed_pp_8_8,inversed_pp_8_7,
    inversed_pp_8_6,inversed_pp_8_5,wallace_tree_cells_8_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_8_io_i_s_hi_lo = {inversed_pp_8_15,inversed_pp_8_14,inversed_pp_8_13,inversed_pp_8_12,
    inversed_pp_8_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_8_io_i_s_hi = {inversed_pp_8_21,inversed_pp_8_20,inversed_pp_8_19,inversed_pp_8_18,
    inversed_pp_8_17,inversed_pp_8_16,wallace_tree_cells_8_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_9_io_i_s_lo_lo = {inversed_pp_9_4,inversed_pp_9_3,inversed_pp_9_2,inversed_pp_9_1,
    inversed_pp_9_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_9_io_i_s_lo = {inversed_pp_9_10,inversed_pp_9_9,inversed_pp_9_8,inversed_pp_9_7,
    inversed_pp_9_6,inversed_pp_9_5,wallace_tree_cells_9_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_9_io_i_s_hi_lo = {inversed_pp_9_15,inversed_pp_9_14,inversed_pp_9_13,inversed_pp_9_12,
    inversed_pp_9_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_9_io_i_s_hi = {inversed_pp_9_21,inversed_pp_9_20,inversed_pp_9_19,inversed_pp_9_18,
    inversed_pp_9_17,inversed_pp_9_16,wallace_tree_cells_9_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_10_io_i_s_lo_lo = {inversed_pp_10_4,inversed_pp_10_3,inversed_pp_10_2,inversed_pp_10_1,
    inversed_pp_10_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_10_io_i_s_lo = {inversed_pp_10_10,inversed_pp_10_9,inversed_pp_10_8,inversed_pp_10_7,
    inversed_pp_10_6,inversed_pp_10_5,wallace_tree_cells_10_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_10_io_i_s_hi_lo = {inversed_pp_10_15,inversed_pp_10_14,inversed_pp_10_13,
    inversed_pp_10_12,inversed_pp_10_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_10_io_i_s_hi = {inversed_pp_10_21,inversed_pp_10_20,inversed_pp_10_19,inversed_pp_10_18
    ,inversed_pp_10_17,inversed_pp_10_16,wallace_tree_cells_10_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_11_io_i_s_lo_lo = {inversed_pp_11_4,inversed_pp_11_3,inversed_pp_11_2,inversed_pp_11_1,
    inversed_pp_11_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_11_io_i_s_lo = {inversed_pp_11_10,inversed_pp_11_9,inversed_pp_11_8,inversed_pp_11_7,
    inversed_pp_11_6,inversed_pp_11_5,wallace_tree_cells_11_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_11_io_i_s_hi_lo = {inversed_pp_11_15,inversed_pp_11_14,inversed_pp_11_13,
    inversed_pp_11_12,inversed_pp_11_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_11_io_i_s_hi = {inversed_pp_11_21,inversed_pp_11_20,inversed_pp_11_19,inversed_pp_11_18
    ,inversed_pp_11_17,inversed_pp_11_16,wallace_tree_cells_11_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_12_io_i_s_lo_lo = {inversed_pp_12_4,inversed_pp_12_3,inversed_pp_12_2,inversed_pp_12_1,
    inversed_pp_12_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_12_io_i_s_lo = {inversed_pp_12_10,inversed_pp_12_9,inversed_pp_12_8,inversed_pp_12_7,
    inversed_pp_12_6,inversed_pp_12_5,wallace_tree_cells_12_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_12_io_i_s_hi_lo = {inversed_pp_12_15,inversed_pp_12_14,inversed_pp_12_13,
    inversed_pp_12_12,inversed_pp_12_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_12_io_i_s_hi = {inversed_pp_12_21,inversed_pp_12_20,inversed_pp_12_19,inversed_pp_12_18
    ,inversed_pp_12_17,inversed_pp_12_16,wallace_tree_cells_12_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_13_io_i_s_lo_lo = {inversed_pp_13_4,inversed_pp_13_3,inversed_pp_13_2,inversed_pp_13_1,
    inversed_pp_13_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_13_io_i_s_lo = {inversed_pp_13_10,inversed_pp_13_9,inversed_pp_13_8,inversed_pp_13_7,
    inversed_pp_13_6,inversed_pp_13_5,wallace_tree_cells_13_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_13_io_i_s_hi_lo = {inversed_pp_13_15,inversed_pp_13_14,inversed_pp_13_13,
    inversed_pp_13_12,inversed_pp_13_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_13_io_i_s_hi = {inversed_pp_13_21,inversed_pp_13_20,inversed_pp_13_19,inversed_pp_13_18
    ,inversed_pp_13_17,inversed_pp_13_16,wallace_tree_cells_13_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_14_io_i_s_lo_lo = {inversed_pp_14_4,inversed_pp_14_3,inversed_pp_14_2,inversed_pp_14_1,
    inversed_pp_14_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_14_io_i_s_lo = {inversed_pp_14_10,inversed_pp_14_9,inversed_pp_14_8,inversed_pp_14_7,
    inversed_pp_14_6,inversed_pp_14_5,wallace_tree_cells_14_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_14_io_i_s_hi_lo = {inversed_pp_14_15,inversed_pp_14_14,inversed_pp_14_13,
    inversed_pp_14_12,inversed_pp_14_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_14_io_i_s_hi = {inversed_pp_14_21,inversed_pp_14_20,inversed_pp_14_19,inversed_pp_14_18
    ,inversed_pp_14_17,inversed_pp_14_16,wallace_tree_cells_14_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_15_io_i_s_lo_lo = {inversed_pp_15_4,inversed_pp_15_3,inversed_pp_15_2,inversed_pp_15_1,
    inversed_pp_15_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_15_io_i_s_lo = {inversed_pp_15_10,inversed_pp_15_9,inversed_pp_15_8,inversed_pp_15_7,
    inversed_pp_15_6,inversed_pp_15_5,wallace_tree_cells_15_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_15_io_i_s_hi_lo = {inversed_pp_15_15,inversed_pp_15_14,inversed_pp_15_13,
    inversed_pp_15_12,inversed_pp_15_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_15_io_i_s_hi = {inversed_pp_15_21,inversed_pp_15_20,inversed_pp_15_19,inversed_pp_15_18
    ,inversed_pp_15_17,inversed_pp_15_16,wallace_tree_cells_15_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_16_io_i_s_lo_lo = {inversed_pp_16_4,inversed_pp_16_3,inversed_pp_16_2,inversed_pp_16_1,
    inversed_pp_16_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_16_io_i_s_lo = {inversed_pp_16_10,inversed_pp_16_9,inversed_pp_16_8,inversed_pp_16_7,
    inversed_pp_16_6,inversed_pp_16_5,wallace_tree_cells_16_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_16_io_i_s_hi_lo = {inversed_pp_16_15,inversed_pp_16_14,inversed_pp_16_13,
    inversed_pp_16_12,inversed_pp_16_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_16_io_i_s_hi = {inversed_pp_16_21,inversed_pp_16_20,inversed_pp_16_19,inversed_pp_16_18
    ,inversed_pp_16_17,inversed_pp_16_16,wallace_tree_cells_16_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_17_io_i_s_lo_lo = {inversed_pp_17_4,inversed_pp_17_3,inversed_pp_17_2,inversed_pp_17_1,
    inversed_pp_17_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_17_io_i_s_lo = {inversed_pp_17_10,inversed_pp_17_9,inversed_pp_17_8,inversed_pp_17_7,
    inversed_pp_17_6,inversed_pp_17_5,wallace_tree_cells_17_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_17_io_i_s_hi_lo = {inversed_pp_17_15,inversed_pp_17_14,inversed_pp_17_13,
    inversed_pp_17_12,inversed_pp_17_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_17_io_i_s_hi = {inversed_pp_17_21,inversed_pp_17_20,inversed_pp_17_19,inversed_pp_17_18
    ,inversed_pp_17_17,inversed_pp_17_16,wallace_tree_cells_17_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_18_io_i_s_lo_lo = {inversed_pp_18_4,inversed_pp_18_3,inversed_pp_18_2,inversed_pp_18_1,
    inversed_pp_18_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_18_io_i_s_lo = {inversed_pp_18_10,inversed_pp_18_9,inversed_pp_18_8,inversed_pp_18_7,
    inversed_pp_18_6,inversed_pp_18_5,wallace_tree_cells_18_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_18_io_i_s_hi_lo = {inversed_pp_18_15,inversed_pp_18_14,inversed_pp_18_13,
    inversed_pp_18_12,inversed_pp_18_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_18_io_i_s_hi = {inversed_pp_18_21,inversed_pp_18_20,inversed_pp_18_19,inversed_pp_18_18
    ,inversed_pp_18_17,inversed_pp_18_16,wallace_tree_cells_18_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_19_io_i_s_lo_lo = {inversed_pp_19_4,inversed_pp_19_3,inversed_pp_19_2,inversed_pp_19_1,
    inversed_pp_19_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_19_io_i_s_lo = {inversed_pp_19_10,inversed_pp_19_9,inversed_pp_19_8,inversed_pp_19_7,
    inversed_pp_19_6,inversed_pp_19_5,wallace_tree_cells_19_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_19_io_i_s_hi_lo = {inversed_pp_19_15,inversed_pp_19_14,inversed_pp_19_13,
    inversed_pp_19_12,inversed_pp_19_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_19_io_i_s_hi = {inversed_pp_19_21,inversed_pp_19_20,inversed_pp_19_19,inversed_pp_19_18
    ,inversed_pp_19_17,inversed_pp_19_16,wallace_tree_cells_19_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_20_io_i_s_lo_lo = {inversed_pp_20_4,inversed_pp_20_3,inversed_pp_20_2,inversed_pp_20_1,
    inversed_pp_20_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_20_io_i_s_lo = {inversed_pp_20_10,inversed_pp_20_9,inversed_pp_20_8,inversed_pp_20_7,
    inversed_pp_20_6,inversed_pp_20_5,wallace_tree_cells_20_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_20_io_i_s_hi_lo = {inversed_pp_20_15,inversed_pp_20_14,inversed_pp_20_13,
    inversed_pp_20_12,inversed_pp_20_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_20_io_i_s_hi = {inversed_pp_20_21,inversed_pp_20_20,inversed_pp_20_19,inversed_pp_20_18
    ,inversed_pp_20_17,inversed_pp_20_16,wallace_tree_cells_20_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_21_io_i_s_lo_lo = {inversed_pp_21_4,inversed_pp_21_3,inversed_pp_21_2,inversed_pp_21_1,
    inversed_pp_21_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_21_io_i_s_lo = {inversed_pp_21_10,inversed_pp_21_9,inversed_pp_21_8,inversed_pp_21_7,
    inversed_pp_21_6,inversed_pp_21_5,wallace_tree_cells_21_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_21_io_i_s_hi_lo = {inversed_pp_21_15,inversed_pp_21_14,inversed_pp_21_13,
    inversed_pp_21_12,inversed_pp_21_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_21_io_i_s_hi = {inversed_pp_21_21,inversed_pp_21_20,inversed_pp_21_19,inversed_pp_21_18
    ,inversed_pp_21_17,inversed_pp_21_16,wallace_tree_cells_21_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_22_io_i_s_lo_lo = {inversed_pp_22_4,inversed_pp_22_3,inversed_pp_22_2,inversed_pp_22_1,
    inversed_pp_22_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_22_io_i_s_lo = {inversed_pp_22_10,inversed_pp_22_9,inversed_pp_22_8,inversed_pp_22_7,
    inversed_pp_22_6,inversed_pp_22_5,wallace_tree_cells_22_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_22_io_i_s_hi_lo = {inversed_pp_22_15,inversed_pp_22_14,inversed_pp_22_13,
    inversed_pp_22_12,inversed_pp_22_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_22_io_i_s_hi = {inversed_pp_22_21,inversed_pp_22_20,inversed_pp_22_19,inversed_pp_22_18
    ,inversed_pp_22_17,inversed_pp_22_16,wallace_tree_cells_22_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_23_io_i_s_lo_lo = {inversed_pp_23_4,inversed_pp_23_3,inversed_pp_23_2,inversed_pp_23_1,
    inversed_pp_23_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_23_io_i_s_lo = {inversed_pp_23_10,inversed_pp_23_9,inversed_pp_23_8,inversed_pp_23_7,
    inversed_pp_23_6,inversed_pp_23_5,wallace_tree_cells_23_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_23_io_i_s_hi_lo = {inversed_pp_23_15,inversed_pp_23_14,inversed_pp_23_13,
    inversed_pp_23_12,inversed_pp_23_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_23_io_i_s_hi = {inversed_pp_23_21,inversed_pp_23_20,inversed_pp_23_19,inversed_pp_23_18
    ,inversed_pp_23_17,inversed_pp_23_16,wallace_tree_cells_23_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_24_io_i_s_lo_lo = {inversed_pp_24_4,inversed_pp_24_3,inversed_pp_24_2,inversed_pp_24_1,
    inversed_pp_24_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_24_io_i_s_lo = {inversed_pp_24_10,inversed_pp_24_9,inversed_pp_24_8,inversed_pp_24_7,
    inversed_pp_24_6,inversed_pp_24_5,wallace_tree_cells_24_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_24_io_i_s_hi_lo = {inversed_pp_24_15,inversed_pp_24_14,inversed_pp_24_13,
    inversed_pp_24_12,inversed_pp_24_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_24_io_i_s_hi = {inversed_pp_24_21,inversed_pp_24_20,inversed_pp_24_19,inversed_pp_24_18
    ,inversed_pp_24_17,inversed_pp_24_16,wallace_tree_cells_24_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_25_io_i_s_lo_lo = {inversed_pp_25_4,inversed_pp_25_3,inversed_pp_25_2,inversed_pp_25_1,
    inversed_pp_25_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_25_io_i_s_lo = {inversed_pp_25_10,inversed_pp_25_9,inversed_pp_25_8,inversed_pp_25_7,
    inversed_pp_25_6,inversed_pp_25_5,wallace_tree_cells_25_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_25_io_i_s_hi_lo = {inversed_pp_25_15,inversed_pp_25_14,inversed_pp_25_13,
    inversed_pp_25_12,inversed_pp_25_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_25_io_i_s_hi = {inversed_pp_25_21,inversed_pp_25_20,inversed_pp_25_19,inversed_pp_25_18
    ,inversed_pp_25_17,inversed_pp_25_16,wallace_tree_cells_25_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_26_io_i_s_lo_lo = {inversed_pp_26_4,inversed_pp_26_3,inversed_pp_26_2,inversed_pp_26_1,
    inversed_pp_26_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_26_io_i_s_lo = {inversed_pp_26_10,inversed_pp_26_9,inversed_pp_26_8,inversed_pp_26_7,
    inversed_pp_26_6,inversed_pp_26_5,wallace_tree_cells_26_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_26_io_i_s_hi_lo = {inversed_pp_26_15,inversed_pp_26_14,inversed_pp_26_13,
    inversed_pp_26_12,inversed_pp_26_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_26_io_i_s_hi = {inversed_pp_26_21,inversed_pp_26_20,inversed_pp_26_19,inversed_pp_26_18
    ,inversed_pp_26_17,inversed_pp_26_16,wallace_tree_cells_26_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_27_io_i_s_lo_lo = {inversed_pp_27_4,inversed_pp_27_3,inversed_pp_27_2,inversed_pp_27_1,
    inversed_pp_27_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_27_io_i_s_lo = {inversed_pp_27_10,inversed_pp_27_9,inversed_pp_27_8,inversed_pp_27_7,
    inversed_pp_27_6,inversed_pp_27_5,wallace_tree_cells_27_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_27_io_i_s_hi_lo = {inversed_pp_27_15,inversed_pp_27_14,inversed_pp_27_13,
    inversed_pp_27_12,inversed_pp_27_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_27_io_i_s_hi = {inversed_pp_27_21,inversed_pp_27_20,inversed_pp_27_19,inversed_pp_27_18
    ,inversed_pp_27_17,inversed_pp_27_16,wallace_tree_cells_27_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_28_io_i_s_lo_lo = {inversed_pp_28_4,inversed_pp_28_3,inversed_pp_28_2,inversed_pp_28_1,
    inversed_pp_28_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_28_io_i_s_lo = {inversed_pp_28_10,inversed_pp_28_9,inversed_pp_28_8,inversed_pp_28_7,
    inversed_pp_28_6,inversed_pp_28_5,wallace_tree_cells_28_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_28_io_i_s_hi_lo = {inversed_pp_28_15,inversed_pp_28_14,inversed_pp_28_13,
    inversed_pp_28_12,inversed_pp_28_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_28_io_i_s_hi = {inversed_pp_28_21,inversed_pp_28_20,inversed_pp_28_19,inversed_pp_28_18
    ,inversed_pp_28_17,inversed_pp_28_16,wallace_tree_cells_28_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_29_io_i_s_lo_lo = {inversed_pp_29_4,inversed_pp_29_3,inversed_pp_29_2,inversed_pp_29_1,
    inversed_pp_29_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_29_io_i_s_lo = {inversed_pp_29_10,inversed_pp_29_9,inversed_pp_29_8,inversed_pp_29_7,
    inversed_pp_29_6,inversed_pp_29_5,wallace_tree_cells_29_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_29_io_i_s_hi_lo = {inversed_pp_29_15,inversed_pp_29_14,inversed_pp_29_13,
    inversed_pp_29_12,inversed_pp_29_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_29_io_i_s_hi = {inversed_pp_29_21,inversed_pp_29_20,inversed_pp_29_19,inversed_pp_29_18
    ,inversed_pp_29_17,inversed_pp_29_16,wallace_tree_cells_29_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_30_io_i_s_lo_lo = {inversed_pp_30_4,inversed_pp_30_3,inversed_pp_30_2,inversed_pp_30_1,
    inversed_pp_30_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_30_io_i_s_lo = {inversed_pp_30_10,inversed_pp_30_9,inversed_pp_30_8,inversed_pp_30_7,
    inversed_pp_30_6,inversed_pp_30_5,wallace_tree_cells_30_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_30_io_i_s_hi_lo = {inversed_pp_30_15,inversed_pp_30_14,inversed_pp_30_13,
    inversed_pp_30_12,inversed_pp_30_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_30_io_i_s_hi = {inversed_pp_30_21,inversed_pp_30_20,inversed_pp_30_19,inversed_pp_30_18
    ,inversed_pp_30_17,inversed_pp_30_16,wallace_tree_cells_30_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_31_io_i_s_lo_lo = {inversed_pp_31_4,inversed_pp_31_3,inversed_pp_31_2,inversed_pp_31_1,
    inversed_pp_31_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_31_io_i_s_lo = {inversed_pp_31_10,inversed_pp_31_9,inversed_pp_31_8,inversed_pp_31_7,
    inversed_pp_31_6,inversed_pp_31_5,wallace_tree_cells_31_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_31_io_i_s_hi_lo = {inversed_pp_31_15,inversed_pp_31_14,inversed_pp_31_13,
    inversed_pp_31_12,inversed_pp_31_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_31_io_i_s_hi = {inversed_pp_31_21,inversed_pp_31_20,inversed_pp_31_19,inversed_pp_31_18
    ,inversed_pp_31_17,inversed_pp_31_16,wallace_tree_cells_31_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_32_io_i_s_lo_lo = {inversed_pp_32_4,inversed_pp_32_3,inversed_pp_32_2,inversed_pp_32_1,
    inversed_pp_32_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_32_io_i_s_lo = {inversed_pp_32_10,inversed_pp_32_9,inversed_pp_32_8,inversed_pp_32_7,
    inversed_pp_32_6,inversed_pp_32_5,wallace_tree_cells_32_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_32_io_i_s_hi_lo = {inversed_pp_32_15,inversed_pp_32_14,inversed_pp_32_13,
    inversed_pp_32_12,inversed_pp_32_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_32_io_i_s_hi = {inversed_pp_32_21,inversed_pp_32_20,inversed_pp_32_19,inversed_pp_32_18
    ,inversed_pp_32_17,inversed_pp_32_16,wallace_tree_cells_32_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_33_io_i_s_lo_lo = {inversed_pp_33_4,inversed_pp_33_3,inversed_pp_33_2,inversed_pp_33_1,
    inversed_pp_33_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_33_io_i_s_lo = {inversed_pp_33_10,inversed_pp_33_9,inversed_pp_33_8,inversed_pp_33_7,
    inversed_pp_33_6,inversed_pp_33_5,wallace_tree_cells_33_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_33_io_i_s_hi_lo = {inversed_pp_33_15,inversed_pp_33_14,inversed_pp_33_13,
    inversed_pp_33_12,inversed_pp_33_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_33_io_i_s_hi = {inversed_pp_33_21,inversed_pp_33_20,inversed_pp_33_19,inversed_pp_33_18
    ,inversed_pp_33_17,inversed_pp_33_16,wallace_tree_cells_33_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_34_io_i_s_lo_lo = {inversed_pp_34_4,inversed_pp_34_3,inversed_pp_34_2,inversed_pp_34_1,
    inversed_pp_34_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_34_io_i_s_lo = {inversed_pp_34_10,inversed_pp_34_9,inversed_pp_34_8,inversed_pp_34_7,
    inversed_pp_34_6,inversed_pp_34_5,wallace_tree_cells_34_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_34_io_i_s_hi_lo = {inversed_pp_34_15,inversed_pp_34_14,inversed_pp_34_13,
    inversed_pp_34_12,inversed_pp_34_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_34_io_i_s_hi = {inversed_pp_34_21,inversed_pp_34_20,inversed_pp_34_19,inversed_pp_34_18
    ,inversed_pp_34_17,inversed_pp_34_16,wallace_tree_cells_34_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_35_io_i_s_lo_lo = {inversed_pp_35_4,inversed_pp_35_3,inversed_pp_35_2,inversed_pp_35_1,
    inversed_pp_35_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_35_io_i_s_lo = {inversed_pp_35_10,inversed_pp_35_9,inversed_pp_35_8,inversed_pp_35_7,
    inversed_pp_35_6,inversed_pp_35_5,wallace_tree_cells_35_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_35_io_i_s_hi_lo = {inversed_pp_35_15,inversed_pp_35_14,inversed_pp_35_13,
    inversed_pp_35_12,inversed_pp_35_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_35_io_i_s_hi = {inversed_pp_35_21,inversed_pp_35_20,inversed_pp_35_19,inversed_pp_35_18
    ,inversed_pp_35_17,inversed_pp_35_16,wallace_tree_cells_35_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_36_io_i_s_lo_lo = {inversed_pp_36_4,inversed_pp_36_3,inversed_pp_36_2,inversed_pp_36_1,
    inversed_pp_36_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_36_io_i_s_lo = {inversed_pp_36_10,inversed_pp_36_9,inversed_pp_36_8,inversed_pp_36_7,
    inversed_pp_36_6,inversed_pp_36_5,wallace_tree_cells_36_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_36_io_i_s_hi_lo = {inversed_pp_36_15,inversed_pp_36_14,inversed_pp_36_13,
    inversed_pp_36_12,inversed_pp_36_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_36_io_i_s_hi = {inversed_pp_36_21,inversed_pp_36_20,inversed_pp_36_19,inversed_pp_36_18
    ,inversed_pp_36_17,inversed_pp_36_16,wallace_tree_cells_36_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_37_io_i_s_lo_lo = {inversed_pp_37_4,inversed_pp_37_3,inversed_pp_37_2,inversed_pp_37_1,
    inversed_pp_37_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_37_io_i_s_lo = {inversed_pp_37_10,inversed_pp_37_9,inversed_pp_37_8,inversed_pp_37_7,
    inversed_pp_37_6,inversed_pp_37_5,wallace_tree_cells_37_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_37_io_i_s_hi_lo = {inversed_pp_37_15,inversed_pp_37_14,inversed_pp_37_13,
    inversed_pp_37_12,inversed_pp_37_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_37_io_i_s_hi = {inversed_pp_37_21,inversed_pp_37_20,inversed_pp_37_19,inversed_pp_37_18
    ,inversed_pp_37_17,inversed_pp_37_16,wallace_tree_cells_37_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_38_io_i_s_lo_lo = {inversed_pp_38_4,inversed_pp_38_3,inversed_pp_38_2,inversed_pp_38_1,
    inversed_pp_38_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_38_io_i_s_lo = {inversed_pp_38_10,inversed_pp_38_9,inversed_pp_38_8,inversed_pp_38_7,
    inversed_pp_38_6,inversed_pp_38_5,wallace_tree_cells_38_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_38_io_i_s_hi_lo = {inversed_pp_38_15,inversed_pp_38_14,inversed_pp_38_13,
    inversed_pp_38_12,inversed_pp_38_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_38_io_i_s_hi = {inversed_pp_38_21,inversed_pp_38_20,inversed_pp_38_19,inversed_pp_38_18
    ,inversed_pp_38_17,inversed_pp_38_16,wallace_tree_cells_38_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_39_io_i_s_lo_lo = {inversed_pp_39_4,inversed_pp_39_3,inversed_pp_39_2,inversed_pp_39_1,
    inversed_pp_39_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_39_io_i_s_lo = {inversed_pp_39_10,inversed_pp_39_9,inversed_pp_39_8,inversed_pp_39_7,
    inversed_pp_39_6,inversed_pp_39_5,wallace_tree_cells_39_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_39_io_i_s_hi_lo = {inversed_pp_39_15,inversed_pp_39_14,inversed_pp_39_13,
    inversed_pp_39_12,inversed_pp_39_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_39_io_i_s_hi = {inversed_pp_39_21,inversed_pp_39_20,inversed_pp_39_19,inversed_pp_39_18
    ,inversed_pp_39_17,inversed_pp_39_16,wallace_tree_cells_39_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_40_io_i_s_lo_lo = {inversed_pp_40_4,inversed_pp_40_3,inversed_pp_40_2,inversed_pp_40_1,
    inversed_pp_40_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_40_io_i_s_lo = {inversed_pp_40_10,inversed_pp_40_9,inversed_pp_40_8,inversed_pp_40_7,
    inversed_pp_40_6,inversed_pp_40_5,wallace_tree_cells_40_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_40_io_i_s_hi_lo = {inversed_pp_40_15,inversed_pp_40_14,inversed_pp_40_13,
    inversed_pp_40_12,inversed_pp_40_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_40_io_i_s_hi = {inversed_pp_40_21,inversed_pp_40_20,inversed_pp_40_19,inversed_pp_40_18
    ,inversed_pp_40_17,inversed_pp_40_16,wallace_tree_cells_40_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_41_io_i_s_lo_lo = {inversed_pp_41_4,inversed_pp_41_3,inversed_pp_41_2,inversed_pp_41_1,
    inversed_pp_41_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_41_io_i_s_lo = {inversed_pp_41_10,inversed_pp_41_9,inversed_pp_41_8,inversed_pp_41_7,
    inversed_pp_41_6,inversed_pp_41_5,wallace_tree_cells_41_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_41_io_i_s_hi_lo = {inversed_pp_41_15,inversed_pp_41_14,inversed_pp_41_13,
    inversed_pp_41_12,inversed_pp_41_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_41_io_i_s_hi = {inversed_pp_41_21,inversed_pp_41_20,inversed_pp_41_19,inversed_pp_41_18
    ,inversed_pp_41_17,inversed_pp_41_16,wallace_tree_cells_41_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_42_io_i_s_lo_lo = {inversed_pp_42_4,inversed_pp_42_3,inversed_pp_42_2,inversed_pp_42_1,
    inversed_pp_42_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_42_io_i_s_lo = {inversed_pp_42_10,inversed_pp_42_9,inversed_pp_42_8,inversed_pp_42_7,
    inversed_pp_42_6,inversed_pp_42_5,wallace_tree_cells_42_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_42_io_i_s_hi_lo = {inversed_pp_42_15,inversed_pp_42_14,inversed_pp_42_13,
    inversed_pp_42_12,inversed_pp_42_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_42_io_i_s_hi = {inversed_pp_42_21,inversed_pp_42_20,inversed_pp_42_19,inversed_pp_42_18
    ,inversed_pp_42_17,inversed_pp_42_16,wallace_tree_cells_42_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_43_io_i_s_lo_lo = {inversed_pp_43_4,inversed_pp_43_3,inversed_pp_43_2,inversed_pp_43_1,
    inversed_pp_43_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_43_io_i_s_lo = {inversed_pp_43_10,inversed_pp_43_9,inversed_pp_43_8,inversed_pp_43_7,
    inversed_pp_43_6,inversed_pp_43_5,wallace_tree_cells_43_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_43_io_i_s_hi_lo = {inversed_pp_43_15,inversed_pp_43_14,inversed_pp_43_13,
    inversed_pp_43_12,inversed_pp_43_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_43_io_i_s_hi = {inversed_pp_43_21,inversed_pp_43_20,inversed_pp_43_19,inversed_pp_43_18
    ,inversed_pp_43_17,inversed_pp_43_16,wallace_tree_cells_43_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_44_io_i_s_lo_lo = {inversed_pp_44_4,inversed_pp_44_3,inversed_pp_44_2,inversed_pp_44_1,
    inversed_pp_44_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_44_io_i_s_lo = {inversed_pp_44_10,inversed_pp_44_9,inversed_pp_44_8,inversed_pp_44_7,
    inversed_pp_44_6,inversed_pp_44_5,wallace_tree_cells_44_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_44_io_i_s_hi_lo = {inversed_pp_44_15,inversed_pp_44_14,inversed_pp_44_13,
    inversed_pp_44_12,inversed_pp_44_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_44_io_i_s_hi = {inversed_pp_44_21,inversed_pp_44_20,inversed_pp_44_19,inversed_pp_44_18
    ,inversed_pp_44_17,inversed_pp_44_16,wallace_tree_cells_44_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_45_io_i_s_lo_lo = {inversed_pp_45_4,inversed_pp_45_3,inversed_pp_45_2,inversed_pp_45_1,
    inversed_pp_45_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_45_io_i_s_lo = {inversed_pp_45_10,inversed_pp_45_9,inversed_pp_45_8,inversed_pp_45_7,
    inversed_pp_45_6,inversed_pp_45_5,wallace_tree_cells_45_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_45_io_i_s_hi_lo = {inversed_pp_45_15,inversed_pp_45_14,inversed_pp_45_13,
    inversed_pp_45_12,inversed_pp_45_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_45_io_i_s_hi = {inversed_pp_45_21,inversed_pp_45_20,inversed_pp_45_19,inversed_pp_45_18
    ,inversed_pp_45_17,inversed_pp_45_16,wallace_tree_cells_45_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_46_io_i_s_lo_lo = {inversed_pp_46_4,inversed_pp_46_3,inversed_pp_46_2,inversed_pp_46_1,
    inversed_pp_46_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_46_io_i_s_lo = {inversed_pp_46_10,inversed_pp_46_9,inversed_pp_46_8,inversed_pp_46_7,
    inversed_pp_46_6,inversed_pp_46_5,wallace_tree_cells_46_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_46_io_i_s_hi_lo = {inversed_pp_46_15,inversed_pp_46_14,inversed_pp_46_13,
    inversed_pp_46_12,inversed_pp_46_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_46_io_i_s_hi = {inversed_pp_46_21,inversed_pp_46_20,inversed_pp_46_19,inversed_pp_46_18
    ,inversed_pp_46_17,inversed_pp_46_16,wallace_tree_cells_46_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_47_io_i_s_lo_lo = {inversed_pp_47_4,inversed_pp_47_3,inversed_pp_47_2,inversed_pp_47_1,
    inversed_pp_47_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_47_io_i_s_lo = {inversed_pp_47_10,inversed_pp_47_9,inversed_pp_47_8,inversed_pp_47_7,
    inversed_pp_47_6,inversed_pp_47_5,wallace_tree_cells_47_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_47_io_i_s_hi_lo = {inversed_pp_47_15,inversed_pp_47_14,inversed_pp_47_13,
    inversed_pp_47_12,inversed_pp_47_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_47_io_i_s_hi = {inversed_pp_47_21,inversed_pp_47_20,inversed_pp_47_19,inversed_pp_47_18
    ,inversed_pp_47_17,inversed_pp_47_16,wallace_tree_cells_47_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_48_io_i_s_lo_lo = {inversed_pp_48_4,inversed_pp_48_3,inversed_pp_48_2,inversed_pp_48_1,
    inversed_pp_48_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_48_io_i_s_lo = {inversed_pp_48_10,inversed_pp_48_9,inversed_pp_48_8,inversed_pp_48_7,
    inversed_pp_48_6,inversed_pp_48_5,wallace_tree_cells_48_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_48_io_i_s_hi_lo = {inversed_pp_48_15,inversed_pp_48_14,inversed_pp_48_13,
    inversed_pp_48_12,inversed_pp_48_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_48_io_i_s_hi = {inversed_pp_48_21,inversed_pp_48_20,inversed_pp_48_19,inversed_pp_48_18
    ,inversed_pp_48_17,inversed_pp_48_16,wallace_tree_cells_48_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_49_io_i_s_lo_lo = {inversed_pp_49_4,inversed_pp_49_3,inversed_pp_49_2,inversed_pp_49_1,
    inversed_pp_49_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_49_io_i_s_lo = {inversed_pp_49_10,inversed_pp_49_9,inversed_pp_49_8,inversed_pp_49_7,
    inversed_pp_49_6,inversed_pp_49_5,wallace_tree_cells_49_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_49_io_i_s_hi_lo = {inversed_pp_49_15,inversed_pp_49_14,inversed_pp_49_13,
    inversed_pp_49_12,inversed_pp_49_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_49_io_i_s_hi = {inversed_pp_49_21,inversed_pp_49_20,inversed_pp_49_19,inversed_pp_49_18
    ,inversed_pp_49_17,inversed_pp_49_16,wallace_tree_cells_49_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_50_io_i_s_lo_lo = {inversed_pp_50_4,inversed_pp_50_3,inversed_pp_50_2,inversed_pp_50_1,
    inversed_pp_50_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_50_io_i_s_lo = {inversed_pp_50_10,inversed_pp_50_9,inversed_pp_50_8,inversed_pp_50_7,
    inversed_pp_50_6,inversed_pp_50_5,wallace_tree_cells_50_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_50_io_i_s_hi_lo = {inversed_pp_50_15,inversed_pp_50_14,inversed_pp_50_13,
    inversed_pp_50_12,inversed_pp_50_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_50_io_i_s_hi = {inversed_pp_50_21,inversed_pp_50_20,inversed_pp_50_19,inversed_pp_50_18
    ,inversed_pp_50_17,inversed_pp_50_16,wallace_tree_cells_50_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_51_io_i_s_lo_lo = {inversed_pp_51_4,inversed_pp_51_3,inversed_pp_51_2,inversed_pp_51_1,
    inversed_pp_51_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_51_io_i_s_lo = {inversed_pp_51_10,inversed_pp_51_9,inversed_pp_51_8,inversed_pp_51_7,
    inversed_pp_51_6,inversed_pp_51_5,wallace_tree_cells_51_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_51_io_i_s_hi_lo = {inversed_pp_51_15,inversed_pp_51_14,inversed_pp_51_13,
    inversed_pp_51_12,inversed_pp_51_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_51_io_i_s_hi = {inversed_pp_51_21,inversed_pp_51_20,inversed_pp_51_19,inversed_pp_51_18
    ,inversed_pp_51_17,inversed_pp_51_16,wallace_tree_cells_51_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_52_io_i_s_lo_lo = {inversed_pp_52_4,inversed_pp_52_3,inversed_pp_52_2,inversed_pp_52_1,
    inversed_pp_52_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_52_io_i_s_lo = {inversed_pp_52_10,inversed_pp_52_9,inversed_pp_52_8,inversed_pp_52_7,
    inversed_pp_52_6,inversed_pp_52_5,wallace_tree_cells_52_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_52_io_i_s_hi_lo = {inversed_pp_52_15,inversed_pp_52_14,inversed_pp_52_13,
    inversed_pp_52_12,inversed_pp_52_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_52_io_i_s_hi = {inversed_pp_52_21,inversed_pp_52_20,inversed_pp_52_19,inversed_pp_52_18
    ,inversed_pp_52_17,inversed_pp_52_16,wallace_tree_cells_52_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_53_io_i_s_lo_lo = {inversed_pp_53_4,inversed_pp_53_3,inversed_pp_53_2,inversed_pp_53_1,
    inversed_pp_53_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_53_io_i_s_lo = {inversed_pp_53_10,inversed_pp_53_9,inversed_pp_53_8,inversed_pp_53_7,
    inversed_pp_53_6,inversed_pp_53_5,wallace_tree_cells_53_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_53_io_i_s_hi_lo = {inversed_pp_53_15,inversed_pp_53_14,inversed_pp_53_13,
    inversed_pp_53_12,inversed_pp_53_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_53_io_i_s_hi = {inversed_pp_53_21,inversed_pp_53_20,inversed_pp_53_19,inversed_pp_53_18
    ,inversed_pp_53_17,inversed_pp_53_16,wallace_tree_cells_53_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_54_io_i_s_lo_lo = {inversed_pp_54_4,inversed_pp_54_3,inversed_pp_54_2,inversed_pp_54_1,
    inversed_pp_54_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_54_io_i_s_lo = {inversed_pp_54_10,inversed_pp_54_9,inversed_pp_54_8,inversed_pp_54_7,
    inversed_pp_54_6,inversed_pp_54_5,wallace_tree_cells_54_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_54_io_i_s_hi_lo = {inversed_pp_54_15,inversed_pp_54_14,inversed_pp_54_13,
    inversed_pp_54_12,inversed_pp_54_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_54_io_i_s_hi = {inversed_pp_54_21,inversed_pp_54_20,inversed_pp_54_19,inversed_pp_54_18
    ,inversed_pp_54_17,inversed_pp_54_16,wallace_tree_cells_54_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_55_io_i_s_lo_lo = {inversed_pp_55_4,inversed_pp_55_3,inversed_pp_55_2,inversed_pp_55_1,
    inversed_pp_55_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_55_io_i_s_lo = {inversed_pp_55_10,inversed_pp_55_9,inversed_pp_55_8,inversed_pp_55_7,
    inversed_pp_55_6,inversed_pp_55_5,wallace_tree_cells_55_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_55_io_i_s_hi_lo = {inversed_pp_55_15,inversed_pp_55_14,inversed_pp_55_13,
    inversed_pp_55_12,inversed_pp_55_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_55_io_i_s_hi = {inversed_pp_55_21,inversed_pp_55_20,inversed_pp_55_19,inversed_pp_55_18
    ,inversed_pp_55_17,inversed_pp_55_16,wallace_tree_cells_55_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_56_io_i_s_lo_lo = {inversed_pp_56_4,inversed_pp_56_3,inversed_pp_56_2,inversed_pp_56_1,
    inversed_pp_56_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_56_io_i_s_lo = {inversed_pp_56_10,inversed_pp_56_9,inversed_pp_56_8,inversed_pp_56_7,
    inversed_pp_56_6,inversed_pp_56_5,wallace_tree_cells_56_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_56_io_i_s_hi_lo = {inversed_pp_56_15,inversed_pp_56_14,inversed_pp_56_13,
    inversed_pp_56_12,inversed_pp_56_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_56_io_i_s_hi = {inversed_pp_56_21,inversed_pp_56_20,inversed_pp_56_19,inversed_pp_56_18
    ,inversed_pp_56_17,inversed_pp_56_16,wallace_tree_cells_56_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_57_io_i_s_lo_lo = {inversed_pp_57_4,inversed_pp_57_3,inversed_pp_57_2,inversed_pp_57_1,
    inversed_pp_57_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_57_io_i_s_lo = {inversed_pp_57_10,inversed_pp_57_9,inversed_pp_57_8,inversed_pp_57_7,
    inversed_pp_57_6,inversed_pp_57_5,wallace_tree_cells_57_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_57_io_i_s_hi_lo = {inversed_pp_57_15,inversed_pp_57_14,inversed_pp_57_13,
    inversed_pp_57_12,inversed_pp_57_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_57_io_i_s_hi = {inversed_pp_57_21,inversed_pp_57_20,inversed_pp_57_19,inversed_pp_57_18
    ,inversed_pp_57_17,inversed_pp_57_16,wallace_tree_cells_57_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_58_io_i_s_lo_lo = {inversed_pp_58_4,inversed_pp_58_3,inversed_pp_58_2,inversed_pp_58_1,
    inversed_pp_58_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_58_io_i_s_lo = {inversed_pp_58_10,inversed_pp_58_9,inversed_pp_58_8,inversed_pp_58_7,
    inversed_pp_58_6,inversed_pp_58_5,wallace_tree_cells_58_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_58_io_i_s_hi_lo = {inversed_pp_58_15,inversed_pp_58_14,inversed_pp_58_13,
    inversed_pp_58_12,inversed_pp_58_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_58_io_i_s_hi = {inversed_pp_58_21,inversed_pp_58_20,inversed_pp_58_19,inversed_pp_58_18
    ,inversed_pp_58_17,inversed_pp_58_16,wallace_tree_cells_58_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_59_io_i_s_lo_lo = {inversed_pp_59_4,inversed_pp_59_3,inversed_pp_59_2,inversed_pp_59_1,
    inversed_pp_59_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_59_io_i_s_lo = {inversed_pp_59_10,inversed_pp_59_9,inversed_pp_59_8,inversed_pp_59_7,
    inversed_pp_59_6,inversed_pp_59_5,wallace_tree_cells_59_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_59_io_i_s_hi_lo = {inversed_pp_59_15,inversed_pp_59_14,inversed_pp_59_13,
    inversed_pp_59_12,inversed_pp_59_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_59_io_i_s_hi = {inversed_pp_59_21,inversed_pp_59_20,inversed_pp_59_19,inversed_pp_59_18
    ,inversed_pp_59_17,inversed_pp_59_16,wallace_tree_cells_59_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_60_io_i_s_lo_lo = {inversed_pp_60_4,inversed_pp_60_3,inversed_pp_60_2,inversed_pp_60_1,
    inversed_pp_60_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_60_io_i_s_lo = {inversed_pp_60_10,inversed_pp_60_9,inversed_pp_60_8,inversed_pp_60_7,
    inversed_pp_60_6,inversed_pp_60_5,wallace_tree_cells_60_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_60_io_i_s_hi_lo = {inversed_pp_60_15,inversed_pp_60_14,inversed_pp_60_13,
    inversed_pp_60_12,inversed_pp_60_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_60_io_i_s_hi = {inversed_pp_60_21,inversed_pp_60_20,inversed_pp_60_19,inversed_pp_60_18
    ,inversed_pp_60_17,inversed_pp_60_16,wallace_tree_cells_60_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_61_io_i_s_lo_lo = {inversed_pp_61_4,inversed_pp_61_3,inversed_pp_61_2,inversed_pp_61_1,
    inversed_pp_61_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_61_io_i_s_lo = {inversed_pp_61_10,inversed_pp_61_9,inversed_pp_61_8,inversed_pp_61_7,
    inversed_pp_61_6,inversed_pp_61_5,wallace_tree_cells_61_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_61_io_i_s_hi_lo = {inversed_pp_61_15,inversed_pp_61_14,inversed_pp_61_13,
    inversed_pp_61_12,inversed_pp_61_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_61_io_i_s_hi = {inversed_pp_61_21,inversed_pp_61_20,inversed_pp_61_19,inversed_pp_61_18
    ,inversed_pp_61_17,inversed_pp_61_16,wallace_tree_cells_61_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_62_io_i_s_lo_lo = {inversed_pp_62_4,inversed_pp_62_3,inversed_pp_62_2,inversed_pp_62_1,
    inversed_pp_62_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_62_io_i_s_lo = {inversed_pp_62_10,inversed_pp_62_9,inversed_pp_62_8,inversed_pp_62_7,
    inversed_pp_62_6,inversed_pp_62_5,wallace_tree_cells_62_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_62_io_i_s_hi_lo = {inversed_pp_62_15,inversed_pp_62_14,inversed_pp_62_13,
    inversed_pp_62_12,inversed_pp_62_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_62_io_i_s_hi = {inversed_pp_62_21,inversed_pp_62_20,inversed_pp_62_19,inversed_pp_62_18
    ,inversed_pp_62_17,inversed_pp_62_16,wallace_tree_cells_62_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_63_io_i_s_lo_lo = {inversed_pp_63_4,inversed_pp_63_3,inversed_pp_63_2,inversed_pp_63_1,
    inversed_pp_63_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_63_io_i_s_lo = {inversed_pp_63_10,inversed_pp_63_9,inversed_pp_63_8,inversed_pp_63_7,
    inversed_pp_63_6,inversed_pp_63_5,wallace_tree_cells_63_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_63_io_i_s_hi_lo = {inversed_pp_63_15,inversed_pp_63_14,inversed_pp_63_13,
    inversed_pp_63_12,inversed_pp_63_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_63_io_i_s_hi = {inversed_pp_63_21,inversed_pp_63_20,inversed_pp_63_19,inversed_pp_63_18
    ,inversed_pp_63_17,inversed_pp_63_16,wallace_tree_cells_63_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_64_io_i_s_lo_lo = {inversed_pp_64_4,inversed_pp_64_3,inversed_pp_64_2,inversed_pp_64_1,
    inversed_pp_64_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_64_io_i_s_lo = {inversed_pp_64_10,inversed_pp_64_9,inversed_pp_64_8,inversed_pp_64_7,
    inversed_pp_64_6,inversed_pp_64_5,wallace_tree_cells_64_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_64_io_i_s_hi_lo = {inversed_pp_64_15,inversed_pp_64_14,inversed_pp_64_13,
    inversed_pp_64_12,inversed_pp_64_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_64_io_i_s_hi = {inversed_pp_64_21,inversed_pp_64_20,inversed_pp_64_19,inversed_pp_64_18
    ,inversed_pp_64_17,inversed_pp_64_16,wallace_tree_cells_64_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_65_io_i_s_lo_lo = {inversed_pp_65_4,inversed_pp_65_3,inversed_pp_65_2,inversed_pp_65_1,
    inversed_pp_65_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_65_io_i_s_lo = {inversed_pp_65_10,inversed_pp_65_9,inversed_pp_65_8,inversed_pp_65_7,
    inversed_pp_65_6,inversed_pp_65_5,wallace_tree_cells_65_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_65_io_i_s_hi_lo = {inversed_pp_65_15,inversed_pp_65_14,inversed_pp_65_13,
    inversed_pp_65_12,inversed_pp_65_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_65_io_i_s_hi = {inversed_pp_65_21,inversed_pp_65_20,inversed_pp_65_19,inversed_pp_65_18
    ,inversed_pp_65_17,inversed_pp_65_16,wallace_tree_cells_65_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_66_io_i_s_lo_lo = {inversed_pp_66_4,inversed_pp_66_3,inversed_pp_66_2,inversed_pp_66_1,
    inversed_pp_66_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_66_io_i_s_lo = {inversed_pp_66_10,inversed_pp_66_9,inversed_pp_66_8,inversed_pp_66_7,
    inversed_pp_66_6,inversed_pp_66_5,wallace_tree_cells_66_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_66_io_i_s_hi_lo = {inversed_pp_66_15,inversed_pp_66_14,inversed_pp_66_13,
    inversed_pp_66_12,inversed_pp_66_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_66_io_i_s_hi = {inversed_pp_66_21,inversed_pp_66_20,inversed_pp_66_19,inversed_pp_66_18
    ,inversed_pp_66_17,inversed_pp_66_16,wallace_tree_cells_66_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_67_io_i_s_lo_lo = {inversed_pp_67_4,inversed_pp_67_3,inversed_pp_67_2,inversed_pp_67_1,
    inversed_pp_67_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_67_io_i_s_lo = {inversed_pp_67_10,inversed_pp_67_9,inversed_pp_67_8,inversed_pp_67_7,
    inversed_pp_67_6,inversed_pp_67_5,wallace_tree_cells_67_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_67_io_i_s_hi_lo = {inversed_pp_67_15,inversed_pp_67_14,inversed_pp_67_13,
    inversed_pp_67_12,inversed_pp_67_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_67_io_i_s_hi = {inversed_pp_67_21,inversed_pp_67_20,inversed_pp_67_19,inversed_pp_67_18
    ,inversed_pp_67_17,inversed_pp_67_16,wallace_tree_cells_67_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_68_io_i_s_lo_lo = {inversed_pp_68_4,inversed_pp_68_3,inversed_pp_68_2,inversed_pp_68_1,
    inversed_pp_68_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_68_io_i_s_lo = {inversed_pp_68_10,inversed_pp_68_9,inversed_pp_68_8,inversed_pp_68_7,
    inversed_pp_68_6,inversed_pp_68_5,wallace_tree_cells_68_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_68_io_i_s_hi_lo = {inversed_pp_68_15,inversed_pp_68_14,inversed_pp_68_13,
    inversed_pp_68_12,inversed_pp_68_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_68_io_i_s_hi = {inversed_pp_68_21,inversed_pp_68_20,inversed_pp_68_19,inversed_pp_68_18
    ,inversed_pp_68_17,inversed_pp_68_16,wallace_tree_cells_68_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_69_io_i_s_lo_lo = {inversed_pp_69_4,inversed_pp_69_3,inversed_pp_69_2,inversed_pp_69_1,
    inversed_pp_69_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_69_io_i_s_lo = {inversed_pp_69_10,inversed_pp_69_9,inversed_pp_69_8,inversed_pp_69_7,
    inversed_pp_69_6,inversed_pp_69_5,wallace_tree_cells_69_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_69_io_i_s_hi_lo = {inversed_pp_69_15,inversed_pp_69_14,inversed_pp_69_13,
    inversed_pp_69_12,inversed_pp_69_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_69_io_i_s_hi = {inversed_pp_69_21,inversed_pp_69_20,inversed_pp_69_19,inversed_pp_69_18
    ,inversed_pp_69_17,inversed_pp_69_16,wallace_tree_cells_69_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_70_io_i_s_lo_lo = {inversed_pp_70_4,inversed_pp_70_3,inversed_pp_70_2,inversed_pp_70_1,
    inversed_pp_70_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_70_io_i_s_lo = {inversed_pp_70_10,inversed_pp_70_9,inversed_pp_70_8,inversed_pp_70_7,
    inversed_pp_70_6,inversed_pp_70_5,wallace_tree_cells_70_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_70_io_i_s_hi_lo = {inversed_pp_70_15,inversed_pp_70_14,inversed_pp_70_13,
    inversed_pp_70_12,inversed_pp_70_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_70_io_i_s_hi = {inversed_pp_70_21,inversed_pp_70_20,inversed_pp_70_19,inversed_pp_70_18
    ,inversed_pp_70_17,inversed_pp_70_16,wallace_tree_cells_70_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_71_io_i_s_lo_lo = {inversed_pp_71_4,inversed_pp_71_3,inversed_pp_71_2,inversed_pp_71_1,
    inversed_pp_71_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_71_io_i_s_lo = {inversed_pp_71_10,inversed_pp_71_9,inversed_pp_71_8,inversed_pp_71_7,
    inversed_pp_71_6,inversed_pp_71_5,wallace_tree_cells_71_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_71_io_i_s_hi_lo = {inversed_pp_71_15,inversed_pp_71_14,inversed_pp_71_13,
    inversed_pp_71_12,inversed_pp_71_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_71_io_i_s_hi = {inversed_pp_71_21,inversed_pp_71_20,inversed_pp_71_19,inversed_pp_71_18
    ,inversed_pp_71_17,inversed_pp_71_16,wallace_tree_cells_71_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_72_io_i_s_lo_lo = {inversed_pp_72_4,inversed_pp_72_3,inversed_pp_72_2,inversed_pp_72_1,
    inversed_pp_72_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_72_io_i_s_lo = {inversed_pp_72_10,inversed_pp_72_9,inversed_pp_72_8,inversed_pp_72_7,
    inversed_pp_72_6,inversed_pp_72_5,wallace_tree_cells_72_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_72_io_i_s_hi_lo = {inversed_pp_72_15,inversed_pp_72_14,inversed_pp_72_13,
    inversed_pp_72_12,inversed_pp_72_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_72_io_i_s_hi = {inversed_pp_72_21,inversed_pp_72_20,inversed_pp_72_19,inversed_pp_72_18
    ,inversed_pp_72_17,inversed_pp_72_16,wallace_tree_cells_72_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_73_io_i_s_lo_lo = {inversed_pp_73_4,inversed_pp_73_3,inversed_pp_73_2,inversed_pp_73_1,
    inversed_pp_73_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_73_io_i_s_lo = {inversed_pp_73_10,inversed_pp_73_9,inversed_pp_73_8,inversed_pp_73_7,
    inversed_pp_73_6,inversed_pp_73_5,wallace_tree_cells_73_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_73_io_i_s_hi_lo = {inversed_pp_73_15,inversed_pp_73_14,inversed_pp_73_13,
    inversed_pp_73_12,inversed_pp_73_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_73_io_i_s_hi = {inversed_pp_73_21,inversed_pp_73_20,inversed_pp_73_19,inversed_pp_73_18
    ,inversed_pp_73_17,inversed_pp_73_16,wallace_tree_cells_73_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_74_io_i_s_lo_lo = {inversed_pp_74_4,inversed_pp_74_3,inversed_pp_74_2,inversed_pp_74_1,
    inversed_pp_74_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_74_io_i_s_lo = {inversed_pp_74_10,inversed_pp_74_9,inversed_pp_74_8,inversed_pp_74_7,
    inversed_pp_74_6,inversed_pp_74_5,wallace_tree_cells_74_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_74_io_i_s_hi_lo = {inversed_pp_74_15,inversed_pp_74_14,inversed_pp_74_13,
    inversed_pp_74_12,inversed_pp_74_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_74_io_i_s_hi = {inversed_pp_74_21,inversed_pp_74_20,inversed_pp_74_19,inversed_pp_74_18
    ,inversed_pp_74_17,inversed_pp_74_16,wallace_tree_cells_74_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_75_io_i_s_lo_lo = {inversed_pp_75_4,inversed_pp_75_3,inversed_pp_75_2,inversed_pp_75_1,
    inversed_pp_75_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_75_io_i_s_lo = {inversed_pp_75_10,inversed_pp_75_9,inversed_pp_75_8,inversed_pp_75_7,
    inversed_pp_75_6,inversed_pp_75_5,wallace_tree_cells_75_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_75_io_i_s_hi_lo = {inversed_pp_75_15,inversed_pp_75_14,inversed_pp_75_13,
    inversed_pp_75_12,inversed_pp_75_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_75_io_i_s_hi = {inversed_pp_75_21,inversed_pp_75_20,inversed_pp_75_19,inversed_pp_75_18
    ,inversed_pp_75_17,inversed_pp_75_16,wallace_tree_cells_75_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_76_io_i_s_lo_lo = {inversed_pp_76_4,inversed_pp_76_3,inversed_pp_76_2,inversed_pp_76_1,
    inversed_pp_76_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_76_io_i_s_lo = {inversed_pp_76_10,inversed_pp_76_9,inversed_pp_76_8,inversed_pp_76_7,
    inversed_pp_76_6,inversed_pp_76_5,wallace_tree_cells_76_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_76_io_i_s_hi_lo = {inversed_pp_76_15,inversed_pp_76_14,inversed_pp_76_13,
    inversed_pp_76_12,inversed_pp_76_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_76_io_i_s_hi = {inversed_pp_76_21,inversed_pp_76_20,inversed_pp_76_19,inversed_pp_76_18
    ,inversed_pp_76_17,inversed_pp_76_16,wallace_tree_cells_76_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_77_io_i_s_lo_lo = {inversed_pp_77_4,inversed_pp_77_3,inversed_pp_77_2,inversed_pp_77_1,
    inversed_pp_77_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_77_io_i_s_lo = {inversed_pp_77_10,inversed_pp_77_9,inversed_pp_77_8,inversed_pp_77_7,
    inversed_pp_77_6,inversed_pp_77_5,wallace_tree_cells_77_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_77_io_i_s_hi_lo = {inversed_pp_77_15,inversed_pp_77_14,inversed_pp_77_13,
    inversed_pp_77_12,inversed_pp_77_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_77_io_i_s_hi = {inversed_pp_77_21,inversed_pp_77_20,inversed_pp_77_19,inversed_pp_77_18
    ,inversed_pp_77_17,inversed_pp_77_16,wallace_tree_cells_77_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_78_io_i_s_lo_lo = {inversed_pp_78_4,inversed_pp_78_3,inversed_pp_78_2,inversed_pp_78_1,
    inversed_pp_78_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_78_io_i_s_lo = {inversed_pp_78_10,inversed_pp_78_9,inversed_pp_78_8,inversed_pp_78_7,
    inversed_pp_78_6,inversed_pp_78_5,wallace_tree_cells_78_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_78_io_i_s_hi_lo = {inversed_pp_78_15,inversed_pp_78_14,inversed_pp_78_13,
    inversed_pp_78_12,inversed_pp_78_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_78_io_i_s_hi = {inversed_pp_78_21,inversed_pp_78_20,inversed_pp_78_19,inversed_pp_78_18
    ,inversed_pp_78_17,inversed_pp_78_16,wallace_tree_cells_78_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_79_io_i_s_lo_lo = {inversed_pp_79_4,inversed_pp_79_3,inversed_pp_79_2,inversed_pp_79_1,
    inversed_pp_79_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_79_io_i_s_lo = {inversed_pp_79_10,inversed_pp_79_9,inversed_pp_79_8,inversed_pp_79_7,
    inversed_pp_79_6,inversed_pp_79_5,wallace_tree_cells_79_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_79_io_i_s_hi_lo = {inversed_pp_79_15,inversed_pp_79_14,inversed_pp_79_13,
    inversed_pp_79_12,inversed_pp_79_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_79_io_i_s_hi = {inversed_pp_79_21,inversed_pp_79_20,inversed_pp_79_19,inversed_pp_79_18
    ,inversed_pp_79_17,inversed_pp_79_16,wallace_tree_cells_79_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_80_io_i_s_lo_lo = {inversed_pp_80_4,inversed_pp_80_3,inversed_pp_80_2,inversed_pp_80_1,
    inversed_pp_80_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_80_io_i_s_lo = {inversed_pp_80_10,inversed_pp_80_9,inversed_pp_80_8,inversed_pp_80_7,
    inversed_pp_80_6,inversed_pp_80_5,wallace_tree_cells_80_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_80_io_i_s_hi_lo = {inversed_pp_80_15,inversed_pp_80_14,inversed_pp_80_13,
    inversed_pp_80_12,inversed_pp_80_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_80_io_i_s_hi = {inversed_pp_80_21,inversed_pp_80_20,inversed_pp_80_19,inversed_pp_80_18
    ,inversed_pp_80_17,inversed_pp_80_16,wallace_tree_cells_80_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_81_io_i_s_lo_lo = {inversed_pp_81_4,inversed_pp_81_3,inversed_pp_81_2,inversed_pp_81_1,
    inversed_pp_81_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_81_io_i_s_lo = {inversed_pp_81_10,inversed_pp_81_9,inversed_pp_81_8,inversed_pp_81_7,
    inversed_pp_81_6,inversed_pp_81_5,wallace_tree_cells_81_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_81_io_i_s_hi_lo = {inversed_pp_81_15,inversed_pp_81_14,inversed_pp_81_13,
    inversed_pp_81_12,inversed_pp_81_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_81_io_i_s_hi = {inversed_pp_81_21,inversed_pp_81_20,inversed_pp_81_19,inversed_pp_81_18
    ,inversed_pp_81_17,inversed_pp_81_16,wallace_tree_cells_81_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_82_io_i_s_lo_lo = {inversed_pp_82_4,inversed_pp_82_3,inversed_pp_82_2,inversed_pp_82_1,
    inversed_pp_82_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_82_io_i_s_lo = {inversed_pp_82_10,inversed_pp_82_9,inversed_pp_82_8,inversed_pp_82_7,
    inversed_pp_82_6,inversed_pp_82_5,wallace_tree_cells_82_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_82_io_i_s_hi_lo = {inversed_pp_82_15,inversed_pp_82_14,inversed_pp_82_13,
    inversed_pp_82_12,inversed_pp_82_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_82_io_i_s_hi = {inversed_pp_82_21,inversed_pp_82_20,inversed_pp_82_19,inversed_pp_82_18
    ,inversed_pp_82_17,inversed_pp_82_16,wallace_tree_cells_82_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_83_io_i_s_lo_lo = {inversed_pp_83_4,inversed_pp_83_3,inversed_pp_83_2,inversed_pp_83_1,
    inversed_pp_83_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_83_io_i_s_lo = {inversed_pp_83_10,inversed_pp_83_9,inversed_pp_83_8,inversed_pp_83_7,
    inversed_pp_83_6,inversed_pp_83_5,wallace_tree_cells_83_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_83_io_i_s_hi_lo = {inversed_pp_83_15,inversed_pp_83_14,inversed_pp_83_13,
    inversed_pp_83_12,inversed_pp_83_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_83_io_i_s_hi = {inversed_pp_83_21,inversed_pp_83_20,inversed_pp_83_19,inversed_pp_83_18
    ,inversed_pp_83_17,inversed_pp_83_16,wallace_tree_cells_83_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_84_io_i_s_lo_lo = {inversed_pp_84_4,inversed_pp_84_3,inversed_pp_84_2,inversed_pp_84_1,
    inversed_pp_84_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_84_io_i_s_lo = {inversed_pp_84_10,inversed_pp_84_9,inversed_pp_84_8,inversed_pp_84_7,
    inversed_pp_84_6,inversed_pp_84_5,wallace_tree_cells_84_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_84_io_i_s_hi_lo = {inversed_pp_84_15,inversed_pp_84_14,inversed_pp_84_13,
    inversed_pp_84_12,inversed_pp_84_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_84_io_i_s_hi = {inversed_pp_84_21,inversed_pp_84_20,inversed_pp_84_19,inversed_pp_84_18
    ,inversed_pp_84_17,inversed_pp_84_16,wallace_tree_cells_84_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_85_io_i_s_lo_lo = {inversed_pp_85_4,inversed_pp_85_3,inversed_pp_85_2,inversed_pp_85_1,
    inversed_pp_85_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_85_io_i_s_lo = {inversed_pp_85_10,inversed_pp_85_9,inversed_pp_85_8,inversed_pp_85_7,
    inversed_pp_85_6,inversed_pp_85_5,wallace_tree_cells_85_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_85_io_i_s_hi_lo = {inversed_pp_85_15,inversed_pp_85_14,inversed_pp_85_13,
    inversed_pp_85_12,inversed_pp_85_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_85_io_i_s_hi = {inversed_pp_85_21,inversed_pp_85_20,inversed_pp_85_19,inversed_pp_85_18
    ,inversed_pp_85_17,inversed_pp_85_16,wallace_tree_cells_85_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_86_io_i_s_lo_lo = {inversed_pp_86_4,inversed_pp_86_3,inversed_pp_86_2,inversed_pp_86_1,
    inversed_pp_86_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_86_io_i_s_lo = {inversed_pp_86_10,inversed_pp_86_9,inversed_pp_86_8,inversed_pp_86_7,
    inversed_pp_86_6,inversed_pp_86_5,wallace_tree_cells_86_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_86_io_i_s_hi_lo = {inversed_pp_86_15,inversed_pp_86_14,inversed_pp_86_13,
    inversed_pp_86_12,inversed_pp_86_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_86_io_i_s_hi = {inversed_pp_86_21,inversed_pp_86_20,inversed_pp_86_19,inversed_pp_86_18
    ,inversed_pp_86_17,inversed_pp_86_16,wallace_tree_cells_86_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_87_io_i_s_lo_lo = {inversed_pp_87_4,inversed_pp_87_3,inversed_pp_87_2,inversed_pp_87_1,
    inversed_pp_87_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_87_io_i_s_lo = {inversed_pp_87_10,inversed_pp_87_9,inversed_pp_87_8,inversed_pp_87_7,
    inversed_pp_87_6,inversed_pp_87_5,wallace_tree_cells_87_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_87_io_i_s_hi_lo = {inversed_pp_87_15,inversed_pp_87_14,inversed_pp_87_13,
    inversed_pp_87_12,inversed_pp_87_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_87_io_i_s_hi = {inversed_pp_87_21,inversed_pp_87_20,inversed_pp_87_19,inversed_pp_87_18
    ,inversed_pp_87_17,inversed_pp_87_16,wallace_tree_cells_87_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_88_io_i_s_lo_lo = {inversed_pp_88_4,inversed_pp_88_3,inversed_pp_88_2,inversed_pp_88_1,
    inversed_pp_88_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_88_io_i_s_lo = {inversed_pp_88_10,inversed_pp_88_9,inversed_pp_88_8,inversed_pp_88_7,
    inversed_pp_88_6,inversed_pp_88_5,wallace_tree_cells_88_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_88_io_i_s_hi_lo = {inversed_pp_88_15,inversed_pp_88_14,inversed_pp_88_13,
    inversed_pp_88_12,inversed_pp_88_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_88_io_i_s_hi = {inversed_pp_88_21,inversed_pp_88_20,inversed_pp_88_19,inversed_pp_88_18
    ,inversed_pp_88_17,inversed_pp_88_16,wallace_tree_cells_88_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_89_io_i_s_lo_lo = {inversed_pp_89_4,inversed_pp_89_3,inversed_pp_89_2,inversed_pp_89_1,
    inversed_pp_89_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_89_io_i_s_lo = {inversed_pp_89_10,inversed_pp_89_9,inversed_pp_89_8,inversed_pp_89_7,
    inversed_pp_89_6,inversed_pp_89_5,wallace_tree_cells_89_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_89_io_i_s_hi_lo = {inversed_pp_89_15,inversed_pp_89_14,inversed_pp_89_13,
    inversed_pp_89_12,inversed_pp_89_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_89_io_i_s_hi = {inversed_pp_89_21,inversed_pp_89_20,inversed_pp_89_19,inversed_pp_89_18
    ,inversed_pp_89_17,inversed_pp_89_16,wallace_tree_cells_89_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_90_io_i_s_lo_lo = {inversed_pp_90_4,inversed_pp_90_3,inversed_pp_90_2,inversed_pp_90_1,
    inversed_pp_90_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_90_io_i_s_lo = {inversed_pp_90_10,inversed_pp_90_9,inversed_pp_90_8,inversed_pp_90_7,
    inversed_pp_90_6,inversed_pp_90_5,wallace_tree_cells_90_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_90_io_i_s_hi_lo = {inversed_pp_90_15,inversed_pp_90_14,inversed_pp_90_13,
    inversed_pp_90_12,inversed_pp_90_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_90_io_i_s_hi = {inversed_pp_90_21,inversed_pp_90_20,inversed_pp_90_19,inversed_pp_90_18
    ,inversed_pp_90_17,inversed_pp_90_16,wallace_tree_cells_90_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_91_io_i_s_lo_lo = {inversed_pp_91_4,inversed_pp_91_3,inversed_pp_91_2,inversed_pp_91_1,
    inversed_pp_91_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_91_io_i_s_lo = {inversed_pp_91_10,inversed_pp_91_9,inversed_pp_91_8,inversed_pp_91_7,
    inversed_pp_91_6,inversed_pp_91_5,wallace_tree_cells_91_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_91_io_i_s_hi_lo = {inversed_pp_91_15,inversed_pp_91_14,inversed_pp_91_13,
    inversed_pp_91_12,inversed_pp_91_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_91_io_i_s_hi = {inversed_pp_91_21,inversed_pp_91_20,inversed_pp_91_19,inversed_pp_91_18
    ,inversed_pp_91_17,inversed_pp_91_16,wallace_tree_cells_91_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_92_io_i_s_lo_lo = {inversed_pp_92_4,inversed_pp_92_3,inversed_pp_92_2,inversed_pp_92_1,
    inversed_pp_92_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_92_io_i_s_lo = {inversed_pp_92_10,inversed_pp_92_9,inversed_pp_92_8,inversed_pp_92_7,
    inversed_pp_92_6,inversed_pp_92_5,wallace_tree_cells_92_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_92_io_i_s_hi_lo = {inversed_pp_92_15,inversed_pp_92_14,inversed_pp_92_13,
    inversed_pp_92_12,inversed_pp_92_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_92_io_i_s_hi = {inversed_pp_92_21,inversed_pp_92_20,inversed_pp_92_19,inversed_pp_92_18
    ,inversed_pp_92_17,inversed_pp_92_16,wallace_tree_cells_92_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_93_io_i_s_lo_lo = {inversed_pp_93_4,inversed_pp_93_3,inversed_pp_93_2,inversed_pp_93_1,
    inversed_pp_93_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_93_io_i_s_lo = {inversed_pp_93_10,inversed_pp_93_9,inversed_pp_93_8,inversed_pp_93_7,
    inversed_pp_93_6,inversed_pp_93_5,wallace_tree_cells_93_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_93_io_i_s_hi_lo = {inversed_pp_93_15,inversed_pp_93_14,inversed_pp_93_13,
    inversed_pp_93_12,inversed_pp_93_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_93_io_i_s_hi = {inversed_pp_93_21,inversed_pp_93_20,inversed_pp_93_19,inversed_pp_93_18
    ,inversed_pp_93_17,inversed_pp_93_16,wallace_tree_cells_93_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_94_io_i_s_lo_lo = {inversed_pp_94_4,inversed_pp_94_3,inversed_pp_94_2,inversed_pp_94_1,
    inversed_pp_94_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_94_io_i_s_lo = {inversed_pp_94_10,inversed_pp_94_9,inversed_pp_94_8,inversed_pp_94_7,
    inversed_pp_94_6,inversed_pp_94_5,wallace_tree_cells_94_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_94_io_i_s_hi_lo = {inversed_pp_94_15,inversed_pp_94_14,inversed_pp_94_13,
    inversed_pp_94_12,inversed_pp_94_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_94_io_i_s_hi = {inversed_pp_94_21,inversed_pp_94_20,inversed_pp_94_19,inversed_pp_94_18
    ,inversed_pp_94_17,inversed_pp_94_16,wallace_tree_cells_94_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_95_io_i_s_lo_lo = {inversed_pp_95_4,inversed_pp_95_3,inversed_pp_95_2,inversed_pp_95_1,
    inversed_pp_95_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_95_io_i_s_lo = {inversed_pp_95_10,inversed_pp_95_9,inversed_pp_95_8,inversed_pp_95_7,
    inversed_pp_95_6,inversed_pp_95_5,wallace_tree_cells_95_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_95_io_i_s_hi_lo = {inversed_pp_95_15,inversed_pp_95_14,inversed_pp_95_13,
    inversed_pp_95_12,inversed_pp_95_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_95_io_i_s_hi = {inversed_pp_95_21,inversed_pp_95_20,inversed_pp_95_19,inversed_pp_95_18
    ,inversed_pp_95_17,inversed_pp_95_16,wallace_tree_cells_95_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_96_io_i_s_lo_lo = {inversed_pp_96_4,inversed_pp_96_3,inversed_pp_96_2,inversed_pp_96_1,
    inversed_pp_96_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_96_io_i_s_lo = {inversed_pp_96_10,inversed_pp_96_9,inversed_pp_96_8,inversed_pp_96_7,
    inversed_pp_96_6,inversed_pp_96_5,wallace_tree_cells_96_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_96_io_i_s_hi_lo = {inversed_pp_96_15,inversed_pp_96_14,inversed_pp_96_13,
    inversed_pp_96_12,inversed_pp_96_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_96_io_i_s_hi = {inversed_pp_96_21,inversed_pp_96_20,inversed_pp_96_19,inversed_pp_96_18
    ,inversed_pp_96_17,inversed_pp_96_16,wallace_tree_cells_96_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_97_io_i_s_lo_lo = {inversed_pp_97_4,inversed_pp_97_3,inversed_pp_97_2,inversed_pp_97_1,
    inversed_pp_97_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_97_io_i_s_lo = {inversed_pp_97_10,inversed_pp_97_9,inversed_pp_97_8,inversed_pp_97_7,
    inversed_pp_97_6,inversed_pp_97_5,wallace_tree_cells_97_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_97_io_i_s_hi_lo = {inversed_pp_97_15,inversed_pp_97_14,inversed_pp_97_13,
    inversed_pp_97_12,inversed_pp_97_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_97_io_i_s_hi = {inversed_pp_97_21,inversed_pp_97_20,inversed_pp_97_19,inversed_pp_97_18
    ,inversed_pp_97_17,inversed_pp_97_16,wallace_tree_cells_97_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_98_io_i_s_lo_lo = {inversed_pp_98_4,inversed_pp_98_3,inversed_pp_98_2,inversed_pp_98_1,
    inversed_pp_98_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_98_io_i_s_lo = {inversed_pp_98_10,inversed_pp_98_9,inversed_pp_98_8,inversed_pp_98_7,
    inversed_pp_98_6,inversed_pp_98_5,wallace_tree_cells_98_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_98_io_i_s_hi_lo = {inversed_pp_98_15,inversed_pp_98_14,inversed_pp_98_13,
    inversed_pp_98_12,inversed_pp_98_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_98_io_i_s_hi = {inversed_pp_98_21,inversed_pp_98_20,inversed_pp_98_19,inversed_pp_98_18
    ,inversed_pp_98_17,inversed_pp_98_16,wallace_tree_cells_98_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_99_io_i_s_lo_lo = {inversed_pp_99_4,inversed_pp_99_3,inversed_pp_99_2,inversed_pp_99_1,
    inversed_pp_99_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_99_io_i_s_lo = {inversed_pp_99_10,inversed_pp_99_9,inversed_pp_99_8,inversed_pp_99_7,
    inversed_pp_99_6,inversed_pp_99_5,wallace_tree_cells_99_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_99_io_i_s_hi_lo = {inversed_pp_99_15,inversed_pp_99_14,inversed_pp_99_13,
    inversed_pp_99_12,inversed_pp_99_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_99_io_i_s_hi = {inversed_pp_99_21,inversed_pp_99_20,inversed_pp_99_19,inversed_pp_99_18
    ,inversed_pp_99_17,inversed_pp_99_16,wallace_tree_cells_99_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_100_io_i_s_lo_lo = {inversed_pp_100_4,inversed_pp_100_3,inversed_pp_100_2,
    inversed_pp_100_1,inversed_pp_100_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_100_io_i_s_lo = {inversed_pp_100_10,inversed_pp_100_9,inversed_pp_100_8,
    inversed_pp_100_7,inversed_pp_100_6,inversed_pp_100_5,wallace_tree_cells_100_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_100_io_i_s_hi_lo = {inversed_pp_100_15,inversed_pp_100_14,inversed_pp_100_13,
    inversed_pp_100_12,inversed_pp_100_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_100_io_i_s_hi = {inversed_pp_100_21,inversed_pp_100_20,inversed_pp_100_19,
    inversed_pp_100_18,inversed_pp_100_17,inversed_pp_100_16,wallace_tree_cells_100_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_101_io_i_s_lo_lo = {inversed_pp_101_4,inversed_pp_101_3,inversed_pp_101_2,
    inversed_pp_101_1,inversed_pp_101_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_101_io_i_s_lo = {inversed_pp_101_10,inversed_pp_101_9,inversed_pp_101_8,
    inversed_pp_101_7,inversed_pp_101_6,inversed_pp_101_5,wallace_tree_cells_101_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_101_io_i_s_hi_lo = {inversed_pp_101_15,inversed_pp_101_14,inversed_pp_101_13,
    inversed_pp_101_12,inversed_pp_101_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_101_io_i_s_hi = {inversed_pp_101_21,inversed_pp_101_20,inversed_pp_101_19,
    inversed_pp_101_18,inversed_pp_101_17,inversed_pp_101_16,wallace_tree_cells_101_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_102_io_i_s_lo_lo = {inversed_pp_102_4,inversed_pp_102_3,inversed_pp_102_2,
    inversed_pp_102_1,inversed_pp_102_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_102_io_i_s_lo = {inversed_pp_102_10,inversed_pp_102_9,inversed_pp_102_8,
    inversed_pp_102_7,inversed_pp_102_6,inversed_pp_102_5,wallace_tree_cells_102_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_102_io_i_s_hi_lo = {inversed_pp_102_15,inversed_pp_102_14,inversed_pp_102_13,
    inversed_pp_102_12,inversed_pp_102_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_102_io_i_s_hi = {inversed_pp_102_21,inversed_pp_102_20,inversed_pp_102_19,
    inversed_pp_102_18,inversed_pp_102_17,inversed_pp_102_16,wallace_tree_cells_102_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_103_io_i_s_lo_lo = {inversed_pp_103_4,inversed_pp_103_3,inversed_pp_103_2,
    inversed_pp_103_1,inversed_pp_103_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_103_io_i_s_lo = {inversed_pp_103_10,inversed_pp_103_9,inversed_pp_103_8,
    inversed_pp_103_7,inversed_pp_103_6,inversed_pp_103_5,wallace_tree_cells_103_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_103_io_i_s_hi_lo = {inversed_pp_103_15,inversed_pp_103_14,inversed_pp_103_13,
    inversed_pp_103_12,inversed_pp_103_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_103_io_i_s_hi = {inversed_pp_103_21,inversed_pp_103_20,inversed_pp_103_19,
    inversed_pp_103_18,inversed_pp_103_17,inversed_pp_103_16,wallace_tree_cells_103_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_104_io_i_s_lo_lo = {inversed_pp_104_4,inversed_pp_104_3,inversed_pp_104_2,
    inversed_pp_104_1,inversed_pp_104_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_104_io_i_s_lo = {inversed_pp_104_10,inversed_pp_104_9,inversed_pp_104_8,
    inversed_pp_104_7,inversed_pp_104_6,inversed_pp_104_5,wallace_tree_cells_104_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_104_io_i_s_hi_lo = {inversed_pp_104_15,inversed_pp_104_14,inversed_pp_104_13,
    inversed_pp_104_12,inversed_pp_104_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_104_io_i_s_hi = {inversed_pp_104_21,inversed_pp_104_20,inversed_pp_104_19,
    inversed_pp_104_18,inversed_pp_104_17,inversed_pp_104_16,wallace_tree_cells_104_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_105_io_i_s_lo_lo = {inversed_pp_105_4,inversed_pp_105_3,inversed_pp_105_2,
    inversed_pp_105_1,inversed_pp_105_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_105_io_i_s_lo = {inversed_pp_105_10,inversed_pp_105_9,inversed_pp_105_8,
    inversed_pp_105_7,inversed_pp_105_6,inversed_pp_105_5,wallace_tree_cells_105_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_105_io_i_s_hi_lo = {inversed_pp_105_15,inversed_pp_105_14,inversed_pp_105_13,
    inversed_pp_105_12,inversed_pp_105_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_105_io_i_s_hi = {inversed_pp_105_21,inversed_pp_105_20,inversed_pp_105_19,
    inversed_pp_105_18,inversed_pp_105_17,inversed_pp_105_16,wallace_tree_cells_105_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_106_io_i_s_lo_lo = {inversed_pp_106_4,inversed_pp_106_3,inversed_pp_106_2,
    inversed_pp_106_1,inversed_pp_106_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_106_io_i_s_lo = {inversed_pp_106_10,inversed_pp_106_9,inversed_pp_106_8,
    inversed_pp_106_7,inversed_pp_106_6,inversed_pp_106_5,wallace_tree_cells_106_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_106_io_i_s_hi_lo = {inversed_pp_106_15,inversed_pp_106_14,inversed_pp_106_13,
    inversed_pp_106_12,inversed_pp_106_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_106_io_i_s_hi = {inversed_pp_106_21,inversed_pp_106_20,inversed_pp_106_19,
    inversed_pp_106_18,inversed_pp_106_17,inversed_pp_106_16,wallace_tree_cells_106_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_107_io_i_s_lo_lo = {inversed_pp_107_4,inversed_pp_107_3,inversed_pp_107_2,
    inversed_pp_107_1,inversed_pp_107_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_107_io_i_s_lo = {inversed_pp_107_10,inversed_pp_107_9,inversed_pp_107_8,
    inversed_pp_107_7,inversed_pp_107_6,inversed_pp_107_5,wallace_tree_cells_107_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_107_io_i_s_hi_lo = {inversed_pp_107_15,inversed_pp_107_14,inversed_pp_107_13,
    inversed_pp_107_12,inversed_pp_107_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_107_io_i_s_hi = {inversed_pp_107_21,inversed_pp_107_20,inversed_pp_107_19,
    inversed_pp_107_18,inversed_pp_107_17,inversed_pp_107_16,wallace_tree_cells_107_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_108_io_i_s_lo_lo = {inversed_pp_108_4,inversed_pp_108_3,inversed_pp_108_2,
    inversed_pp_108_1,inversed_pp_108_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_108_io_i_s_lo = {inversed_pp_108_10,inversed_pp_108_9,inversed_pp_108_8,
    inversed_pp_108_7,inversed_pp_108_6,inversed_pp_108_5,wallace_tree_cells_108_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_108_io_i_s_hi_lo = {inversed_pp_108_15,inversed_pp_108_14,inversed_pp_108_13,
    inversed_pp_108_12,inversed_pp_108_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_108_io_i_s_hi = {inversed_pp_108_21,inversed_pp_108_20,inversed_pp_108_19,
    inversed_pp_108_18,inversed_pp_108_17,inversed_pp_108_16,wallace_tree_cells_108_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_109_io_i_s_lo_lo = {inversed_pp_109_4,inversed_pp_109_3,inversed_pp_109_2,
    inversed_pp_109_1,inversed_pp_109_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_109_io_i_s_lo = {inversed_pp_109_10,inversed_pp_109_9,inversed_pp_109_8,
    inversed_pp_109_7,inversed_pp_109_6,inversed_pp_109_5,wallace_tree_cells_109_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_109_io_i_s_hi_lo = {inversed_pp_109_15,inversed_pp_109_14,inversed_pp_109_13,
    inversed_pp_109_12,inversed_pp_109_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_109_io_i_s_hi = {inversed_pp_109_21,inversed_pp_109_20,inversed_pp_109_19,
    inversed_pp_109_18,inversed_pp_109_17,inversed_pp_109_16,wallace_tree_cells_109_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_110_io_i_s_lo_lo = {inversed_pp_110_4,inversed_pp_110_3,inversed_pp_110_2,
    inversed_pp_110_1,inversed_pp_110_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_110_io_i_s_lo = {inversed_pp_110_10,inversed_pp_110_9,inversed_pp_110_8,
    inversed_pp_110_7,inversed_pp_110_6,inversed_pp_110_5,wallace_tree_cells_110_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_110_io_i_s_hi_lo = {inversed_pp_110_15,inversed_pp_110_14,inversed_pp_110_13,
    inversed_pp_110_12,inversed_pp_110_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_110_io_i_s_hi = {inversed_pp_110_21,inversed_pp_110_20,inversed_pp_110_19,
    inversed_pp_110_18,inversed_pp_110_17,inversed_pp_110_16,wallace_tree_cells_110_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_111_io_i_s_lo_lo = {inversed_pp_111_4,inversed_pp_111_3,inversed_pp_111_2,
    inversed_pp_111_1,inversed_pp_111_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_111_io_i_s_lo = {inversed_pp_111_10,inversed_pp_111_9,inversed_pp_111_8,
    inversed_pp_111_7,inversed_pp_111_6,inversed_pp_111_5,wallace_tree_cells_111_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_111_io_i_s_hi_lo = {inversed_pp_111_15,inversed_pp_111_14,inversed_pp_111_13,
    inversed_pp_111_12,inversed_pp_111_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_111_io_i_s_hi = {inversed_pp_111_21,inversed_pp_111_20,inversed_pp_111_19,
    inversed_pp_111_18,inversed_pp_111_17,inversed_pp_111_16,wallace_tree_cells_111_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_112_io_i_s_lo_lo = {inversed_pp_112_4,inversed_pp_112_3,inversed_pp_112_2,
    inversed_pp_112_1,inversed_pp_112_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_112_io_i_s_lo = {inversed_pp_112_10,inversed_pp_112_9,inversed_pp_112_8,
    inversed_pp_112_7,inversed_pp_112_6,inversed_pp_112_5,wallace_tree_cells_112_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_112_io_i_s_hi_lo = {inversed_pp_112_15,inversed_pp_112_14,inversed_pp_112_13,
    inversed_pp_112_12,inversed_pp_112_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_112_io_i_s_hi = {inversed_pp_112_21,inversed_pp_112_20,inversed_pp_112_19,
    inversed_pp_112_18,inversed_pp_112_17,inversed_pp_112_16,wallace_tree_cells_112_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_113_io_i_s_lo_lo = {inversed_pp_113_4,inversed_pp_113_3,inversed_pp_113_2,
    inversed_pp_113_1,inversed_pp_113_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_113_io_i_s_lo = {inversed_pp_113_10,inversed_pp_113_9,inversed_pp_113_8,
    inversed_pp_113_7,inversed_pp_113_6,inversed_pp_113_5,wallace_tree_cells_113_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_113_io_i_s_hi_lo = {inversed_pp_113_15,inversed_pp_113_14,inversed_pp_113_13,
    inversed_pp_113_12,inversed_pp_113_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_113_io_i_s_hi = {inversed_pp_113_21,inversed_pp_113_20,inversed_pp_113_19,
    inversed_pp_113_18,inversed_pp_113_17,inversed_pp_113_16,wallace_tree_cells_113_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_114_io_i_s_lo_lo = {inversed_pp_114_4,inversed_pp_114_3,inversed_pp_114_2,
    inversed_pp_114_1,inversed_pp_114_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_114_io_i_s_lo = {inversed_pp_114_10,inversed_pp_114_9,inversed_pp_114_8,
    inversed_pp_114_7,inversed_pp_114_6,inversed_pp_114_5,wallace_tree_cells_114_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_114_io_i_s_hi_lo = {inversed_pp_114_15,inversed_pp_114_14,inversed_pp_114_13,
    inversed_pp_114_12,inversed_pp_114_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_114_io_i_s_hi = {inversed_pp_114_21,inversed_pp_114_20,inversed_pp_114_19,
    inversed_pp_114_18,inversed_pp_114_17,inversed_pp_114_16,wallace_tree_cells_114_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_115_io_i_s_lo_lo = {inversed_pp_115_4,inversed_pp_115_3,inversed_pp_115_2,
    inversed_pp_115_1,inversed_pp_115_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_115_io_i_s_lo = {inversed_pp_115_10,inversed_pp_115_9,inversed_pp_115_8,
    inversed_pp_115_7,inversed_pp_115_6,inversed_pp_115_5,wallace_tree_cells_115_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_115_io_i_s_hi_lo = {inversed_pp_115_15,inversed_pp_115_14,inversed_pp_115_13,
    inversed_pp_115_12,inversed_pp_115_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_115_io_i_s_hi = {inversed_pp_115_21,inversed_pp_115_20,inversed_pp_115_19,
    inversed_pp_115_18,inversed_pp_115_17,inversed_pp_115_16,wallace_tree_cells_115_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_116_io_i_s_lo_lo = {inversed_pp_116_4,inversed_pp_116_3,inversed_pp_116_2,
    inversed_pp_116_1,inversed_pp_116_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_116_io_i_s_lo = {inversed_pp_116_10,inversed_pp_116_9,inversed_pp_116_8,
    inversed_pp_116_7,inversed_pp_116_6,inversed_pp_116_5,wallace_tree_cells_116_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_116_io_i_s_hi_lo = {inversed_pp_116_15,inversed_pp_116_14,inversed_pp_116_13,
    inversed_pp_116_12,inversed_pp_116_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_116_io_i_s_hi = {inversed_pp_116_21,inversed_pp_116_20,inversed_pp_116_19,
    inversed_pp_116_18,inversed_pp_116_17,inversed_pp_116_16,wallace_tree_cells_116_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_117_io_i_s_lo_lo = {inversed_pp_117_4,inversed_pp_117_3,inversed_pp_117_2,
    inversed_pp_117_1,inversed_pp_117_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_117_io_i_s_lo = {inversed_pp_117_10,inversed_pp_117_9,inversed_pp_117_8,
    inversed_pp_117_7,inversed_pp_117_6,inversed_pp_117_5,wallace_tree_cells_117_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_117_io_i_s_hi_lo = {inversed_pp_117_15,inversed_pp_117_14,inversed_pp_117_13,
    inversed_pp_117_12,inversed_pp_117_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_117_io_i_s_hi = {inversed_pp_117_21,inversed_pp_117_20,inversed_pp_117_19,
    inversed_pp_117_18,inversed_pp_117_17,inversed_pp_117_16,wallace_tree_cells_117_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_118_io_i_s_lo_lo = {inversed_pp_118_4,inversed_pp_118_3,inversed_pp_118_2,
    inversed_pp_118_1,inversed_pp_118_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_118_io_i_s_lo = {inversed_pp_118_10,inversed_pp_118_9,inversed_pp_118_8,
    inversed_pp_118_7,inversed_pp_118_6,inversed_pp_118_5,wallace_tree_cells_118_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_118_io_i_s_hi_lo = {inversed_pp_118_15,inversed_pp_118_14,inversed_pp_118_13,
    inversed_pp_118_12,inversed_pp_118_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_118_io_i_s_hi = {inversed_pp_118_21,inversed_pp_118_20,inversed_pp_118_19,
    inversed_pp_118_18,inversed_pp_118_17,inversed_pp_118_16,wallace_tree_cells_118_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_119_io_i_s_lo_lo = {inversed_pp_119_4,inversed_pp_119_3,inversed_pp_119_2,
    inversed_pp_119_1,inversed_pp_119_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_119_io_i_s_lo = {inversed_pp_119_10,inversed_pp_119_9,inversed_pp_119_8,
    inversed_pp_119_7,inversed_pp_119_6,inversed_pp_119_5,wallace_tree_cells_119_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_119_io_i_s_hi_lo = {inversed_pp_119_15,inversed_pp_119_14,inversed_pp_119_13,
    inversed_pp_119_12,inversed_pp_119_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_119_io_i_s_hi = {inversed_pp_119_21,inversed_pp_119_20,inversed_pp_119_19,
    inversed_pp_119_18,inversed_pp_119_17,inversed_pp_119_16,wallace_tree_cells_119_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_120_io_i_s_lo_lo = {inversed_pp_120_4,inversed_pp_120_3,inversed_pp_120_2,
    inversed_pp_120_1,inversed_pp_120_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_120_io_i_s_lo = {inversed_pp_120_10,inversed_pp_120_9,inversed_pp_120_8,
    inversed_pp_120_7,inversed_pp_120_6,inversed_pp_120_5,wallace_tree_cells_120_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_120_io_i_s_hi_lo = {inversed_pp_120_15,inversed_pp_120_14,inversed_pp_120_13,
    inversed_pp_120_12,inversed_pp_120_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_120_io_i_s_hi = {inversed_pp_120_21,inversed_pp_120_20,inversed_pp_120_19,
    inversed_pp_120_18,inversed_pp_120_17,inversed_pp_120_16,wallace_tree_cells_120_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_121_io_i_s_lo_lo = {inversed_pp_121_4,inversed_pp_121_3,inversed_pp_121_2,
    inversed_pp_121_1,inversed_pp_121_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_121_io_i_s_lo = {inversed_pp_121_10,inversed_pp_121_9,inversed_pp_121_8,
    inversed_pp_121_7,inversed_pp_121_6,inversed_pp_121_5,wallace_tree_cells_121_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_121_io_i_s_hi_lo = {inversed_pp_121_15,inversed_pp_121_14,inversed_pp_121_13,
    inversed_pp_121_12,inversed_pp_121_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_121_io_i_s_hi = {inversed_pp_121_21,inversed_pp_121_20,inversed_pp_121_19,
    inversed_pp_121_18,inversed_pp_121_17,inversed_pp_121_16,wallace_tree_cells_121_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_122_io_i_s_lo_lo = {inversed_pp_122_4,inversed_pp_122_3,inversed_pp_122_2,
    inversed_pp_122_1,inversed_pp_122_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_122_io_i_s_lo = {inversed_pp_122_10,inversed_pp_122_9,inversed_pp_122_8,
    inversed_pp_122_7,inversed_pp_122_6,inversed_pp_122_5,wallace_tree_cells_122_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_122_io_i_s_hi_lo = {inversed_pp_122_15,inversed_pp_122_14,inversed_pp_122_13,
    inversed_pp_122_12,inversed_pp_122_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_122_io_i_s_hi = {inversed_pp_122_21,inversed_pp_122_20,inversed_pp_122_19,
    inversed_pp_122_18,inversed_pp_122_17,inversed_pp_122_16,wallace_tree_cells_122_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_123_io_i_s_lo_lo = {inversed_pp_123_4,inversed_pp_123_3,inversed_pp_123_2,
    inversed_pp_123_1,inversed_pp_123_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_123_io_i_s_lo = {inversed_pp_123_10,inversed_pp_123_9,inversed_pp_123_8,
    inversed_pp_123_7,inversed_pp_123_6,inversed_pp_123_5,wallace_tree_cells_123_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_123_io_i_s_hi_lo = {inversed_pp_123_15,inversed_pp_123_14,inversed_pp_123_13,
    inversed_pp_123_12,inversed_pp_123_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_123_io_i_s_hi = {inversed_pp_123_21,inversed_pp_123_20,inversed_pp_123_19,
    inversed_pp_123_18,inversed_pp_123_17,inversed_pp_123_16,wallace_tree_cells_123_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_124_io_i_s_lo_lo = {inversed_pp_124_4,inversed_pp_124_3,inversed_pp_124_2,
    inversed_pp_124_1,inversed_pp_124_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_124_io_i_s_lo = {inversed_pp_124_10,inversed_pp_124_9,inversed_pp_124_8,
    inversed_pp_124_7,inversed_pp_124_6,inversed_pp_124_5,wallace_tree_cells_124_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_124_io_i_s_hi_lo = {inversed_pp_124_15,inversed_pp_124_14,inversed_pp_124_13,
    inversed_pp_124_12,inversed_pp_124_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_124_io_i_s_hi = {inversed_pp_124_21,inversed_pp_124_20,inversed_pp_124_19,
    inversed_pp_124_18,inversed_pp_124_17,inversed_pp_124_16,wallace_tree_cells_124_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_125_io_i_s_lo_lo = {inversed_pp_125_4,inversed_pp_125_3,inversed_pp_125_2,
    inversed_pp_125_1,inversed_pp_125_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_125_io_i_s_lo = {inversed_pp_125_10,inversed_pp_125_9,inversed_pp_125_8,
    inversed_pp_125_7,inversed_pp_125_6,inversed_pp_125_5,wallace_tree_cells_125_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_125_io_i_s_hi_lo = {inversed_pp_125_15,inversed_pp_125_14,inversed_pp_125_13,
    inversed_pp_125_12,inversed_pp_125_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_125_io_i_s_hi = {inversed_pp_125_21,inversed_pp_125_20,inversed_pp_125_19,
    inversed_pp_125_18,inversed_pp_125_17,inversed_pp_125_16,wallace_tree_cells_125_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_126_io_i_s_lo_lo = {inversed_pp_126_4,inversed_pp_126_3,inversed_pp_126_2,
    inversed_pp_126_1,inversed_pp_126_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_126_io_i_s_lo = {inversed_pp_126_10,inversed_pp_126_9,inversed_pp_126_8,
    inversed_pp_126_7,inversed_pp_126_6,inversed_pp_126_5,wallace_tree_cells_126_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_126_io_i_s_hi_lo = {inversed_pp_126_15,inversed_pp_126_14,inversed_pp_126_13,
    inversed_pp_126_12,inversed_pp_126_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_126_io_i_s_hi = {inversed_pp_126_21,inversed_pp_126_20,inversed_pp_126_19,
    inversed_pp_126_18,inversed_pp_126_17,inversed_pp_126_16,wallace_tree_cells_126_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_127_io_i_s_lo_lo = {inversed_pp_127_4,inversed_pp_127_3,inversed_pp_127_2,
    inversed_pp_127_1,inversed_pp_127_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_127_io_i_s_lo = {inversed_pp_127_10,inversed_pp_127_9,inversed_pp_127_8,
    inversed_pp_127_7,inversed_pp_127_6,inversed_pp_127_5,wallace_tree_cells_127_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_127_io_i_s_hi_lo = {inversed_pp_127_15,inversed_pp_127_14,inversed_pp_127_13,
    inversed_pp_127_12,inversed_pp_127_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_127_io_i_s_hi = {inversed_pp_127_21,inversed_pp_127_20,inversed_pp_127_19,
    inversed_pp_127_18,inversed_pp_127_17,inversed_pp_127_16,wallace_tree_cells_127_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_128_io_i_s_lo_lo = {inversed_pp_128_4,inversed_pp_128_3,inversed_pp_128_2,
    inversed_pp_128_1,inversed_pp_128_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_128_io_i_s_lo = {inversed_pp_128_10,inversed_pp_128_9,inversed_pp_128_8,
    inversed_pp_128_7,inversed_pp_128_6,inversed_pp_128_5,wallace_tree_cells_128_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_128_io_i_s_hi_lo = {inversed_pp_128_15,inversed_pp_128_14,inversed_pp_128_13,
    inversed_pp_128_12,inversed_pp_128_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_128_io_i_s_hi = {inversed_pp_128_21,inversed_pp_128_20,inversed_pp_128_19,
    inversed_pp_128_18,inversed_pp_128_17,inversed_pp_128_16,wallace_tree_cells_128_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_129_io_i_s_lo_lo = {inversed_pp_129_4,inversed_pp_129_3,inversed_pp_129_2,
    inversed_pp_129_1,inversed_pp_129_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_129_io_i_s_lo = {inversed_pp_129_10,inversed_pp_129_9,inversed_pp_129_8,
    inversed_pp_129_7,inversed_pp_129_6,inversed_pp_129_5,wallace_tree_cells_129_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_129_io_i_s_hi_lo = {inversed_pp_129_15,inversed_pp_129_14,inversed_pp_129_13,
    inversed_pp_129_12,inversed_pp_129_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_129_io_i_s_hi = {inversed_pp_129_21,inversed_pp_129_20,inversed_pp_129_19,
    inversed_pp_129_18,inversed_pp_129_17,inversed_pp_129_16,wallace_tree_cells_129_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_130_io_i_s_lo_lo = {inversed_pp_130_4,inversed_pp_130_3,inversed_pp_130_2,
    inversed_pp_130_1,inversed_pp_130_0}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_130_io_i_s_lo = {inversed_pp_130_10,inversed_pp_130_9,inversed_pp_130_8,
    inversed_pp_130_7,inversed_pp_130_6,inversed_pp_130_5,wallace_tree_cells_130_io_i_s_lo_lo}; // @[wallace_tree.scala 147:56]
  wire [4:0] wallace_tree_cells_130_io_i_s_hi_lo = {inversed_pp_130_15,inversed_pp_130_14,inversed_pp_130_13,
    inversed_pp_130_12,inversed_pp_130_11}; // @[wallace_tree.scala 147:56]
  wire [10:0] wallace_tree_cells_130_io_i_s_hi = {inversed_pp_130_21,inversed_pp_130_20,inversed_pp_130_19,
    inversed_pp_130_18,inversed_pp_130_17,inversed_pp_130_16,wallace_tree_cells_130_io_i_s_hi_lo}; // @[wallace_tree.scala 147:56]
  wire  s_1 = wallace_tree_cells_1_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_0 = wallace_tree_cells_0_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_3 = wallace_tree_cells_3_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_2 = wallace_tree_cells_2_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_5 = wallace_tree_cells_5_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_4 = wallace_tree_cells_4_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_7 = wallace_tree_cells_7_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_6 = wallace_tree_cells_6_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_lo_lo_lo_lo = {s_7,s_6,s_5,s_4,s_3,s_2,s_1,s_0}; // @[wallace_tree.scala 156:17]
  wire  s_9 = wallace_tree_cells_9_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_8 = wallace_tree_cells_8_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_11 = wallace_tree_cells_11_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_10 = wallace_tree_cells_10_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_13 = wallace_tree_cells_13_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_12 = wallace_tree_cells_12_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_15 = wallace_tree_cells_15_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_14 = wallace_tree_cells_14_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [15:0] io_o_s_lo_lo_lo = {s_15,s_14,s_13,s_12,s_11,s_10,s_9,s_8,io_o_s_lo_lo_lo_lo}; // @[wallace_tree.scala 156:17]
  wire  s_17 = wallace_tree_cells_17_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_16 = wallace_tree_cells_16_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_19 = wallace_tree_cells_19_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_18 = wallace_tree_cells_18_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_21 = wallace_tree_cells_21_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_20 = wallace_tree_cells_20_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_23 = wallace_tree_cells_23_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_22 = wallace_tree_cells_22_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_lo_lo_hi_lo = {s_23,s_22,s_21,s_20,s_19,s_18,s_17,s_16}; // @[wallace_tree.scala 156:17]
  wire  s_25 = wallace_tree_cells_25_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_24 = wallace_tree_cells_24_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_27 = wallace_tree_cells_27_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_26 = wallace_tree_cells_26_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_29 = wallace_tree_cells_29_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_28 = wallace_tree_cells_28_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_31 = wallace_tree_cells_31_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_30 = wallace_tree_cells_30_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [31:0] io_o_s_lo_lo = {s_31,s_30,s_29,s_28,s_27,s_26,s_25,s_24,io_o_s_lo_lo_hi_lo,io_o_s_lo_lo_lo}; // @[wallace_tree.scala 156:17]
  wire  s_33 = wallace_tree_cells_33_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_32 = wallace_tree_cells_32_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_35 = wallace_tree_cells_35_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_34 = wallace_tree_cells_34_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_37 = wallace_tree_cells_37_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_36 = wallace_tree_cells_36_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_39 = wallace_tree_cells_39_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_38 = wallace_tree_cells_38_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_lo_hi_lo_lo = {s_39,s_38,s_37,s_36,s_35,s_34,s_33,s_32}; // @[wallace_tree.scala 156:17]
  wire  s_41 = wallace_tree_cells_41_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_40 = wallace_tree_cells_40_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_43 = wallace_tree_cells_43_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_42 = wallace_tree_cells_42_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_45 = wallace_tree_cells_45_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_44 = wallace_tree_cells_44_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_47 = wallace_tree_cells_47_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_46 = wallace_tree_cells_46_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_49 = wallace_tree_cells_49_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_48 = wallace_tree_cells_48_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_51 = wallace_tree_cells_51_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_50 = wallace_tree_cells_50_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_53 = wallace_tree_cells_53_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_52 = wallace_tree_cells_52_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_55 = wallace_tree_cells_55_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_54 = wallace_tree_cells_54_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_lo_hi_hi_lo = {s_55,s_54,s_53,s_52,s_51,s_50,s_49,s_48}; // @[wallace_tree.scala 156:17]
  wire  s_57 = wallace_tree_cells_57_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_56 = wallace_tree_cells_56_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_59 = wallace_tree_cells_59_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_58 = wallace_tree_cells_58_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_61 = wallace_tree_cells_61_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_60 = wallace_tree_cells_60_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_64 = wallace_tree_cells_64_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_63 = wallace_tree_cells_63_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_62 = wallace_tree_cells_62_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [16:0] io_o_s_lo_hi_hi = {s_64,s_63,s_62,s_61,s_60,s_59,s_58,s_57,s_56,io_o_s_lo_hi_hi_lo}; // @[wallace_tree.scala 156:17]
  wire [32:0] io_o_s_lo_hi = {io_o_s_lo_hi_hi,s_47,s_46,s_45,s_44,s_43,s_42,s_41,s_40,io_o_s_lo_hi_lo_lo}; // @[wallace_tree.scala 156:17]
  wire [64:0] io_o_s_lo = {io_o_s_lo_hi,io_o_s_lo_lo}; // @[wallace_tree.scala 156:17]
  wire  s_66 = wallace_tree_cells_66_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_65 = wallace_tree_cells_65_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_68 = wallace_tree_cells_68_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_67 = wallace_tree_cells_67_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_70 = wallace_tree_cells_70_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_69 = wallace_tree_cells_69_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_72 = wallace_tree_cells_72_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_71 = wallace_tree_cells_71_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_hi_lo_lo_lo = {s_72,s_71,s_70,s_69,s_68,s_67,s_66,s_65}; // @[wallace_tree.scala 156:17]
  wire  s_74 = wallace_tree_cells_74_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_73 = wallace_tree_cells_73_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_76 = wallace_tree_cells_76_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_75 = wallace_tree_cells_75_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_78 = wallace_tree_cells_78_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_77 = wallace_tree_cells_77_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_80 = wallace_tree_cells_80_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_79 = wallace_tree_cells_79_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_82 = wallace_tree_cells_82_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_81 = wallace_tree_cells_81_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_84 = wallace_tree_cells_84_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_83 = wallace_tree_cells_83_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_86 = wallace_tree_cells_86_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_85 = wallace_tree_cells_85_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_88 = wallace_tree_cells_88_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_87 = wallace_tree_cells_87_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_hi_lo_hi_lo = {s_88,s_87,s_86,s_85,s_84,s_83,s_82,s_81}; // @[wallace_tree.scala 156:17]
  wire  s_90 = wallace_tree_cells_90_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_89 = wallace_tree_cells_89_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_92 = wallace_tree_cells_92_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_91 = wallace_tree_cells_91_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_94 = wallace_tree_cells_94_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_93 = wallace_tree_cells_93_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_97 = wallace_tree_cells_97_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_96 = wallace_tree_cells_96_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_95 = wallace_tree_cells_95_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [16:0] io_o_s_hi_lo_hi = {s_97,s_96,s_95,s_94,s_93,s_92,s_91,s_90,s_89,io_o_s_hi_lo_hi_lo}; // @[wallace_tree.scala 156:17]
  wire [32:0] io_o_s_hi_lo = {io_o_s_hi_lo_hi,s_80,s_79,s_78,s_77,s_76,s_75,s_74,s_73,io_o_s_hi_lo_lo_lo}; // @[wallace_tree.scala 156:17]
  wire  s_99 = wallace_tree_cells_99_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_98 = wallace_tree_cells_98_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_101 = wallace_tree_cells_101_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_100 = wallace_tree_cells_100_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_103 = wallace_tree_cells_103_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_102 = wallace_tree_cells_102_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_105 = wallace_tree_cells_105_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_104 = wallace_tree_cells_104_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_hi_hi_lo_lo = {s_105,s_104,s_103,s_102,s_101,s_100,s_99,s_98}; // @[wallace_tree.scala 156:17]
  wire  s_107 = wallace_tree_cells_107_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_106 = wallace_tree_cells_106_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_109 = wallace_tree_cells_109_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_108 = wallace_tree_cells_108_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_111 = wallace_tree_cells_111_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_110 = wallace_tree_cells_110_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_113 = wallace_tree_cells_113_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_112 = wallace_tree_cells_112_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_115 = wallace_tree_cells_115_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_114 = wallace_tree_cells_114_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_117 = wallace_tree_cells_117_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_116 = wallace_tree_cells_116_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_119 = wallace_tree_cells_119_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_118 = wallace_tree_cells_118_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_121 = wallace_tree_cells_121_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_120 = wallace_tree_cells_120_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [7:0] io_o_s_hi_hi_hi_lo = {s_121,s_120,s_119,s_118,s_117,s_116,s_115,s_114}; // @[wallace_tree.scala 156:17]
  wire  s_123 = wallace_tree_cells_123_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_122 = wallace_tree_cells_122_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_125 = wallace_tree_cells_125_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_124 = wallace_tree_cells_124_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_127 = wallace_tree_cells_127_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_126 = wallace_tree_cells_126_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_130 = wallace_tree_cells_130_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_129 = wallace_tree_cells_129_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire  s_128 = wallace_tree_cells_128_io_o_s; // @[wallace_tree.scala 154:17 160:14]
  wire [16:0] io_o_s_hi_hi_hi = {s_130,s_129,s_128,s_127,s_126,s_125,s_124,s_123,s_122,io_o_s_hi_hi_hi_lo}; // @[wallace_tree.scala 156:17]
  wire [32:0] io_o_s_hi_hi = {io_o_s_hi_hi_hi,s_113,s_112,s_111,s_110,s_109,s_108,s_107,s_106,io_o_s_hi_hi_lo_lo}; // @[wallace_tree.scala 156:17]
  wire [65:0] io_o_s_hi = {io_o_s_hi_hi,io_o_s_hi_lo}; // @[wallace_tree.scala 156:17]
  wire  c_1 = wallace_tree_cells_1_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_0 = wallace_tree_cells_0_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_3 = wallace_tree_cells_3_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_2 = wallace_tree_cells_2_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_5 = wallace_tree_cells_5_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_4 = wallace_tree_cells_4_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_7 = wallace_tree_cells_7_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_6 = wallace_tree_cells_6_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_lo_lo_lo_lo = {c_7,c_6,c_5,c_4,c_3,c_2,c_1,c_0}; // @[wallace_tree.scala 157:17]
  wire  c_9 = wallace_tree_cells_9_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_8 = wallace_tree_cells_8_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_11 = wallace_tree_cells_11_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_10 = wallace_tree_cells_10_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_13 = wallace_tree_cells_13_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_12 = wallace_tree_cells_12_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_15 = wallace_tree_cells_15_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_14 = wallace_tree_cells_14_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [15:0] io_o_c_lo_lo_lo = {c_15,c_14,c_13,c_12,c_11,c_10,c_9,c_8,io_o_c_lo_lo_lo_lo}; // @[wallace_tree.scala 157:17]
  wire  c_17 = wallace_tree_cells_17_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_16 = wallace_tree_cells_16_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_19 = wallace_tree_cells_19_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_18 = wallace_tree_cells_18_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_21 = wallace_tree_cells_21_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_20 = wallace_tree_cells_20_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_23 = wallace_tree_cells_23_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_22 = wallace_tree_cells_22_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_lo_lo_hi_lo = {c_23,c_22,c_21,c_20,c_19,c_18,c_17,c_16}; // @[wallace_tree.scala 157:17]
  wire  c_25 = wallace_tree_cells_25_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_24 = wallace_tree_cells_24_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_27 = wallace_tree_cells_27_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_26 = wallace_tree_cells_26_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_29 = wallace_tree_cells_29_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_28 = wallace_tree_cells_28_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_31 = wallace_tree_cells_31_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_30 = wallace_tree_cells_30_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [31:0] io_o_c_lo_lo = {c_31,c_30,c_29,c_28,c_27,c_26,c_25,c_24,io_o_c_lo_lo_hi_lo,io_o_c_lo_lo_lo}; // @[wallace_tree.scala 157:17]
  wire  c_33 = wallace_tree_cells_33_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_32 = wallace_tree_cells_32_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_35 = wallace_tree_cells_35_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_34 = wallace_tree_cells_34_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_37 = wallace_tree_cells_37_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_36 = wallace_tree_cells_36_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_39 = wallace_tree_cells_39_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_38 = wallace_tree_cells_38_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_lo_hi_lo_lo = {c_39,c_38,c_37,c_36,c_35,c_34,c_33,c_32}; // @[wallace_tree.scala 157:17]
  wire  c_41 = wallace_tree_cells_41_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_40 = wallace_tree_cells_40_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_43 = wallace_tree_cells_43_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_42 = wallace_tree_cells_42_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_45 = wallace_tree_cells_45_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_44 = wallace_tree_cells_44_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_47 = wallace_tree_cells_47_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_46 = wallace_tree_cells_46_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_49 = wallace_tree_cells_49_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_48 = wallace_tree_cells_48_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_51 = wallace_tree_cells_51_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_50 = wallace_tree_cells_50_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_53 = wallace_tree_cells_53_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_52 = wallace_tree_cells_52_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_55 = wallace_tree_cells_55_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_54 = wallace_tree_cells_54_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_lo_hi_hi_lo = {c_55,c_54,c_53,c_52,c_51,c_50,c_49,c_48}; // @[wallace_tree.scala 157:17]
  wire  c_57 = wallace_tree_cells_57_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_56 = wallace_tree_cells_56_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_59 = wallace_tree_cells_59_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_58 = wallace_tree_cells_58_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_61 = wallace_tree_cells_61_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_60 = wallace_tree_cells_60_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_64 = wallace_tree_cells_64_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_63 = wallace_tree_cells_63_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_62 = wallace_tree_cells_62_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [16:0] io_o_c_lo_hi_hi = {c_64,c_63,c_62,c_61,c_60,c_59,c_58,c_57,c_56,io_o_c_lo_hi_hi_lo}; // @[wallace_tree.scala 157:17]
  wire [32:0] io_o_c_lo_hi = {io_o_c_lo_hi_hi,c_47,c_46,c_45,c_44,c_43,c_42,c_41,c_40,io_o_c_lo_hi_lo_lo}; // @[wallace_tree.scala 157:17]
  wire [64:0] io_o_c_lo = {io_o_c_lo_hi,io_o_c_lo_lo}; // @[wallace_tree.scala 157:17]
  wire  c_66 = wallace_tree_cells_66_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_65 = wallace_tree_cells_65_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_68 = wallace_tree_cells_68_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_67 = wallace_tree_cells_67_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_70 = wallace_tree_cells_70_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_69 = wallace_tree_cells_69_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_72 = wallace_tree_cells_72_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_71 = wallace_tree_cells_71_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_hi_lo_lo_lo = {c_72,c_71,c_70,c_69,c_68,c_67,c_66,c_65}; // @[wallace_tree.scala 157:17]
  wire  c_74 = wallace_tree_cells_74_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_73 = wallace_tree_cells_73_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_76 = wallace_tree_cells_76_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_75 = wallace_tree_cells_75_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_78 = wallace_tree_cells_78_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_77 = wallace_tree_cells_77_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_80 = wallace_tree_cells_80_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_79 = wallace_tree_cells_79_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_82 = wallace_tree_cells_82_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_81 = wallace_tree_cells_81_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_84 = wallace_tree_cells_84_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_83 = wallace_tree_cells_83_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_86 = wallace_tree_cells_86_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_85 = wallace_tree_cells_85_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_88 = wallace_tree_cells_88_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_87 = wallace_tree_cells_87_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_hi_lo_hi_lo = {c_88,c_87,c_86,c_85,c_84,c_83,c_82,c_81}; // @[wallace_tree.scala 157:17]
  wire  c_90 = wallace_tree_cells_90_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_89 = wallace_tree_cells_89_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_92 = wallace_tree_cells_92_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_91 = wallace_tree_cells_91_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_94 = wallace_tree_cells_94_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_93 = wallace_tree_cells_93_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_97 = wallace_tree_cells_97_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_96 = wallace_tree_cells_96_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_95 = wallace_tree_cells_95_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [16:0] io_o_c_hi_lo_hi = {c_97,c_96,c_95,c_94,c_93,c_92,c_91,c_90,c_89,io_o_c_hi_lo_hi_lo}; // @[wallace_tree.scala 157:17]
  wire [32:0] io_o_c_hi_lo = {io_o_c_hi_lo_hi,c_80,c_79,c_78,c_77,c_76,c_75,c_74,c_73,io_o_c_hi_lo_lo_lo}; // @[wallace_tree.scala 157:17]
  wire  c_99 = wallace_tree_cells_99_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_98 = wallace_tree_cells_98_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_101 = wallace_tree_cells_101_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_100 = wallace_tree_cells_100_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_103 = wallace_tree_cells_103_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_102 = wallace_tree_cells_102_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_105 = wallace_tree_cells_105_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_104 = wallace_tree_cells_104_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_hi_hi_lo_lo = {c_105,c_104,c_103,c_102,c_101,c_100,c_99,c_98}; // @[wallace_tree.scala 157:17]
  wire  c_107 = wallace_tree_cells_107_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_106 = wallace_tree_cells_106_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_109 = wallace_tree_cells_109_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_108 = wallace_tree_cells_108_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_111 = wallace_tree_cells_111_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_110 = wallace_tree_cells_110_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_113 = wallace_tree_cells_113_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_112 = wallace_tree_cells_112_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_115 = wallace_tree_cells_115_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_114 = wallace_tree_cells_114_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_117 = wallace_tree_cells_117_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_116 = wallace_tree_cells_116_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_119 = wallace_tree_cells_119_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_118 = wallace_tree_cells_118_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_121 = wallace_tree_cells_121_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_120 = wallace_tree_cells_120_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [7:0] io_o_c_hi_hi_hi_lo = {c_121,c_120,c_119,c_118,c_117,c_116,c_115,c_114}; // @[wallace_tree.scala 157:17]
  wire  c_123 = wallace_tree_cells_123_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_122 = wallace_tree_cells_122_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_125 = wallace_tree_cells_125_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_124 = wallace_tree_cells_124_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_127 = wallace_tree_cells_127_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_126 = wallace_tree_cells_126_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_130 = wallace_tree_cells_130_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_129 = wallace_tree_cells_129_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire  c_128 = wallace_tree_cells_128_io_o_c; // @[wallace_tree.scala 155:17 161:14]
  wire [16:0] io_o_c_hi_hi_hi = {c_130,c_129,c_128,c_127,c_126,c_125,c_124,c_123,c_122,io_o_c_hi_hi_hi_lo}; // @[wallace_tree.scala 157:17]
  wire [32:0] io_o_c_hi_hi = {io_o_c_hi_hi_hi,c_113,c_112,c_111,c_110,c_109,c_108,c_107,c_106,io_o_c_hi_hi_lo_lo}; // @[wallace_tree.scala 157:17]
  wire [65:0] io_o_c_hi = {io_o_c_hi_hi,io_o_c_hi_lo}; // @[wallace_tree.scala 157:17]
  Wallace_Tree_Cell wallace_tree_cells_0 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_0_io_i_inter_c),
    .io_i_s(wallace_tree_cells_0_io_i_s),
    .io_o_inter_c(wallace_tree_cells_0_io_o_inter_c),
    .io_o_c(wallace_tree_cells_0_io_o_c),
    .io_o_s(wallace_tree_cells_0_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_1 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_1_io_i_inter_c),
    .io_i_s(wallace_tree_cells_1_io_i_s),
    .io_o_inter_c(wallace_tree_cells_1_io_o_inter_c),
    .io_o_c(wallace_tree_cells_1_io_o_c),
    .io_o_s(wallace_tree_cells_1_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_2 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_2_io_i_inter_c),
    .io_i_s(wallace_tree_cells_2_io_i_s),
    .io_o_inter_c(wallace_tree_cells_2_io_o_inter_c),
    .io_o_c(wallace_tree_cells_2_io_o_c),
    .io_o_s(wallace_tree_cells_2_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_3 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_3_io_i_inter_c),
    .io_i_s(wallace_tree_cells_3_io_i_s),
    .io_o_inter_c(wallace_tree_cells_3_io_o_inter_c),
    .io_o_c(wallace_tree_cells_3_io_o_c),
    .io_o_s(wallace_tree_cells_3_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_4 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_4_io_i_inter_c),
    .io_i_s(wallace_tree_cells_4_io_i_s),
    .io_o_inter_c(wallace_tree_cells_4_io_o_inter_c),
    .io_o_c(wallace_tree_cells_4_io_o_c),
    .io_o_s(wallace_tree_cells_4_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_5 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_5_io_i_inter_c),
    .io_i_s(wallace_tree_cells_5_io_i_s),
    .io_o_inter_c(wallace_tree_cells_5_io_o_inter_c),
    .io_o_c(wallace_tree_cells_5_io_o_c),
    .io_o_s(wallace_tree_cells_5_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_6 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_6_io_i_inter_c),
    .io_i_s(wallace_tree_cells_6_io_i_s),
    .io_o_inter_c(wallace_tree_cells_6_io_o_inter_c),
    .io_o_c(wallace_tree_cells_6_io_o_c),
    .io_o_s(wallace_tree_cells_6_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_7 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_7_io_i_inter_c),
    .io_i_s(wallace_tree_cells_7_io_i_s),
    .io_o_inter_c(wallace_tree_cells_7_io_o_inter_c),
    .io_o_c(wallace_tree_cells_7_io_o_c),
    .io_o_s(wallace_tree_cells_7_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_8 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_8_io_i_inter_c),
    .io_i_s(wallace_tree_cells_8_io_i_s),
    .io_o_inter_c(wallace_tree_cells_8_io_o_inter_c),
    .io_o_c(wallace_tree_cells_8_io_o_c),
    .io_o_s(wallace_tree_cells_8_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_9 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_9_io_i_inter_c),
    .io_i_s(wallace_tree_cells_9_io_i_s),
    .io_o_inter_c(wallace_tree_cells_9_io_o_inter_c),
    .io_o_c(wallace_tree_cells_9_io_o_c),
    .io_o_s(wallace_tree_cells_9_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_10 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_10_io_i_inter_c),
    .io_i_s(wallace_tree_cells_10_io_i_s),
    .io_o_inter_c(wallace_tree_cells_10_io_o_inter_c),
    .io_o_c(wallace_tree_cells_10_io_o_c),
    .io_o_s(wallace_tree_cells_10_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_11 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_11_io_i_inter_c),
    .io_i_s(wallace_tree_cells_11_io_i_s),
    .io_o_inter_c(wallace_tree_cells_11_io_o_inter_c),
    .io_o_c(wallace_tree_cells_11_io_o_c),
    .io_o_s(wallace_tree_cells_11_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_12 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_12_io_i_inter_c),
    .io_i_s(wallace_tree_cells_12_io_i_s),
    .io_o_inter_c(wallace_tree_cells_12_io_o_inter_c),
    .io_o_c(wallace_tree_cells_12_io_o_c),
    .io_o_s(wallace_tree_cells_12_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_13 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_13_io_i_inter_c),
    .io_i_s(wallace_tree_cells_13_io_i_s),
    .io_o_inter_c(wallace_tree_cells_13_io_o_inter_c),
    .io_o_c(wallace_tree_cells_13_io_o_c),
    .io_o_s(wallace_tree_cells_13_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_14 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_14_io_i_inter_c),
    .io_i_s(wallace_tree_cells_14_io_i_s),
    .io_o_inter_c(wallace_tree_cells_14_io_o_inter_c),
    .io_o_c(wallace_tree_cells_14_io_o_c),
    .io_o_s(wallace_tree_cells_14_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_15 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_15_io_i_inter_c),
    .io_i_s(wallace_tree_cells_15_io_i_s),
    .io_o_inter_c(wallace_tree_cells_15_io_o_inter_c),
    .io_o_c(wallace_tree_cells_15_io_o_c),
    .io_o_s(wallace_tree_cells_15_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_16 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_16_io_i_inter_c),
    .io_i_s(wallace_tree_cells_16_io_i_s),
    .io_o_inter_c(wallace_tree_cells_16_io_o_inter_c),
    .io_o_c(wallace_tree_cells_16_io_o_c),
    .io_o_s(wallace_tree_cells_16_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_17 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_17_io_i_inter_c),
    .io_i_s(wallace_tree_cells_17_io_i_s),
    .io_o_inter_c(wallace_tree_cells_17_io_o_inter_c),
    .io_o_c(wallace_tree_cells_17_io_o_c),
    .io_o_s(wallace_tree_cells_17_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_18 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_18_io_i_inter_c),
    .io_i_s(wallace_tree_cells_18_io_i_s),
    .io_o_inter_c(wallace_tree_cells_18_io_o_inter_c),
    .io_o_c(wallace_tree_cells_18_io_o_c),
    .io_o_s(wallace_tree_cells_18_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_19 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_19_io_i_inter_c),
    .io_i_s(wallace_tree_cells_19_io_i_s),
    .io_o_inter_c(wallace_tree_cells_19_io_o_inter_c),
    .io_o_c(wallace_tree_cells_19_io_o_c),
    .io_o_s(wallace_tree_cells_19_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_20 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_20_io_i_inter_c),
    .io_i_s(wallace_tree_cells_20_io_i_s),
    .io_o_inter_c(wallace_tree_cells_20_io_o_inter_c),
    .io_o_c(wallace_tree_cells_20_io_o_c),
    .io_o_s(wallace_tree_cells_20_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_21 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_21_io_i_inter_c),
    .io_i_s(wallace_tree_cells_21_io_i_s),
    .io_o_inter_c(wallace_tree_cells_21_io_o_inter_c),
    .io_o_c(wallace_tree_cells_21_io_o_c),
    .io_o_s(wallace_tree_cells_21_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_22 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_22_io_i_inter_c),
    .io_i_s(wallace_tree_cells_22_io_i_s),
    .io_o_inter_c(wallace_tree_cells_22_io_o_inter_c),
    .io_o_c(wallace_tree_cells_22_io_o_c),
    .io_o_s(wallace_tree_cells_22_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_23 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_23_io_i_inter_c),
    .io_i_s(wallace_tree_cells_23_io_i_s),
    .io_o_inter_c(wallace_tree_cells_23_io_o_inter_c),
    .io_o_c(wallace_tree_cells_23_io_o_c),
    .io_o_s(wallace_tree_cells_23_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_24 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_24_io_i_inter_c),
    .io_i_s(wallace_tree_cells_24_io_i_s),
    .io_o_inter_c(wallace_tree_cells_24_io_o_inter_c),
    .io_o_c(wallace_tree_cells_24_io_o_c),
    .io_o_s(wallace_tree_cells_24_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_25 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_25_io_i_inter_c),
    .io_i_s(wallace_tree_cells_25_io_i_s),
    .io_o_inter_c(wallace_tree_cells_25_io_o_inter_c),
    .io_o_c(wallace_tree_cells_25_io_o_c),
    .io_o_s(wallace_tree_cells_25_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_26 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_26_io_i_inter_c),
    .io_i_s(wallace_tree_cells_26_io_i_s),
    .io_o_inter_c(wallace_tree_cells_26_io_o_inter_c),
    .io_o_c(wallace_tree_cells_26_io_o_c),
    .io_o_s(wallace_tree_cells_26_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_27 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_27_io_i_inter_c),
    .io_i_s(wallace_tree_cells_27_io_i_s),
    .io_o_inter_c(wallace_tree_cells_27_io_o_inter_c),
    .io_o_c(wallace_tree_cells_27_io_o_c),
    .io_o_s(wallace_tree_cells_27_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_28 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_28_io_i_inter_c),
    .io_i_s(wallace_tree_cells_28_io_i_s),
    .io_o_inter_c(wallace_tree_cells_28_io_o_inter_c),
    .io_o_c(wallace_tree_cells_28_io_o_c),
    .io_o_s(wallace_tree_cells_28_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_29 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_29_io_i_inter_c),
    .io_i_s(wallace_tree_cells_29_io_i_s),
    .io_o_inter_c(wallace_tree_cells_29_io_o_inter_c),
    .io_o_c(wallace_tree_cells_29_io_o_c),
    .io_o_s(wallace_tree_cells_29_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_30 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_30_io_i_inter_c),
    .io_i_s(wallace_tree_cells_30_io_i_s),
    .io_o_inter_c(wallace_tree_cells_30_io_o_inter_c),
    .io_o_c(wallace_tree_cells_30_io_o_c),
    .io_o_s(wallace_tree_cells_30_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_31 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_31_io_i_inter_c),
    .io_i_s(wallace_tree_cells_31_io_i_s),
    .io_o_inter_c(wallace_tree_cells_31_io_o_inter_c),
    .io_o_c(wallace_tree_cells_31_io_o_c),
    .io_o_s(wallace_tree_cells_31_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_32 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_32_io_i_inter_c),
    .io_i_s(wallace_tree_cells_32_io_i_s),
    .io_o_inter_c(wallace_tree_cells_32_io_o_inter_c),
    .io_o_c(wallace_tree_cells_32_io_o_c),
    .io_o_s(wallace_tree_cells_32_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_33 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_33_io_i_inter_c),
    .io_i_s(wallace_tree_cells_33_io_i_s),
    .io_o_inter_c(wallace_tree_cells_33_io_o_inter_c),
    .io_o_c(wallace_tree_cells_33_io_o_c),
    .io_o_s(wallace_tree_cells_33_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_34 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_34_io_i_inter_c),
    .io_i_s(wallace_tree_cells_34_io_i_s),
    .io_o_inter_c(wallace_tree_cells_34_io_o_inter_c),
    .io_o_c(wallace_tree_cells_34_io_o_c),
    .io_o_s(wallace_tree_cells_34_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_35 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_35_io_i_inter_c),
    .io_i_s(wallace_tree_cells_35_io_i_s),
    .io_o_inter_c(wallace_tree_cells_35_io_o_inter_c),
    .io_o_c(wallace_tree_cells_35_io_o_c),
    .io_o_s(wallace_tree_cells_35_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_36 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_36_io_i_inter_c),
    .io_i_s(wallace_tree_cells_36_io_i_s),
    .io_o_inter_c(wallace_tree_cells_36_io_o_inter_c),
    .io_o_c(wallace_tree_cells_36_io_o_c),
    .io_o_s(wallace_tree_cells_36_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_37 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_37_io_i_inter_c),
    .io_i_s(wallace_tree_cells_37_io_i_s),
    .io_o_inter_c(wallace_tree_cells_37_io_o_inter_c),
    .io_o_c(wallace_tree_cells_37_io_o_c),
    .io_o_s(wallace_tree_cells_37_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_38 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_38_io_i_inter_c),
    .io_i_s(wallace_tree_cells_38_io_i_s),
    .io_o_inter_c(wallace_tree_cells_38_io_o_inter_c),
    .io_o_c(wallace_tree_cells_38_io_o_c),
    .io_o_s(wallace_tree_cells_38_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_39 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_39_io_i_inter_c),
    .io_i_s(wallace_tree_cells_39_io_i_s),
    .io_o_inter_c(wallace_tree_cells_39_io_o_inter_c),
    .io_o_c(wallace_tree_cells_39_io_o_c),
    .io_o_s(wallace_tree_cells_39_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_40 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_40_io_i_inter_c),
    .io_i_s(wallace_tree_cells_40_io_i_s),
    .io_o_inter_c(wallace_tree_cells_40_io_o_inter_c),
    .io_o_c(wallace_tree_cells_40_io_o_c),
    .io_o_s(wallace_tree_cells_40_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_41 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_41_io_i_inter_c),
    .io_i_s(wallace_tree_cells_41_io_i_s),
    .io_o_inter_c(wallace_tree_cells_41_io_o_inter_c),
    .io_o_c(wallace_tree_cells_41_io_o_c),
    .io_o_s(wallace_tree_cells_41_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_42 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_42_io_i_inter_c),
    .io_i_s(wallace_tree_cells_42_io_i_s),
    .io_o_inter_c(wallace_tree_cells_42_io_o_inter_c),
    .io_o_c(wallace_tree_cells_42_io_o_c),
    .io_o_s(wallace_tree_cells_42_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_43 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_43_io_i_inter_c),
    .io_i_s(wallace_tree_cells_43_io_i_s),
    .io_o_inter_c(wallace_tree_cells_43_io_o_inter_c),
    .io_o_c(wallace_tree_cells_43_io_o_c),
    .io_o_s(wallace_tree_cells_43_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_44 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_44_io_i_inter_c),
    .io_i_s(wallace_tree_cells_44_io_i_s),
    .io_o_inter_c(wallace_tree_cells_44_io_o_inter_c),
    .io_o_c(wallace_tree_cells_44_io_o_c),
    .io_o_s(wallace_tree_cells_44_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_45 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_45_io_i_inter_c),
    .io_i_s(wallace_tree_cells_45_io_i_s),
    .io_o_inter_c(wallace_tree_cells_45_io_o_inter_c),
    .io_o_c(wallace_tree_cells_45_io_o_c),
    .io_o_s(wallace_tree_cells_45_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_46 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_46_io_i_inter_c),
    .io_i_s(wallace_tree_cells_46_io_i_s),
    .io_o_inter_c(wallace_tree_cells_46_io_o_inter_c),
    .io_o_c(wallace_tree_cells_46_io_o_c),
    .io_o_s(wallace_tree_cells_46_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_47 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_47_io_i_inter_c),
    .io_i_s(wallace_tree_cells_47_io_i_s),
    .io_o_inter_c(wallace_tree_cells_47_io_o_inter_c),
    .io_o_c(wallace_tree_cells_47_io_o_c),
    .io_o_s(wallace_tree_cells_47_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_48 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_48_io_i_inter_c),
    .io_i_s(wallace_tree_cells_48_io_i_s),
    .io_o_inter_c(wallace_tree_cells_48_io_o_inter_c),
    .io_o_c(wallace_tree_cells_48_io_o_c),
    .io_o_s(wallace_tree_cells_48_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_49 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_49_io_i_inter_c),
    .io_i_s(wallace_tree_cells_49_io_i_s),
    .io_o_inter_c(wallace_tree_cells_49_io_o_inter_c),
    .io_o_c(wallace_tree_cells_49_io_o_c),
    .io_o_s(wallace_tree_cells_49_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_50 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_50_io_i_inter_c),
    .io_i_s(wallace_tree_cells_50_io_i_s),
    .io_o_inter_c(wallace_tree_cells_50_io_o_inter_c),
    .io_o_c(wallace_tree_cells_50_io_o_c),
    .io_o_s(wallace_tree_cells_50_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_51 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_51_io_i_inter_c),
    .io_i_s(wallace_tree_cells_51_io_i_s),
    .io_o_inter_c(wallace_tree_cells_51_io_o_inter_c),
    .io_o_c(wallace_tree_cells_51_io_o_c),
    .io_o_s(wallace_tree_cells_51_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_52 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_52_io_i_inter_c),
    .io_i_s(wallace_tree_cells_52_io_i_s),
    .io_o_inter_c(wallace_tree_cells_52_io_o_inter_c),
    .io_o_c(wallace_tree_cells_52_io_o_c),
    .io_o_s(wallace_tree_cells_52_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_53 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_53_io_i_inter_c),
    .io_i_s(wallace_tree_cells_53_io_i_s),
    .io_o_inter_c(wallace_tree_cells_53_io_o_inter_c),
    .io_o_c(wallace_tree_cells_53_io_o_c),
    .io_o_s(wallace_tree_cells_53_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_54 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_54_io_i_inter_c),
    .io_i_s(wallace_tree_cells_54_io_i_s),
    .io_o_inter_c(wallace_tree_cells_54_io_o_inter_c),
    .io_o_c(wallace_tree_cells_54_io_o_c),
    .io_o_s(wallace_tree_cells_54_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_55 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_55_io_i_inter_c),
    .io_i_s(wallace_tree_cells_55_io_i_s),
    .io_o_inter_c(wallace_tree_cells_55_io_o_inter_c),
    .io_o_c(wallace_tree_cells_55_io_o_c),
    .io_o_s(wallace_tree_cells_55_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_56 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_56_io_i_inter_c),
    .io_i_s(wallace_tree_cells_56_io_i_s),
    .io_o_inter_c(wallace_tree_cells_56_io_o_inter_c),
    .io_o_c(wallace_tree_cells_56_io_o_c),
    .io_o_s(wallace_tree_cells_56_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_57 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_57_io_i_inter_c),
    .io_i_s(wallace_tree_cells_57_io_i_s),
    .io_o_inter_c(wallace_tree_cells_57_io_o_inter_c),
    .io_o_c(wallace_tree_cells_57_io_o_c),
    .io_o_s(wallace_tree_cells_57_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_58 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_58_io_i_inter_c),
    .io_i_s(wallace_tree_cells_58_io_i_s),
    .io_o_inter_c(wallace_tree_cells_58_io_o_inter_c),
    .io_o_c(wallace_tree_cells_58_io_o_c),
    .io_o_s(wallace_tree_cells_58_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_59 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_59_io_i_inter_c),
    .io_i_s(wallace_tree_cells_59_io_i_s),
    .io_o_inter_c(wallace_tree_cells_59_io_o_inter_c),
    .io_o_c(wallace_tree_cells_59_io_o_c),
    .io_o_s(wallace_tree_cells_59_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_60 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_60_io_i_inter_c),
    .io_i_s(wallace_tree_cells_60_io_i_s),
    .io_o_inter_c(wallace_tree_cells_60_io_o_inter_c),
    .io_o_c(wallace_tree_cells_60_io_o_c),
    .io_o_s(wallace_tree_cells_60_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_61 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_61_io_i_inter_c),
    .io_i_s(wallace_tree_cells_61_io_i_s),
    .io_o_inter_c(wallace_tree_cells_61_io_o_inter_c),
    .io_o_c(wallace_tree_cells_61_io_o_c),
    .io_o_s(wallace_tree_cells_61_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_62 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_62_io_i_inter_c),
    .io_i_s(wallace_tree_cells_62_io_i_s),
    .io_o_inter_c(wallace_tree_cells_62_io_o_inter_c),
    .io_o_c(wallace_tree_cells_62_io_o_c),
    .io_o_s(wallace_tree_cells_62_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_63 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_63_io_i_inter_c),
    .io_i_s(wallace_tree_cells_63_io_i_s),
    .io_o_inter_c(wallace_tree_cells_63_io_o_inter_c),
    .io_o_c(wallace_tree_cells_63_io_o_c),
    .io_o_s(wallace_tree_cells_63_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_64 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_64_io_i_inter_c),
    .io_i_s(wallace_tree_cells_64_io_i_s),
    .io_o_inter_c(wallace_tree_cells_64_io_o_inter_c),
    .io_o_c(wallace_tree_cells_64_io_o_c),
    .io_o_s(wallace_tree_cells_64_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_65 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_65_io_i_inter_c),
    .io_i_s(wallace_tree_cells_65_io_i_s),
    .io_o_inter_c(wallace_tree_cells_65_io_o_inter_c),
    .io_o_c(wallace_tree_cells_65_io_o_c),
    .io_o_s(wallace_tree_cells_65_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_66 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_66_io_i_inter_c),
    .io_i_s(wallace_tree_cells_66_io_i_s),
    .io_o_inter_c(wallace_tree_cells_66_io_o_inter_c),
    .io_o_c(wallace_tree_cells_66_io_o_c),
    .io_o_s(wallace_tree_cells_66_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_67 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_67_io_i_inter_c),
    .io_i_s(wallace_tree_cells_67_io_i_s),
    .io_o_inter_c(wallace_tree_cells_67_io_o_inter_c),
    .io_o_c(wallace_tree_cells_67_io_o_c),
    .io_o_s(wallace_tree_cells_67_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_68 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_68_io_i_inter_c),
    .io_i_s(wallace_tree_cells_68_io_i_s),
    .io_o_inter_c(wallace_tree_cells_68_io_o_inter_c),
    .io_o_c(wallace_tree_cells_68_io_o_c),
    .io_o_s(wallace_tree_cells_68_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_69 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_69_io_i_inter_c),
    .io_i_s(wallace_tree_cells_69_io_i_s),
    .io_o_inter_c(wallace_tree_cells_69_io_o_inter_c),
    .io_o_c(wallace_tree_cells_69_io_o_c),
    .io_o_s(wallace_tree_cells_69_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_70 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_70_io_i_inter_c),
    .io_i_s(wallace_tree_cells_70_io_i_s),
    .io_o_inter_c(wallace_tree_cells_70_io_o_inter_c),
    .io_o_c(wallace_tree_cells_70_io_o_c),
    .io_o_s(wallace_tree_cells_70_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_71 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_71_io_i_inter_c),
    .io_i_s(wallace_tree_cells_71_io_i_s),
    .io_o_inter_c(wallace_tree_cells_71_io_o_inter_c),
    .io_o_c(wallace_tree_cells_71_io_o_c),
    .io_o_s(wallace_tree_cells_71_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_72 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_72_io_i_inter_c),
    .io_i_s(wallace_tree_cells_72_io_i_s),
    .io_o_inter_c(wallace_tree_cells_72_io_o_inter_c),
    .io_o_c(wallace_tree_cells_72_io_o_c),
    .io_o_s(wallace_tree_cells_72_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_73 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_73_io_i_inter_c),
    .io_i_s(wallace_tree_cells_73_io_i_s),
    .io_o_inter_c(wallace_tree_cells_73_io_o_inter_c),
    .io_o_c(wallace_tree_cells_73_io_o_c),
    .io_o_s(wallace_tree_cells_73_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_74 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_74_io_i_inter_c),
    .io_i_s(wallace_tree_cells_74_io_i_s),
    .io_o_inter_c(wallace_tree_cells_74_io_o_inter_c),
    .io_o_c(wallace_tree_cells_74_io_o_c),
    .io_o_s(wallace_tree_cells_74_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_75 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_75_io_i_inter_c),
    .io_i_s(wallace_tree_cells_75_io_i_s),
    .io_o_inter_c(wallace_tree_cells_75_io_o_inter_c),
    .io_o_c(wallace_tree_cells_75_io_o_c),
    .io_o_s(wallace_tree_cells_75_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_76 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_76_io_i_inter_c),
    .io_i_s(wallace_tree_cells_76_io_i_s),
    .io_o_inter_c(wallace_tree_cells_76_io_o_inter_c),
    .io_o_c(wallace_tree_cells_76_io_o_c),
    .io_o_s(wallace_tree_cells_76_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_77 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_77_io_i_inter_c),
    .io_i_s(wallace_tree_cells_77_io_i_s),
    .io_o_inter_c(wallace_tree_cells_77_io_o_inter_c),
    .io_o_c(wallace_tree_cells_77_io_o_c),
    .io_o_s(wallace_tree_cells_77_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_78 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_78_io_i_inter_c),
    .io_i_s(wallace_tree_cells_78_io_i_s),
    .io_o_inter_c(wallace_tree_cells_78_io_o_inter_c),
    .io_o_c(wallace_tree_cells_78_io_o_c),
    .io_o_s(wallace_tree_cells_78_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_79 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_79_io_i_inter_c),
    .io_i_s(wallace_tree_cells_79_io_i_s),
    .io_o_inter_c(wallace_tree_cells_79_io_o_inter_c),
    .io_o_c(wallace_tree_cells_79_io_o_c),
    .io_o_s(wallace_tree_cells_79_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_80 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_80_io_i_inter_c),
    .io_i_s(wallace_tree_cells_80_io_i_s),
    .io_o_inter_c(wallace_tree_cells_80_io_o_inter_c),
    .io_o_c(wallace_tree_cells_80_io_o_c),
    .io_o_s(wallace_tree_cells_80_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_81 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_81_io_i_inter_c),
    .io_i_s(wallace_tree_cells_81_io_i_s),
    .io_o_inter_c(wallace_tree_cells_81_io_o_inter_c),
    .io_o_c(wallace_tree_cells_81_io_o_c),
    .io_o_s(wallace_tree_cells_81_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_82 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_82_io_i_inter_c),
    .io_i_s(wallace_tree_cells_82_io_i_s),
    .io_o_inter_c(wallace_tree_cells_82_io_o_inter_c),
    .io_o_c(wallace_tree_cells_82_io_o_c),
    .io_o_s(wallace_tree_cells_82_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_83 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_83_io_i_inter_c),
    .io_i_s(wallace_tree_cells_83_io_i_s),
    .io_o_inter_c(wallace_tree_cells_83_io_o_inter_c),
    .io_o_c(wallace_tree_cells_83_io_o_c),
    .io_o_s(wallace_tree_cells_83_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_84 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_84_io_i_inter_c),
    .io_i_s(wallace_tree_cells_84_io_i_s),
    .io_o_inter_c(wallace_tree_cells_84_io_o_inter_c),
    .io_o_c(wallace_tree_cells_84_io_o_c),
    .io_o_s(wallace_tree_cells_84_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_85 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_85_io_i_inter_c),
    .io_i_s(wallace_tree_cells_85_io_i_s),
    .io_o_inter_c(wallace_tree_cells_85_io_o_inter_c),
    .io_o_c(wallace_tree_cells_85_io_o_c),
    .io_o_s(wallace_tree_cells_85_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_86 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_86_io_i_inter_c),
    .io_i_s(wallace_tree_cells_86_io_i_s),
    .io_o_inter_c(wallace_tree_cells_86_io_o_inter_c),
    .io_o_c(wallace_tree_cells_86_io_o_c),
    .io_o_s(wallace_tree_cells_86_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_87 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_87_io_i_inter_c),
    .io_i_s(wallace_tree_cells_87_io_i_s),
    .io_o_inter_c(wallace_tree_cells_87_io_o_inter_c),
    .io_o_c(wallace_tree_cells_87_io_o_c),
    .io_o_s(wallace_tree_cells_87_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_88 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_88_io_i_inter_c),
    .io_i_s(wallace_tree_cells_88_io_i_s),
    .io_o_inter_c(wallace_tree_cells_88_io_o_inter_c),
    .io_o_c(wallace_tree_cells_88_io_o_c),
    .io_o_s(wallace_tree_cells_88_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_89 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_89_io_i_inter_c),
    .io_i_s(wallace_tree_cells_89_io_i_s),
    .io_o_inter_c(wallace_tree_cells_89_io_o_inter_c),
    .io_o_c(wallace_tree_cells_89_io_o_c),
    .io_o_s(wallace_tree_cells_89_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_90 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_90_io_i_inter_c),
    .io_i_s(wallace_tree_cells_90_io_i_s),
    .io_o_inter_c(wallace_tree_cells_90_io_o_inter_c),
    .io_o_c(wallace_tree_cells_90_io_o_c),
    .io_o_s(wallace_tree_cells_90_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_91 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_91_io_i_inter_c),
    .io_i_s(wallace_tree_cells_91_io_i_s),
    .io_o_inter_c(wallace_tree_cells_91_io_o_inter_c),
    .io_o_c(wallace_tree_cells_91_io_o_c),
    .io_o_s(wallace_tree_cells_91_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_92 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_92_io_i_inter_c),
    .io_i_s(wallace_tree_cells_92_io_i_s),
    .io_o_inter_c(wallace_tree_cells_92_io_o_inter_c),
    .io_o_c(wallace_tree_cells_92_io_o_c),
    .io_o_s(wallace_tree_cells_92_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_93 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_93_io_i_inter_c),
    .io_i_s(wallace_tree_cells_93_io_i_s),
    .io_o_inter_c(wallace_tree_cells_93_io_o_inter_c),
    .io_o_c(wallace_tree_cells_93_io_o_c),
    .io_o_s(wallace_tree_cells_93_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_94 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_94_io_i_inter_c),
    .io_i_s(wallace_tree_cells_94_io_i_s),
    .io_o_inter_c(wallace_tree_cells_94_io_o_inter_c),
    .io_o_c(wallace_tree_cells_94_io_o_c),
    .io_o_s(wallace_tree_cells_94_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_95 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_95_io_i_inter_c),
    .io_i_s(wallace_tree_cells_95_io_i_s),
    .io_o_inter_c(wallace_tree_cells_95_io_o_inter_c),
    .io_o_c(wallace_tree_cells_95_io_o_c),
    .io_o_s(wallace_tree_cells_95_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_96 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_96_io_i_inter_c),
    .io_i_s(wallace_tree_cells_96_io_i_s),
    .io_o_inter_c(wallace_tree_cells_96_io_o_inter_c),
    .io_o_c(wallace_tree_cells_96_io_o_c),
    .io_o_s(wallace_tree_cells_96_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_97 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_97_io_i_inter_c),
    .io_i_s(wallace_tree_cells_97_io_i_s),
    .io_o_inter_c(wallace_tree_cells_97_io_o_inter_c),
    .io_o_c(wallace_tree_cells_97_io_o_c),
    .io_o_s(wallace_tree_cells_97_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_98 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_98_io_i_inter_c),
    .io_i_s(wallace_tree_cells_98_io_i_s),
    .io_o_inter_c(wallace_tree_cells_98_io_o_inter_c),
    .io_o_c(wallace_tree_cells_98_io_o_c),
    .io_o_s(wallace_tree_cells_98_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_99 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_99_io_i_inter_c),
    .io_i_s(wallace_tree_cells_99_io_i_s),
    .io_o_inter_c(wallace_tree_cells_99_io_o_inter_c),
    .io_o_c(wallace_tree_cells_99_io_o_c),
    .io_o_s(wallace_tree_cells_99_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_100 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_100_io_i_inter_c),
    .io_i_s(wallace_tree_cells_100_io_i_s),
    .io_o_inter_c(wallace_tree_cells_100_io_o_inter_c),
    .io_o_c(wallace_tree_cells_100_io_o_c),
    .io_o_s(wallace_tree_cells_100_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_101 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_101_io_i_inter_c),
    .io_i_s(wallace_tree_cells_101_io_i_s),
    .io_o_inter_c(wallace_tree_cells_101_io_o_inter_c),
    .io_o_c(wallace_tree_cells_101_io_o_c),
    .io_o_s(wallace_tree_cells_101_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_102 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_102_io_i_inter_c),
    .io_i_s(wallace_tree_cells_102_io_i_s),
    .io_o_inter_c(wallace_tree_cells_102_io_o_inter_c),
    .io_o_c(wallace_tree_cells_102_io_o_c),
    .io_o_s(wallace_tree_cells_102_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_103 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_103_io_i_inter_c),
    .io_i_s(wallace_tree_cells_103_io_i_s),
    .io_o_inter_c(wallace_tree_cells_103_io_o_inter_c),
    .io_o_c(wallace_tree_cells_103_io_o_c),
    .io_o_s(wallace_tree_cells_103_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_104 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_104_io_i_inter_c),
    .io_i_s(wallace_tree_cells_104_io_i_s),
    .io_o_inter_c(wallace_tree_cells_104_io_o_inter_c),
    .io_o_c(wallace_tree_cells_104_io_o_c),
    .io_o_s(wallace_tree_cells_104_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_105 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_105_io_i_inter_c),
    .io_i_s(wallace_tree_cells_105_io_i_s),
    .io_o_inter_c(wallace_tree_cells_105_io_o_inter_c),
    .io_o_c(wallace_tree_cells_105_io_o_c),
    .io_o_s(wallace_tree_cells_105_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_106 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_106_io_i_inter_c),
    .io_i_s(wallace_tree_cells_106_io_i_s),
    .io_o_inter_c(wallace_tree_cells_106_io_o_inter_c),
    .io_o_c(wallace_tree_cells_106_io_o_c),
    .io_o_s(wallace_tree_cells_106_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_107 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_107_io_i_inter_c),
    .io_i_s(wallace_tree_cells_107_io_i_s),
    .io_o_inter_c(wallace_tree_cells_107_io_o_inter_c),
    .io_o_c(wallace_tree_cells_107_io_o_c),
    .io_o_s(wallace_tree_cells_107_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_108 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_108_io_i_inter_c),
    .io_i_s(wallace_tree_cells_108_io_i_s),
    .io_o_inter_c(wallace_tree_cells_108_io_o_inter_c),
    .io_o_c(wallace_tree_cells_108_io_o_c),
    .io_o_s(wallace_tree_cells_108_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_109 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_109_io_i_inter_c),
    .io_i_s(wallace_tree_cells_109_io_i_s),
    .io_o_inter_c(wallace_tree_cells_109_io_o_inter_c),
    .io_o_c(wallace_tree_cells_109_io_o_c),
    .io_o_s(wallace_tree_cells_109_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_110 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_110_io_i_inter_c),
    .io_i_s(wallace_tree_cells_110_io_i_s),
    .io_o_inter_c(wallace_tree_cells_110_io_o_inter_c),
    .io_o_c(wallace_tree_cells_110_io_o_c),
    .io_o_s(wallace_tree_cells_110_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_111 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_111_io_i_inter_c),
    .io_i_s(wallace_tree_cells_111_io_i_s),
    .io_o_inter_c(wallace_tree_cells_111_io_o_inter_c),
    .io_o_c(wallace_tree_cells_111_io_o_c),
    .io_o_s(wallace_tree_cells_111_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_112 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_112_io_i_inter_c),
    .io_i_s(wallace_tree_cells_112_io_i_s),
    .io_o_inter_c(wallace_tree_cells_112_io_o_inter_c),
    .io_o_c(wallace_tree_cells_112_io_o_c),
    .io_o_s(wallace_tree_cells_112_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_113 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_113_io_i_inter_c),
    .io_i_s(wallace_tree_cells_113_io_i_s),
    .io_o_inter_c(wallace_tree_cells_113_io_o_inter_c),
    .io_o_c(wallace_tree_cells_113_io_o_c),
    .io_o_s(wallace_tree_cells_113_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_114 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_114_io_i_inter_c),
    .io_i_s(wallace_tree_cells_114_io_i_s),
    .io_o_inter_c(wallace_tree_cells_114_io_o_inter_c),
    .io_o_c(wallace_tree_cells_114_io_o_c),
    .io_o_s(wallace_tree_cells_114_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_115 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_115_io_i_inter_c),
    .io_i_s(wallace_tree_cells_115_io_i_s),
    .io_o_inter_c(wallace_tree_cells_115_io_o_inter_c),
    .io_o_c(wallace_tree_cells_115_io_o_c),
    .io_o_s(wallace_tree_cells_115_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_116 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_116_io_i_inter_c),
    .io_i_s(wallace_tree_cells_116_io_i_s),
    .io_o_inter_c(wallace_tree_cells_116_io_o_inter_c),
    .io_o_c(wallace_tree_cells_116_io_o_c),
    .io_o_s(wallace_tree_cells_116_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_117 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_117_io_i_inter_c),
    .io_i_s(wallace_tree_cells_117_io_i_s),
    .io_o_inter_c(wallace_tree_cells_117_io_o_inter_c),
    .io_o_c(wallace_tree_cells_117_io_o_c),
    .io_o_s(wallace_tree_cells_117_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_118 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_118_io_i_inter_c),
    .io_i_s(wallace_tree_cells_118_io_i_s),
    .io_o_inter_c(wallace_tree_cells_118_io_o_inter_c),
    .io_o_c(wallace_tree_cells_118_io_o_c),
    .io_o_s(wallace_tree_cells_118_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_119 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_119_io_i_inter_c),
    .io_i_s(wallace_tree_cells_119_io_i_s),
    .io_o_inter_c(wallace_tree_cells_119_io_o_inter_c),
    .io_o_c(wallace_tree_cells_119_io_o_c),
    .io_o_s(wallace_tree_cells_119_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_120 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_120_io_i_inter_c),
    .io_i_s(wallace_tree_cells_120_io_i_s),
    .io_o_inter_c(wallace_tree_cells_120_io_o_inter_c),
    .io_o_c(wallace_tree_cells_120_io_o_c),
    .io_o_s(wallace_tree_cells_120_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_121 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_121_io_i_inter_c),
    .io_i_s(wallace_tree_cells_121_io_i_s),
    .io_o_inter_c(wallace_tree_cells_121_io_o_inter_c),
    .io_o_c(wallace_tree_cells_121_io_o_c),
    .io_o_s(wallace_tree_cells_121_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_122 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_122_io_i_inter_c),
    .io_i_s(wallace_tree_cells_122_io_i_s),
    .io_o_inter_c(wallace_tree_cells_122_io_o_inter_c),
    .io_o_c(wallace_tree_cells_122_io_o_c),
    .io_o_s(wallace_tree_cells_122_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_123 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_123_io_i_inter_c),
    .io_i_s(wallace_tree_cells_123_io_i_s),
    .io_o_inter_c(wallace_tree_cells_123_io_o_inter_c),
    .io_o_c(wallace_tree_cells_123_io_o_c),
    .io_o_s(wallace_tree_cells_123_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_124 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_124_io_i_inter_c),
    .io_i_s(wallace_tree_cells_124_io_i_s),
    .io_o_inter_c(wallace_tree_cells_124_io_o_inter_c),
    .io_o_c(wallace_tree_cells_124_io_o_c),
    .io_o_s(wallace_tree_cells_124_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_125 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_125_io_i_inter_c),
    .io_i_s(wallace_tree_cells_125_io_i_s),
    .io_o_inter_c(wallace_tree_cells_125_io_o_inter_c),
    .io_o_c(wallace_tree_cells_125_io_o_c),
    .io_o_s(wallace_tree_cells_125_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_126 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_126_io_i_inter_c),
    .io_i_s(wallace_tree_cells_126_io_i_s),
    .io_o_inter_c(wallace_tree_cells_126_io_o_inter_c),
    .io_o_c(wallace_tree_cells_126_io_o_c),
    .io_o_s(wallace_tree_cells_126_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_127 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_127_io_i_inter_c),
    .io_i_s(wallace_tree_cells_127_io_i_s),
    .io_o_inter_c(wallace_tree_cells_127_io_o_inter_c),
    .io_o_c(wallace_tree_cells_127_io_o_c),
    .io_o_s(wallace_tree_cells_127_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_128 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_128_io_i_inter_c),
    .io_i_s(wallace_tree_cells_128_io_i_s),
    .io_o_inter_c(wallace_tree_cells_128_io_o_inter_c),
    .io_o_c(wallace_tree_cells_128_io_o_c),
    .io_o_s(wallace_tree_cells_128_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_129 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_129_io_i_inter_c),
    .io_i_s(wallace_tree_cells_129_io_i_s),
    .io_o_inter_c(wallace_tree_cells_129_io_o_inter_c),
    .io_o_c(wallace_tree_cells_129_io_o_c),
    .io_o_s(wallace_tree_cells_129_io_o_s)
  );
  Wallace_Tree_Cell wallace_tree_cells_130 ( // @[wallace_tree.scala 137:50]
    .io_i_inter_c(wallace_tree_cells_130_io_i_inter_c),
    .io_i_s(wallace_tree_cells_130_io_i_s),
    .io_o_inter_c(wallace_tree_cells_130_io_o_inter_c),
    .io_o_c(wallace_tree_cells_130_io_o_c),
    .io_o_s(wallace_tree_cells_130_io_o_s)
  );
  assign io_o_s = {io_o_s_hi,io_o_s_lo}; // @[wallace_tree.scala 156:17]
  assign io_o_c = {io_o_c_hi,io_o_c_lo}; // @[wallace_tree.scala 157:17]
  assign wallace_tree_cells_0_io_i_inter_c = 19'h0; // @[wallace_tree.scala 150:40]
  assign wallace_tree_cells_0_io_i_s = {wallace_tree_cells_0_io_i_s_hi,wallace_tree_cells_0_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_1_io_i_inter_c = wallace_tree_cells_0_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_1_io_i_s = {wallace_tree_cells_1_io_i_s_hi,wallace_tree_cells_1_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_2_io_i_inter_c = wallace_tree_cells_1_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_2_io_i_s = {wallace_tree_cells_2_io_i_s_hi,wallace_tree_cells_2_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_3_io_i_inter_c = wallace_tree_cells_2_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_3_io_i_s = {wallace_tree_cells_3_io_i_s_hi,wallace_tree_cells_3_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_4_io_i_inter_c = wallace_tree_cells_3_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_4_io_i_s = {wallace_tree_cells_4_io_i_s_hi,wallace_tree_cells_4_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_5_io_i_inter_c = wallace_tree_cells_4_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_5_io_i_s = {wallace_tree_cells_5_io_i_s_hi,wallace_tree_cells_5_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_6_io_i_inter_c = wallace_tree_cells_5_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_6_io_i_s = {wallace_tree_cells_6_io_i_s_hi,wallace_tree_cells_6_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_7_io_i_inter_c = wallace_tree_cells_6_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_7_io_i_s = {wallace_tree_cells_7_io_i_s_hi,wallace_tree_cells_7_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_8_io_i_inter_c = wallace_tree_cells_7_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_8_io_i_s = {wallace_tree_cells_8_io_i_s_hi,wallace_tree_cells_8_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_9_io_i_inter_c = wallace_tree_cells_8_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_9_io_i_s = {wallace_tree_cells_9_io_i_s_hi,wallace_tree_cells_9_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_10_io_i_inter_c = wallace_tree_cells_9_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_10_io_i_s = {wallace_tree_cells_10_io_i_s_hi,wallace_tree_cells_10_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_11_io_i_inter_c = wallace_tree_cells_10_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_11_io_i_s = {wallace_tree_cells_11_io_i_s_hi,wallace_tree_cells_11_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_12_io_i_inter_c = wallace_tree_cells_11_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_12_io_i_s = {wallace_tree_cells_12_io_i_s_hi,wallace_tree_cells_12_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_13_io_i_inter_c = wallace_tree_cells_12_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_13_io_i_s = {wallace_tree_cells_13_io_i_s_hi,wallace_tree_cells_13_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_14_io_i_inter_c = wallace_tree_cells_13_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_14_io_i_s = {wallace_tree_cells_14_io_i_s_hi,wallace_tree_cells_14_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_15_io_i_inter_c = wallace_tree_cells_14_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_15_io_i_s = {wallace_tree_cells_15_io_i_s_hi,wallace_tree_cells_15_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_16_io_i_inter_c = wallace_tree_cells_15_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_16_io_i_s = {wallace_tree_cells_16_io_i_s_hi,wallace_tree_cells_16_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_17_io_i_inter_c = wallace_tree_cells_16_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_17_io_i_s = {wallace_tree_cells_17_io_i_s_hi,wallace_tree_cells_17_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_18_io_i_inter_c = wallace_tree_cells_17_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_18_io_i_s = {wallace_tree_cells_18_io_i_s_hi,wallace_tree_cells_18_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_19_io_i_inter_c = wallace_tree_cells_18_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_19_io_i_s = {wallace_tree_cells_19_io_i_s_hi,wallace_tree_cells_19_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_20_io_i_inter_c = wallace_tree_cells_19_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_20_io_i_s = {wallace_tree_cells_20_io_i_s_hi,wallace_tree_cells_20_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_21_io_i_inter_c = wallace_tree_cells_20_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_21_io_i_s = {wallace_tree_cells_21_io_i_s_hi,wallace_tree_cells_21_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_22_io_i_inter_c = wallace_tree_cells_21_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_22_io_i_s = {wallace_tree_cells_22_io_i_s_hi,wallace_tree_cells_22_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_23_io_i_inter_c = wallace_tree_cells_22_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_23_io_i_s = {wallace_tree_cells_23_io_i_s_hi,wallace_tree_cells_23_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_24_io_i_inter_c = wallace_tree_cells_23_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_24_io_i_s = {wallace_tree_cells_24_io_i_s_hi,wallace_tree_cells_24_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_25_io_i_inter_c = wallace_tree_cells_24_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_25_io_i_s = {wallace_tree_cells_25_io_i_s_hi,wallace_tree_cells_25_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_26_io_i_inter_c = wallace_tree_cells_25_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_26_io_i_s = {wallace_tree_cells_26_io_i_s_hi,wallace_tree_cells_26_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_27_io_i_inter_c = wallace_tree_cells_26_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_27_io_i_s = {wallace_tree_cells_27_io_i_s_hi,wallace_tree_cells_27_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_28_io_i_inter_c = wallace_tree_cells_27_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_28_io_i_s = {wallace_tree_cells_28_io_i_s_hi,wallace_tree_cells_28_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_29_io_i_inter_c = wallace_tree_cells_28_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_29_io_i_s = {wallace_tree_cells_29_io_i_s_hi,wallace_tree_cells_29_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_30_io_i_inter_c = wallace_tree_cells_29_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_30_io_i_s = {wallace_tree_cells_30_io_i_s_hi,wallace_tree_cells_30_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_31_io_i_inter_c = wallace_tree_cells_30_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_31_io_i_s = {wallace_tree_cells_31_io_i_s_hi,wallace_tree_cells_31_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_32_io_i_inter_c = wallace_tree_cells_31_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_32_io_i_s = {wallace_tree_cells_32_io_i_s_hi,wallace_tree_cells_32_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_33_io_i_inter_c = wallace_tree_cells_32_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_33_io_i_s = {wallace_tree_cells_33_io_i_s_hi,wallace_tree_cells_33_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_34_io_i_inter_c = wallace_tree_cells_33_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_34_io_i_s = {wallace_tree_cells_34_io_i_s_hi,wallace_tree_cells_34_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_35_io_i_inter_c = wallace_tree_cells_34_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_35_io_i_s = {wallace_tree_cells_35_io_i_s_hi,wallace_tree_cells_35_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_36_io_i_inter_c = wallace_tree_cells_35_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_36_io_i_s = {wallace_tree_cells_36_io_i_s_hi,wallace_tree_cells_36_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_37_io_i_inter_c = wallace_tree_cells_36_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_37_io_i_s = {wallace_tree_cells_37_io_i_s_hi,wallace_tree_cells_37_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_38_io_i_inter_c = wallace_tree_cells_37_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_38_io_i_s = {wallace_tree_cells_38_io_i_s_hi,wallace_tree_cells_38_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_39_io_i_inter_c = wallace_tree_cells_38_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_39_io_i_s = {wallace_tree_cells_39_io_i_s_hi,wallace_tree_cells_39_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_40_io_i_inter_c = wallace_tree_cells_39_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_40_io_i_s = {wallace_tree_cells_40_io_i_s_hi,wallace_tree_cells_40_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_41_io_i_inter_c = wallace_tree_cells_40_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_41_io_i_s = {wallace_tree_cells_41_io_i_s_hi,wallace_tree_cells_41_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_42_io_i_inter_c = wallace_tree_cells_41_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_42_io_i_s = {wallace_tree_cells_42_io_i_s_hi,wallace_tree_cells_42_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_43_io_i_inter_c = wallace_tree_cells_42_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_43_io_i_s = {wallace_tree_cells_43_io_i_s_hi,wallace_tree_cells_43_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_44_io_i_inter_c = wallace_tree_cells_43_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_44_io_i_s = {wallace_tree_cells_44_io_i_s_hi,wallace_tree_cells_44_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_45_io_i_inter_c = wallace_tree_cells_44_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_45_io_i_s = {wallace_tree_cells_45_io_i_s_hi,wallace_tree_cells_45_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_46_io_i_inter_c = wallace_tree_cells_45_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_46_io_i_s = {wallace_tree_cells_46_io_i_s_hi,wallace_tree_cells_46_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_47_io_i_inter_c = wallace_tree_cells_46_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_47_io_i_s = {wallace_tree_cells_47_io_i_s_hi,wallace_tree_cells_47_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_48_io_i_inter_c = wallace_tree_cells_47_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_48_io_i_s = {wallace_tree_cells_48_io_i_s_hi,wallace_tree_cells_48_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_49_io_i_inter_c = wallace_tree_cells_48_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_49_io_i_s = {wallace_tree_cells_49_io_i_s_hi,wallace_tree_cells_49_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_50_io_i_inter_c = wallace_tree_cells_49_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_50_io_i_s = {wallace_tree_cells_50_io_i_s_hi,wallace_tree_cells_50_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_51_io_i_inter_c = wallace_tree_cells_50_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_51_io_i_s = {wallace_tree_cells_51_io_i_s_hi,wallace_tree_cells_51_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_52_io_i_inter_c = wallace_tree_cells_51_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_52_io_i_s = {wallace_tree_cells_52_io_i_s_hi,wallace_tree_cells_52_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_53_io_i_inter_c = wallace_tree_cells_52_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_53_io_i_s = {wallace_tree_cells_53_io_i_s_hi,wallace_tree_cells_53_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_54_io_i_inter_c = wallace_tree_cells_53_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_54_io_i_s = {wallace_tree_cells_54_io_i_s_hi,wallace_tree_cells_54_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_55_io_i_inter_c = wallace_tree_cells_54_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_55_io_i_s = {wallace_tree_cells_55_io_i_s_hi,wallace_tree_cells_55_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_56_io_i_inter_c = wallace_tree_cells_55_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_56_io_i_s = {wallace_tree_cells_56_io_i_s_hi,wallace_tree_cells_56_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_57_io_i_inter_c = wallace_tree_cells_56_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_57_io_i_s = {wallace_tree_cells_57_io_i_s_hi,wallace_tree_cells_57_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_58_io_i_inter_c = wallace_tree_cells_57_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_58_io_i_s = {wallace_tree_cells_58_io_i_s_hi,wallace_tree_cells_58_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_59_io_i_inter_c = wallace_tree_cells_58_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_59_io_i_s = {wallace_tree_cells_59_io_i_s_hi,wallace_tree_cells_59_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_60_io_i_inter_c = wallace_tree_cells_59_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_60_io_i_s = {wallace_tree_cells_60_io_i_s_hi,wallace_tree_cells_60_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_61_io_i_inter_c = wallace_tree_cells_60_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_61_io_i_s = {wallace_tree_cells_61_io_i_s_hi,wallace_tree_cells_61_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_62_io_i_inter_c = wallace_tree_cells_61_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_62_io_i_s = {wallace_tree_cells_62_io_i_s_hi,wallace_tree_cells_62_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_63_io_i_inter_c = wallace_tree_cells_62_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_63_io_i_s = {wallace_tree_cells_63_io_i_s_hi,wallace_tree_cells_63_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_64_io_i_inter_c = wallace_tree_cells_63_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_64_io_i_s = {wallace_tree_cells_64_io_i_s_hi,wallace_tree_cells_64_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_65_io_i_inter_c = wallace_tree_cells_64_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_65_io_i_s = {wallace_tree_cells_65_io_i_s_hi,wallace_tree_cells_65_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_66_io_i_inter_c = wallace_tree_cells_65_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_66_io_i_s = {wallace_tree_cells_66_io_i_s_hi,wallace_tree_cells_66_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_67_io_i_inter_c = wallace_tree_cells_66_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_67_io_i_s = {wallace_tree_cells_67_io_i_s_hi,wallace_tree_cells_67_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_68_io_i_inter_c = wallace_tree_cells_67_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_68_io_i_s = {wallace_tree_cells_68_io_i_s_hi,wallace_tree_cells_68_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_69_io_i_inter_c = wallace_tree_cells_68_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_69_io_i_s = {wallace_tree_cells_69_io_i_s_hi,wallace_tree_cells_69_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_70_io_i_inter_c = wallace_tree_cells_69_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_70_io_i_s = {wallace_tree_cells_70_io_i_s_hi,wallace_tree_cells_70_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_71_io_i_inter_c = wallace_tree_cells_70_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_71_io_i_s = {wallace_tree_cells_71_io_i_s_hi,wallace_tree_cells_71_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_72_io_i_inter_c = wallace_tree_cells_71_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_72_io_i_s = {wallace_tree_cells_72_io_i_s_hi,wallace_tree_cells_72_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_73_io_i_inter_c = wallace_tree_cells_72_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_73_io_i_s = {wallace_tree_cells_73_io_i_s_hi,wallace_tree_cells_73_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_74_io_i_inter_c = wallace_tree_cells_73_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_74_io_i_s = {wallace_tree_cells_74_io_i_s_hi,wallace_tree_cells_74_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_75_io_i_inter_c = wallace_tree_cells_74_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_75_io_i_s = {wallace_tree_cells_75_io_i_s_hi,wallace_tree_cells_75_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_76_io_i_inter_c = wallace_tree_cells_75_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_76_io_i_s = {wallace_tree_cells_76_io_i_s_hi,wallace_tree_cells_76_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_77_io_i_inter_c = wallace_tree_cells_76_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_77_io_i_s = {wallace_tree_cells_77_io_i_s_hi,wallace_tree_cells_77_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_78_io_i_inter_c = wallace_tree_cells_77_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_78_io_i_s = {wallace_tree_cells_78_io_i_s_hi,wallace_tree_cells_78_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_79_io_i_inter_c = wallace_tree_cells_78_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_79_io_i_s = {wallace_tree_cells_79_io_i_s_hi,wallace_tree_cells_79_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_80_io_i_inter_c = wallace_tree_cells_79_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_80_io_i_s = {wallace_tree_cells_80_io_i_s_hi,wallace_tree_cells_80_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_81_io_i_inter_c = wallace_tree_cells_80_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_81_io_i_s = {wallace_tree_cells_81_io_i_s_hi,wallace_tree_cells_81_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_82_io_i_inter_c = wallace_tree_cells_81_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_82_io_i_s = {wallace_tree_cells_82_io_i_s_hi,wallace_tree_cells_82_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_83_io_i_inter_c = wallace_tree_cells_82_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_83_io_i_s = {wallace_tree_cells_83_io_i_s_hi,wallace_tree_cells_83_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_84_io_i_inter_c = wallace_tree_cells_83_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_84_io_i_s = {wallace_tree_cells_84_io_i_s_hi,wallace_tree_cells_84_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_85_io_i_inter_c = wallace_tree_cells_84_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_85_io_i_s = {wallace_tree_cells_85_io_i_s_hi,wallace_tree_cells_85_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_86_io_i_inter_c = wallace_tree_cells_85_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_86_io_i_s = {wallace_tree_cells_86_io_i_s_hi,wallace_tree_cells_86_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_87_io_i_inter_c = wallace_tree_cells_86_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_87_io_i_s = {wallace_tree_cells_87_io_i_s_hi,wallace_tree_cells_87_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_88_io_i_inter_c = wallace_tree_cells_87_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_88_io_i_s = {wallace_tree_cells_88_io_i_s_hi,wallace_tree_cells_88_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_89_io_i_inter_c = wallace_tree_cells_88_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_89_io_i_s = {wallace_tree_cells_89_io_i_s_hi,wallace_tree_cells_89_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_90_io_i_inter_c = wallace_tree_cells_89_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_90_io_i_s = {wallace_tree_cells_90_io_i_s_hi,wallace_tree_cells_90_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_91_io_i_inter_c = wallace_tree_cells_90_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_91_io_i_s = {wallace_tree_cells_91_io_i_s_hi,wallace_tree_cells_91_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_92_io_i_inter_c = wallace_tree_cells_91_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_92_io_i_s = {wallace_tree_cells_92_io_i_s_hi,wallace_tree_cells_92_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_93_io_i_inter_c = wallace_tree_cells_92_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_93_io_i_s = {wallace_tree_cells_93_io_i_s_hi,wallace_tree_cells_93_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_94_io_i_inter_c = wallace_tree_cells_93_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_94_io_i_s = {wallace_tree_cells_94_io_i_s_hi,wallace_tree_cells_94_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_95_io_i_inter_c = wallace_tree_cells_94_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_95_io_i_s = {wallace_tree_cells_95_io_i_s_hi,wallace_tree_cells_95_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_96_io_i_inter_c = wallace_tree_cells_95_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_96_io_i_s = {wallace_tree_cells_96_io_i_s_hi,wallace_tree_cells_96_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_97_io_i_inter_c = wallace_tree_cells_96_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_97_io_i_s = {wallace_tree_cells_97_io_i_s_hi,wallace_tree_cells_97_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_98_io_i_inter_c = wallace_tree_cells_97_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_98_io_i_s = {wallace_tree_cells_98_io_i_s_hi,wallace_tree_cells_98_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_99_io_i_inter_c = wallace_tree_cells_98_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_99_io_i_s = {wallace_tree_cells_99_io_i_s_hi,wallace_tree_cells_99_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_100_io_i_inter_c = wallace_tree_cells_99_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_100_io_i_s = {wallace_tree_cells_100_io_i_s_hi,wallace_tree_cells_100_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_101_io_i_inter_c = wallace_tree_cells_100_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_101_io_i_s = {wallace_tree_cells_101_io_i_s_hi,wallace_tree_cells_101_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_102_io_i_inter_c = wallace_tree_cells_101_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_102_io_i_s = {wallace_tree_cells_102_io_i_s_hi,wallace_tree_cells_102_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_103_io_i_inter_c = wallace_tree_cells_102_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_103_io_i_s = {wallace_tree_cells_103_io_i_s_hi,wallace_tree_cells_103_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_104_io_i_inter_c = wallace_tree_cells_103_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_104_io_i_s = {wallace_tree_cells_104_io_i_s_hi,wallace_tree_cells_104_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_105_io_i_inter_c = wallace_tree_cells_104_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_105_io_i_s = {wallace_tree_cells_105_io_i_s_hi,wallace_tree_cells_105_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_106_io_i_inter_c = wallace_tree_cells_105_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_106_io_i_s = {wallace_tree_cells_106_io_i_s_hi,wallace_tree_cells_106_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_107_io_i_inter_c = wallace_tree_cells_106_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_107_io_i_s = {wallace_tree_cells_107_io_i_s_hi,wallace_tree_cells_107_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_108_io_i_inter_c = wallace_tree_cells_107_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_108_io_i_s = {wallace_tree_cells_108_io_i_s_hi,wallace_tree_cells_108_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_109_io_i_inter_c = wallace_tree_cells_108_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_109_io_i_s = {wallace_tree_cells_109_io_i_s_hi,wallace_tree_cells_109_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_110_io_i_inter_c = wallace_tree_cells_109_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_110_io_i_s = {wallace_tree_cells_110_io_i_s_hi,wallace_tree_cells_110_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_111_io_i_inter_c = wallace_tree_cells_110_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_111_io_i_s = {wallace_tree_cells_111_io_i_s_hi,wallace_tree_cells_111_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_112_io_i_inter_c = wallace_tree_cells_111_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_112_io_i_s = {wallace_tree_cells_112_io_i_s_hi,wallace_tree_cells_112_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_113_io_i_inter_c = wallace_tree_cells_112_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_113_io_i_s = {wallace_tree_cells_113_io_i_s_hi,wallace_tree_cells_113_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_114_io_i_inter_c = wallace_tree_cells_113_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_114_io_i_s = {wallace_tree_cells_114_io_i_s_hi,wallace_tree_cells_114_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_115_io_i_inter_c = wallace_tree_cells_114_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_115_io_i_s = {wallace_tree_cells_115_io_i_s_hi,wallace_tree_cells_115_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_116_io_i_inter_c = wallace_tree_cells_115_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_116_io_i_s = {wallace_tree_cells_116_io_i_s_hi,wallace_tree_cells_116_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_117_io_i_inter_c = wallace_tree_cells_116_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_117_io_i_s = {wallace_tree_cells_117_io_i_s_hi,wallace_tree_cells_117_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_118_io_i_inter_c = wallace_tree_cells_117_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_118_io_i_s = {wallace_tree_cells_118_io_i_s_hi,wallace_tree_cells_118_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_119_io_i_inter_c = wallace_tree_cells_118_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_119_io_i_s = {wallace_tree_cells_119_io_i_s_hi,wallace_tree_cells_119_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_120_io_i_inter_c = wallace_tree_cells_119_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_120_io_i_s = {wallace_tree_cells_120_io_i_s_hi,wallace_tree_cells_120_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_121_io_i_inter_c = wallace_tree_cells_120_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_121_io_i_s = {wallace_tree_cells_121_io_i_s_hi,wallace_tree_cells_121_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_122_io_i_inter_c = wallace_tree_cells_121_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_122_io_i_s = {wallace_tree_cells_122_io_i_s_hi,wallace_tree_cells_122_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_123_io_i_inter_c = wallace_tree_cells_122_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_123_io_i_s = {wallace_tree_cells_123_io_i_s_hi,wallace_tree_cells_123_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_124_io_i_inter_c = wallace_tree_cells_123_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_124_io_i_s = {wallace_tree_cells_124_io_i_s_hi,wallace_tree_cells_124_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_125_io_i_inter_c = wallace_tree_cells_124_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_125_io_i_s = {wallace_tree_cells_125_io_i_s_hi,wallace_tree_cells_125_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_126_io_i_inter_c = wallace_tree_cells_125_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_126_io_i_s = {wallace_tree_cells_126_io_i_s_hi,wallace_tree_cells_126_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_127_io_i_inter_c = wallace_tree_cells_126_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_127_io_i_s = {wallace_tree_cells_127_io_i_s_hi,wallace_tree_cells_127_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_128_io_i_inter_c = wallace_tree_cells_127_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_128_io_i_s = {wallace_tree_cells_128_io_i_s_hi,wallace_tree_cells_128_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_129_io_i_inter_c = wallace_tree_cells_128_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_129_io_i_s = {wallace_tree_cells_129_io_i_s_hi,wallace_tree_cells_129_io_i_s_lo}; // @[wallace_tree.scala 147:56]
  assign wallace_tree_cells_130_io_i_inter_c = wallace_tree_cells_129_io_o_inter_c; // @[wallace_tree.scala 152:44]
  assign wallace_tree_cells_130_io_i_s = {wallace_tree_cells_130_io_i_s_hi,wallace_tree_cells_130_io_i_s_lo}; // @[wallace_tree.scala 147:56]
endmodule

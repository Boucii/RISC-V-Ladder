module BPU(
  input         clock,
  input         reset,
  input  [63:0] io_i_addr,
  input         io_i_branch_resolve_pack_valid,
  input         io_i_branch_resolve_pack_taken,
  input  [63:0] io_i_branch_resolve_pack_pc,
  input  [63:0] io_i_branch_resolve_pack_target,
  input         io_i_branch_resolve_pack_prediction_valid,
  input         io_i_branch_presolve_pack_valid,
  input  [63:0] io_i_branch_presolve_pack_pc,
  output        io_o_branch_predict_pack_valid,
  output [63:0] io_o_branch_predict_pack_target,
  output        io_o_branch_predict_pack_taken
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [63:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [63:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [63:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [63:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [63:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [63:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [63:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [63:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [63:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [63:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [63:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [63:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [63:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [63:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [63:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [63:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [63:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [63:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [63:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [63:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [63:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [63:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [63:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [63:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [63:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [63:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [63:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [63:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [63:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [63:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [63:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [63:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [63:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [63:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [63:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [63:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [63:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [63:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [63:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [63:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [63:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [63:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [63:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [63:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [63:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [63:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [63:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [63:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [63:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [63:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [63:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [63:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [63:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [63:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [63:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [63:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [63:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [63:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [63:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [63:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [63:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [63:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [63:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [63:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [63:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [63:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [63:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [63:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [63:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [63:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [63:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [63:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [63:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [63:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [63:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [63:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [63:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [63:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [63:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [63:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [63:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [63:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [63:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [63:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [63:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [63:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [63:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [63:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [63:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [63:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [63:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [63:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [63:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [63:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [63:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [63:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [63:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [63:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [63:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [63:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [63:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [63:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [63:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [63:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [63:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [63:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [63:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [63:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [63:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [63:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [63:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [63:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [63:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [63:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [63:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [63:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [63:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [63:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [63:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [63:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [63:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [63:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [63:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [63:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [63:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [63:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [63:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [63:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [63:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [63:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [63:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [63:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [63:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [63:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [63:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [63:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [63:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [63:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [63:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [63:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [63:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [63:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [63:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [63:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [63:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [63:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [63:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [63:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [63:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [63:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [63:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [63:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [63:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [63:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [63:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [63:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [63:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [63:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [63:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [63:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [63:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [63:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [63:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [63:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [63:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [63:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [63:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [63:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [63:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [63:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [63:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [63:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [63:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [63:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [63:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [63:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [63:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [63:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [63:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [63:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [63:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [63:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [63:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [63:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [63:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [63:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [63:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [63:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [63:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [63:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [63:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [63:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [63:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [63:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [63:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [63:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [63:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [63:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [63:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [63:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [63:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [63:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [63:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [63:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [63:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [63:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [63:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [63:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [63:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [63:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [63:0] _RAND_1038;
  reg [31:0] _RAND_1039;
  reg [31:0] _RAND_1040;
  reg [31:0] _RAND_1041;
  reg [63:0] _RAND_1042;
  reg [31:0] _RAND_1043;
  reg [31:0] _RAND_1044;
  reg [31:0] _RAND_1045;
  reg [63:0] _RAND_1046;
  reg [31:0] _RAND_1047;
  reg [31:0] _RAND_1048;
  reg [31:0] _RAND_1049;
  reg [63:0] _RAND_1050;
  reg [31:0] _RAND_1051;
  reg [31:0] _RAND_1052;
  reg [31:0] _RAND_1053;
  reg [63:0] _RAND_1054;
  reg [31:0] _RAND_1055;
  reg [31:0] _RAND_1056;
  reg [31:0] _RAND_1057;
  reg [63:0] _RAND_1058;
  reg [31:0] _RAND_1059;
  reg [31:0] _RAND_1060;
  reg [31:0] _RAND_1061;
  reg [63:0] _RAND_1062;
  reg [31:0] _RAND_1063;
  reg [31:0] _RAND_1064;
  reg [31:0] _RAND_1065;
  reg [63:0] _RAND_1066;
  reg [31:0] _RAND_1067;
  reg [31:0] _RAND_1068;
  reg [31:0] _RAND_1069;
  reg [63:0] _RAND_1070;
  reg [31:0] _RAND_1071;
  reg [31:0] _RAND_1072;
  reg [31:0] _RAND_1073;
  reg [63:0] _RAND_1074;
  reg [31:0] _RAND_1075;
  reg [31:0] _RAND_1076;
  reg [31:0] _RAND_1077;
  reg [63:0] _RAND_1078;
  reg [31:0] _RAND_1079;
  reg [31:0] _RAND_1080;
  reg [31:0] _RAND_1081;
  reg [63:0] _RAND_1082;
  reg [31:0] _RAND_1083;
  reg [31:0] _RAND_1084;
  reg [31:0] _RAND_1085;
  reg [63:0] _RAND_1086;
  reg [31:0] _RAND_1087;
  reg [31:0] _RAND_1088;
  reg [31:0] _RAND_1089;
  reg [63:0] _RAND_1090;
  reg [31:0] _RAND_1091;
  reg [31:0] _RAND_1092;
  reg [31:0] _RAND_1093;
  reg [63:0] _RAND_1094;
  reg [31:0] _RAND_1095;
  reg [31:0] _RAND_1096;
  reg [31:0] _RAND_1097;
  reg [63:0] _RAND_1098;
  reg [31:0] _RAND_1099;
  reg [31:0] _RAND_1100;
  reg [31:0] _RAND_1101;
  reg [63:0] _RAND_1102;
  reg [31:0] _RAND_1103;
  reg [31:0] _RAND_1104;
  reg [31:0] _RAND_1105;
  reg [63:0] _RAND_1106;
  reg [31:0] _RAND_1107;
  reg [31:0] _RAND_1108;
  reg [31:0] _RAND_1109;
  reg [63:0] _RAND_1110;
  reg [31:0] _RAND_1111;
  reg [31:0] _RAND_1112;
  reg [31:0] _RAND_1113;
  reg [63:0] _RAND_1114;
  reg [31:0] _RAND_1115;
  reg [31:0] _RAND_1116;
  reg [31:0] _RAND_1117;
  reg [63:0] _RAND_1118;
  reg [31:0] _RAND_1119;
  reg [31:0] _RAND_1120;
  reg [31:0] _RAND_1121;
  reg [63:0] _RAND_1122;
  reg [31:0] _RAND_1123;
  reg [31:0] _RAND_1124;
  reg [31:0] _RAND_1125;
  reg [63:0] _RAND_1126;
  reg [31:0] _RAND_1127;
  reg [31:0] _RAND_1128;
  reg [31:0] _RAND_1129;
  reg [63:0] _RAND_1130;
  reg [31:0] _RAND_1131;
  reg [31:0] _RAND_1132;
  reg [31:0] _RAND_1133;
  reg [63:0] _RAND_1134;
  reg [31:0] _RAND_1135;
  reg [31:0] _RAND_1136;
  reg [31:0] _RAND_1137;
  reg [63:0] _RAND_1138;
  reg [31:0] _RAND_1139;
  reg [31:0] _RAND_1140;
  reg [31:0] _RAND_1141;
  reg [63:0] _RAND_1142;
  reg [31:0] _RAND_1143;
  reg [31:0] _RAND_1144;
  reg [31:0] _RAND_1145;
  reg [63:0] _RAND_1146;
  reg [31:0] _RAND_1147;
  reg [31:0] _RAND_1148;
  reg [31:0] _RAND_1149;
  reg [63:0] _RAND_1150;
  reg [31:0] _RAND_1151;
  reg [31:0] _RAND_1152;
  reg [31:0] _RAND_1153;
  reg [63:0] _RAND_1154;
  reg [31:0] _RAND_1155;
  reg [31:0] _RAND_1156;
  reg [31:0] _RAND_1157;
  reg [63:0] _RAND_1158;
  reg [31:0] _RAND_1159;
  reg [31:0] _RAND_1160;
  reg [31:0] _RAND_1161;
  reg [63:0] _RAND_1162;
  reg [31:0] _RAND_1163;
  reg [31:0] _RAND_1164;
  reg [31:0] _RAND_1165;
  reg [63:0] _RAND_1166;
  reg [31:0] _RAND_1167;
  reg [31:0] _RAND_1168;
  reg [31:0] _RAND_1169;
  reg [63:0] _RAND_1170;
  reg [31:0] _RAND_1171;
  reg [31:0] _RAND_1172;
  reg [31:0] _RAND_1173;
  reg [63:0] _RAND_1174;
  reg [31:0] _RAND_1175;
  reg [31:0] _RAND_1176;
  reg [31:0] _RAND_1177;
  reg [63:0] _RAND_1178;
  reg [31:0] _RAND_1179;
  reg [31:0] _RAND_1180;
  reg [31:0] _RAND_1181;
  reg [63:0] _RAND_1182;
  reg [31:0] _RAND_1183;
  reg [31:0] _RAND_1184;
  reg [31:0] _RAND_1185;
  reg [63:0] _RAND_1186;
  reg [31:0] _RAND_1187;
  reg [31:0] _RAND_1188;
  reg [31:0] _RAND_1189;
  reg [63:0] _RAND_1190;
  reg [31:0] _RAND_1191;
  reg [31:0] _RAND_1192;
  reg [31:0] _RAND_1193;
  reg [63:0] _RAND_1194;
  reg [31:0] _RAND_1195;
  reg [31:0] _RAND_1196;
  reg [31:0] _RAND_1197;
  reg [63:0] _RAND_1198;
  reg [31:0] _RAND_1199;
  reg [31:0] _RAND_1200;
  reg [31:0] _RAND_1201;
  reg [63:0] _RAND_1202;
  reg [31:0] _RAND_1203;
  reg [31:0] _RAND_1204;
  reg [31:0] _RAND_1205;
  reg [63:0] _RAND_1206;
  reg [31:0] _RAND_1207;
  reg [31:0] _RAND_1208;
  reg [31:0] _RAND_1209;
  reg [63:0] _RAND_1210;
  reg [31:0] _RAND_1211;
  reg [31:0] _RAND_1212;
  reg [31:0] _RAND_1213;
  reg [63:0] _RAND_1214;
  reg [31:0] _RAND_1215;
  reg [31:0] _RAND_1216;
  reg [31:0] _RAND_1217;
  reg [63:0] _RAND_1218;
  reg [31:0] _RAND_1219;
  reg [31:0] _RAND_1220;
  reg [31:0] _RAND_1221;
  reg [63:0] _RAND_1222;
  reg [31:0] _RAND_1223;
  reg [31:0] _RAND_1224;
  reg [31:0] _RAND_1225;
  reg [63:0] _RAND_1226;
  reg [31:0] _RAND_1227;
  reg [31:0] _RAND_1228;
  reg [31:0] _RAND_1229;
  reg [63:0] _RAND_1230;
  reg [31:0] _RAND_1231;
  reg [31:0] _RAND_1232;
  reg [31:0] _RAND_1233;
  reg [63:0] _RAND_1234;
  reg [31:0] _RAND_1235;
  reg [31:0] _RAND_1236;
  reg [31:0] _RAND_1237;
  reg [63:0] _RAND_1238;
  reg [31:0] _RAND_1239;
  reg [31:0] _RAND_1240;
  reg [31:0] _RAND_1241;
  reg [63:0] _RAND_1242;
  reg [31:0] _RAND_1243;
  reg [31:0] _RAND_1244;
  reg [31:0] _RAND_1245;
  reg [63:0] _RAND_1246;
  reg [31:0] _RAND_1247;
  reg [31:0] _RAND_1248;
  reg [31:0] _RAND_1249;
  reg [63:0] _RAND_1250;
  reg [31:0] _RAND_1251;
  reg [31:0] _RAND_1252;
  reg [31:0] _RAND_1253;
  reg [63:0] _RAND_1254;
  reg [31:0] _RAND_1255;
  reg [31:0] _RAND_1256;
  reg [31:0] _RAND_1257;
  reg [63:0] _RAND_1258;
  reg [31:0] _RAND_1259;
  reg [31:0] _RAND_1260;
  reg [31:0] _RAND_1261;
  reg [63:0] _RAND_1262;
  reg [31:0] _RAND_1263;
  reg [31:0] _RAND_1264;
  reg [31:0] _RAND_1265;
  reg [63:0] _RAND_1266;
  reg [31:0] _RAND_1267;
  reg [31:0] _RAND_1268;
  reg [31:0] _RAND_1269;
  reg [63:0] _RAND_1270;
  reg [31:0] _RAND_1271;
  reg [31:0] _RAND_1272;
  reg [31:0] _RAND_1273;
  reg [63:0] _RAND_1274;
  reg [31:0] _RAND_1275;
  reg [31:0] _RAND_1276;
  reg [31:0] _RAND_1277;
  reg [63:0] _RAND_1278;
  reg [31:0] _RAND_1279;
  reg [31:0] _RAND_1280;
  reg [31:0] _RAND_1281;
  reg [63:0] _RAND_1282;
  reg [31:0] _RAND_1283;
  reg [31:0] _RAND_1284;
  reg [31:0] _RAND_1285;
  reg [63:0] _RAND_1286;
  reg [31:0] _RAND_1287;
  reg [31:0] _RAND_1288;
  reg [31:0] _RAND_1289;
  reg [63:0] _RAND_1290;
  reg [31:0] _RAND_1291;
  reg [31:0] _RAND_1292;
  reg [31:0] _RAND_1293;
  reg [63:0] _RAND_1294;
  reg [31:0] _RAND_1295;
  reg [31:0] _RAND_1296;
  reg [31:0] _RAND_1297;
  reg [63:0] _RAND_1298;
  reg [31:0] _RAND_1299;
  reg [31:0] _RAND_1300;
  reg [31:0] _RAND_1301;
  reg [63:0] _RAND_1302;
  reg [31:0] _RAND_1303;
  reg [31:0] _RAND_1304;
  reg [31:0] _RAND_1305;
  reg [63:0] _RAND_1306;
  reg [31:0] _RAND_1307;
  reg [31:0] _RAND_1308;
  reg [31:0] _RAND_1309;
  reg [63:0] _RAND_1310;
  reg [31:0] _RAND_1311;
  reg [31:0] _RAND_1312;
  reg [31:0] _RAND_1313;
  reg [63:0] _RAND_1314;
  reg [31:0] _RAND_1315;
  reg [31:0] _RAND_1316;
  reg [31:0] _RAND_1317;
  reg [63:0] _RAND_1318;
  reg [31:0] _RAND_1319;
  reg [31:0] _RAND_1320;
  reg [31:0] _RAND_1321;
  reg [63:0] _RAND_1322;
  reg [31:0] _RAND_1323;
  reg [31:0] _RAND_1324;
  reg [31:0] _RAND_1325;
  reg [63:0] _RAND_1326;
  reg [31:0] _RAND_1327;
  reg [31:0] _RAND_1328;
  reg [31:0] _RAND_1329;
  reg [63:0] _RAND_1330;
  reg [31:0] _RAND_1331;
  reg [31:0] _RAND_1332;
  reg [31:0] _RAND_1333;
  reg [63:0] _RAND_1334;
  reg [31:0] _RAND_1335;
  reg [31:0] _RAND_1336;
  reg [31:0] _RAND_1337;
  reg [63:0] _RAND_1338;
  reg [31:0] _RAND_1339;
  reg [31:0] _RAND_1340;
  reg [31:0] _RAND_1341;
  reg [63:0] _RAND_1342;
  reg [31:0] _RAND_1343;
  reg [31:0] _RAND_1344;
  reg [31:0] _RAND_1345;
  reg [63:0] _RAND_1346;
  reg [31:0] _RAND_1347;
  reg [31:0] _RAND_1348;
  reg [31:0] _RAND_1349;
  reg [63:0] _RAND_1350;
  reg [31:0] _RAND_1351;
  reg [31:0] _RAND_1352;
  reg [31:0] _RAND_1353;
  reg [63:0] _RAND_1354;
  reg [31:0] _RAND_1355;
  reg [31:0] _RAND_1356;
  reg [31:0] _RAND_1357;
  reg [63:0] _RAND_1358;
  reg [31:0] _RAND_1359;
  reg [31:0] _RAND_1360;
  reg [31:0] _RAND_1361;
  reg [63:0] _RAND_1362;
  reg [31:0] _RAND_1363;
  reg [31:0] _RAND_1364;
  reg [31:0] _RAND_1365;
  reg [63:0] _RAND_1366;
  reg [31:0] _RAND_1367;
  reg [31:0] _RAND_1368;
  reg [31:0] _RAND_1369;
  reg [63:0] _RAND_1370;
  reg [31:0] _RAND_1371;
  reg [31:0] _RAND_1372;
  reg [31:0] _RAND_1373;
  reg [63:0] _RAND_1374;
  reg [31:0] _RAND_1375;
  reg [31:0] _RAND_1376;
  reg [31:0] _RAND_1377;
  reg [63:0] _RAND_1378;
  reg [31:0] _RAND_1379;
  reg [31:0] _RAND_1380;
  reg [31:0] _RAND_1381;
  reg [63:0] _RAND_1382;
  reg [31:0] _RAND_1383;
  reg [31:0] _RAND_1384;
  reg [31:0] _RAND_1385;
  reg [63:0] _RAND_1386;
  reg [31:0] _RAND_1387;
  reg [31:0] _RAND_1388;
  reg [31:0] _RAND_1389;
  reg [63:0] _RAND_1390;
  reg [31:0] _RAND_1391;
  reg [31:0] _RAND_1392;
  reg [31:0] _RAND_1393;
  reg [63:0] _RAND_1394;
  reg [31:0] _RAND_1395;
  reg [31:0] _RAND_1396;
  reg [31:0] _RAND_1397;
  reg [63:0] _RAND_1398;
  reg [31:0] _RAND_1399;
  reg [31:0] _RAND_1400;
  reg [31:0] _RAND_1401;
  reg [63:0] _RAND_1402;
  reg [31:0] _RAND_1403;
  reg [31:0] _RAND_1404;
  reg [31:0] _RAND_1405;
  reg [63:0] _RAND_1406;
  reg [31:0] _RAND_1407;
  reg [31:0] _RAND_1408;
  reg [31:0] _RAND_1409;
  reg [63:0] _RAND_1410;
  reg [31:0] _RAND_1411;
  reg [31:0] _RAND_1412;
  reg [31:0] _RAND_1413;
  reg [63:0] _RAND_1414;
  reg [31:0] _RAND_1415;
  reg [31:0] _RAND_1416;
  reg [31:0] _RAND_1417;
  reg [63:0] _RAND_1418;
  reg [31:0] _RAND_1419;
  reg [31:0] _RAND_1420;
  reg [31:0] _RAND_1421;
  reg [63:0] _RAND_1422;
  reg [31:0] _RAND_1423;
  reg [31:0] _RAND_1424;
  reg [31:0] _RAND_1425;
  reg [63:0] _RAND_1426;
  reg [31:0] _RAND_1427;
  reg [31:0] _RAND_1428;
  reg [31:0] _RAND_1429;
  reg [63:0] _RAND_1430;
  reg [31:0] _RAND_1431;
  reg [31:0] _RAND_1432;
  reg [31:0] _RAND_1433;
  reg [63:0] _RAND_1434;
  reg [31:0] _RAND_1435;
  reg [31:0] _RAND_1436;
  reg [31:0] _RAND_1437;
  reg [63:0] _RAND_1438;
  reg [31:0] _RAND_1439;
  reg [31:0] _RAND_1440;
  reg [31:0] _RAND_1441;
  reg [63:0] _RAND_1442;
  reg [31:0] _RAND_1443;
  reg [31:0] _RAND_1444;
  reg [31:0] _RAND_1445;
  reg [63:0] _RAND_1446;
  reg [31:0] _RAND_1447;
  reg [31:0] _RAND_1448;
  reg [31:0] _RAND_1449;
  reg [63:0] _RAND_1450;
  reg [31:0] _RAND_1451;
  reg [31:0] _RAND_1452;
  reg [31:0] _RAND_1453;
  reg [63:0] _RAND_1454;
  reg [31:0] _RAND_1455;
  reg [31:0] _RAND_1456;
  reg [31:0] _RAND_1457;
  reg [63:0] _RAND_1458;
  reg [31:0] _RAND_1459;
  reg [31:0] _RAND_1460;
  reg [31:0] _RAND_1461;
  reg [63:0] _RAND_1462;
  reg [31:0] _RAND_1463;
  reg [31:0] _RAND_1464;
  reg [31:0] _RAND_1465;
  reg [63:0] _RAND_1466;
  reg [31:0] _RAND_1467;
  reg [31:0] _RAND_1468;
  reg [31:0] _RAND_1469;
  reg [63:0] _RAND_1470;
  reg [31:0] _RAND_1471;
  reg [31:0] _RAND_1472;
  reg [31:0] _RAND_1473;
  reg [63:0] _RAND_1474;
  reg [31:0] _RAND_1475;
  reg [31:0] _RAND_1476;
  reg [31:0] _RAND_1477;
  reg [63:0] _RAND_1478;
  reg [31:0] _RAND_1479;
  reg [31:0] _RAND_1480;
  reg [31:0] _RAND_1481;
  reg [63:0] _RAND_1482;
  reg [31:0] _RAND_1483;
  reg [31:0] _RAND_1484;
  reg [31:0] _RAND_1485;
  reg [63:0] _RAND_1486;
  reg [31:0] _RAND_1487;
  reg [31:0] _RAND_1488;
  reg [31:0] _RAND_1489;
  reg [63:0] _RAND_1490;
  reg [31:0] _RAND_1491;
  reg [31:0] _RAND_1492;
  reg [31:0] _RAND_1493;
  reg [63:0] _RAND_1494;
  reg [31:0] _RAND_1495;
  reg [31:0] _RAND_1496;
  reg [31:0] _RAND_1497;
  reg [63:0] _RAND_1498;
  reg [31:0] _RAND_1499;
  reg [31:0] _RAND_1500;
  reg [31:0] _RAND_1501;
  reg [63:0] _RAND_1502;
  reg [31:0] _RAND_1503;
  reg [31:0] _RAND_1504;
  reg [31:0] _RAND_1505;
  reg [63:0] _RAND_1506;
  reg [31:0] _RAND_1507;
  reg [31:0] _RAND_1508;
  reg [31:0] _RAND_1509;
  reg [63:0] _RAND_1510;
  reg [31:0] _RAND_1511;
  reg [31:0] _RAND_1512;
  reg [31:0] _RAND_1513;
  reg [63:0] _RAND_1514;
  reg [31:0] _RAND_1515;
  reg [31:0] _RAND_1516;
  reg [31:0] _RAND_1517;
  reg [63:0] _RAND_1518;
  reg [31:0] _RAND_1519;
  reg [31:0] _RAND_1520;
  reg [31:0] _RAND_1521;
  reg [63:0] _RAND_1522;
  reg [31:0] _RAND_1523;
  reg [31:0] _RAND_1524;
  reg [31:0] _RAND_1525;
  reg [63:0] _RAND_1526;
  reg [31:0] _RAND_1527;
  reg [31:0] _RAND_1528;
  reg [31:0] _RAND_1529;
  reg [63:0] _RAND_1530;
  reg [31:0] _RAND_1531;
  reg [31:0] _RAND_1532;
  reg [31:0] _RAND_1533;
  reg [63:0] _RAND_1534;
  reg [31:0] _RAND_1535;
  reg [31:0] _RAND_1536;
  reg [31:0] _RAND_1537;
  reg [63:0] _RAND_1538;
  reg [31:0] _RAND_1539;
  reg [31:0] _RAND_1540;
  reg [31:0] _RAND_1541;
  reg [63:0] _RAND_1542;
  reg [31:0] _RAND_1543;
  reg [31:0] _RAND_1544;
  reg [31:0] _RAND_1545;
  reg [63:0] _RAND_1546;
  reg [31:0] _RAND_1547;
  reg [31:0] _RAND_1548;
  reg [31:0] _RAND_1549;
  reg [63:0] _RAND_1550;
  reg [31:0] _RAND_1551;
  reg [31:0] _RAND_1552;
  reg [31:0] _RAND_1553;
  reg [63:0] _RAND_1554;
  reg [31:0] _RAND_1555;
  reg [31:0] _RAND_1556;
  reg [31:0] _RAND_1557;
  reg [63:0] _RAND_1558;
  reg [31:0] _RAND_1559;
  reg [31:0] _RAND_1560;
  reg [31:0] _RAND_1561;
  reg [63:0] _RAND_1562;
  reg [31:0] _RAND_1563;
  reg [31:0] _RAND_1564;
  reg [31:0] _RAND_1565;
  reg [63:0] _RAND_1566;
  reg [31:0] _RAND_1567;
  reg [31:0] _RAND_1568;
  reg [31:0] _RAND_1569;
  reg [63:0] _RAND_1570;
  reg [31:0] _RAND_1571;
  reg [31:0] _RAND_1572;
  reg [31:0] _RAND_1573;
  reg [63:0] _RAND_1574;
  reg [31:0] _RAND_1575;
  reg [31:0] _RAND_1576;
  reg [31:0] _RAND_1577;
  reg [63:0] _RAND_1578;
  reg [31:0] _RAND_1579;
  reg [31:0] _RAND_1580;
  reg [31:0] _RAND_1581;
  reg [63:0] _RAND_1582;
  reg [31:0] _RAND_1583;
  reg [31:0] _RAND_1584;
  reg [31:0] _RAND_1585;
  reg [63:0] _RAND_1586;
  reg [31:0] _RAND_1587;
  reg [31:0] _RAND_1588;
  reg [31:0] _RAND_1589;
  reg [63:0] _RAND_1590;
  reg [31:0] _RAND_1591;
  reg [31:0] _RAND_1592;
  reg [31:0] _RAND_1593;
  reg [63:0] _RAND_1594;
  reg [31:0] _RAND_1595;
  reg [31:0] _RAND_1596;
  reg [31:0] _RAND_1597;
  reg [63:0] _RAND_1598;
  reg [31:0] _RAND_1599;
  reg [31:0] _RAND_1600;
  reg [31:0] _RAND_1601;
  reg [63:0] _RAND_1602;
  reg [31:0] _RAND_1603;
  reg [31:0] _RAND_1604;
  reg [31:0] _RAND_1605;
  reg [63:0] _RAND_1606;
  reg [31:0] _RAND_1607;
  reg [31:0] _RAND_1608;
  reg [31:0] _RAND_1609;
  reg [63:0] _RAND_1610;
  reg [31:0] _RAND_1611;
  reg [31:0] _RAND_1612;
  reg [31:0] _RAND_1613;
  reg [63:0] _RAND_1614;
  reg [31:0] _RAND_1615;
  reg [31:0] _RAND_1616;
  reg [31:0] _RAND_1617;
  reg [63:0] _RAND_1618;
  reg [31:0] _RAND_1619;
  reg [31:0] _RAND_1620;
  reg [31:0] _RAND_1621;
  reg [63:0] _RAND_1622;
  reg [31:0] _RAND_1623;
  reg [31:0] _RAND_1624;
  reg [31:0] _RAND_1625;
  reg [63:0] _RAND_1626;
  reg [31:0] _RAND_1627;
  reg [31:0] _RAND_1628;
  reg [31:0] _RAND_1629;
  reg [63:0] _RAND_1630;
  reg [31:0] _RAND_1631;
  reg [31:0] _RAND_1632;
  reg [31:0] _RAND_1633;
  reg [63:0] _RAND_1634;
  reg [31:0] _RAND_1635;
  reg [31:0] _RAND_1636;
  reg [31:0] _RAND_1637;
  reg [63:0] _RAND_1638;
  reg [31:0] _RAND_1639;
  reg [31:0] _RAND_1640;
  reg [31:0] _RAND_1641;
  reg [63:0] _RAND_1642;
  reg [31:0] _RAND_1643;
  reg [31:0] _RAND_1644;
  reg [31:0] _RAND_1645;
  reg [63:0] _RAND_1646;
  reg [31:0] _RAND_1647;
  reg [31:0] _RAND_1648;
  reg [31:0] _RAND_1649;
  reg [63:0] _RAND_1650;
  reg [31:0] _RAND_1651;
  reg [31:0] _RAND_1652;
  reg [31:0] _RAND_1653;
  reg [63:0] _RAND_1654;
  reg [31:0] _RAND_1655;
  reg [31:0] _RAND_1656;
  reg [31:0] _RAND_1657;
  reg [63:0] _RAND_1658;
  reg [31:0] _RAND_1659;
  reg [31:0] _RAND_1660;
  reg [31:0] _RAND_1661;
  reg [63:0] _RAND_1662;
  reg [31:0] _RAND_1663;
  reg [31:0] _RAND_1664;
  reg [31:0] _RAND_1665;
  reg [63:0] _RAND_1666;
  reg [31:0] _RAND_1667;
  reg [31:0] _RAND_1668;
  reg [31:0] _RAND_1669;
  reg [63:0] _RAND_1670;
  reg [31:0] _RAND_1671;
  reg [31:0] _RAND_1672;
  reg [31:0] _RAND_1673;
  reg [63:0] _RAND_1674;
  reg [31:0] _RAND_1675;
  reg [31:0] _RAND_1676;
  reg [31:0] _RAND_1677;
  reg [63:0] _RAND_1678;
  reg [31:0] _RAND_1679;
  reg [31:0] _RAND_1680;
  reg [31:0] _RAND_1681;
  reg [63:0] _RAND_1682;
  reg [31:0] _RAND_1683;
  reg [31:0] _RAND_1684;
  reg [31:0] _RAND_1685;
  reg [63:0] _RAND_1686;
  reg [31:0] _RAND_1687;
  reg [31:0] _RAND_1688;
  reg [31:0] _RAND_1689;
  reg [63:0] _RAND_1690;
  reg [31:0] _RAND_1691;
  reg [31:0] _RAND_1692;
  reg [31:0] _RAND_1693;
  reg [63:0] _RAND_1694;
  reg [31:0] _RAND_1695;
  reg [31:0] _RAND_1696;
  reg [31:0] _RAND_1697;
  reg [63:0] _RAND_1698;
  reg [31:0] _RAND_1699;
  reg [31:0] _RAND_1700;
  reg [31:0] _RAND_1701;
  reg [63:0] _RAND_1702;
  reg [31:0] _RAND_1703;
  reg [31:0] _RAND_1704;
  reg [31:0] _RAND_1705;
  reg [63:0] _RAND_1706;
  reg [31:0] _RAND_1707;
  reg [31:0] _RAND_1708;
  reg [31:0] _RAND_1709;
  reg [63:0] _RAND_1710;
  reg [31:0] _RAND_1711;
  reg [31:0] _RAND_1712;
  reg [31:0] _RAND_1713;
  reg [63:0] _RAND_1714;
  reg [31:0] _RAND_1715;
  reg [31:0] _RAND_1716;
  reg [31:0] _RAND_1717;
  reg [63:0] _RAND_1718;
  reg [31:0] _RAND_1719;
  reg [31:0] _RAND_1720;
  reg [31:0] _RAND_1721;
  reg [63:0] _RAND_1722;
  reg [31:0] _RAND_1723;
  reg [31:0] _RAND_1724;
  reg [31:0] _RAND_1725;
  reg [63:0] _RAND_1726;
  reg [31:0] _RAND_1727;
  reg [31:0] _RAND_1728;
  reg [31:0] _RAND_1729;
  reg [63:0] _RAND_1730;
  reg [31:0] _RAND_1731;
  reg [31:0] _RAND_1732;
  reg [31:0] _RAND_1733;
  reg [63:0] _RAND_1734;
  reg [31:0] _RAND_1735;
  reg [31:0] _RAND_1736;
  reg [31:0] _RAND_1737;
  reg [63:0] _RAND_1738;
  reg [31:0] _RAND_1739;
  reg [31:0] _RAND_1740;
  reg [31:0] _RAND_1741;
  reg [63:0] _RAND_1742;
  reg [31:0] _RAND_1743;
  reg [31:0] _RAND_1744;
  reg [31:0] _RAND_1745;
  reg [63:0] _RAND_1746;
  reg [31:0] _RAND_1747;
  reg [31:0] _RAND_1748;
  reg [31:0] _RAND_1749;
  reg [63:0] _RAND_1750;
  reg [31:0] _RAND_1751;
  reg [31:0] _RAND_1752;
  reg [31:0] _RAND_1753;
  reg [63:0] _RAND_1754;
  reg [31:0] _RAND_1755;
  reg [31:0] _RAND_1756;
  reg [31:0] _RAND_1757;
  reg [63:0] _RAND_1758;
  reg [31:0] _RAND_1759;
  reg [31:0] _RAND_1760;
  reg [31:0] _RAND_1761;
  reg [63:0] _RAND_1762;
  reg [31:0] _RAND_1763;
  reg [31:0] _RAND_1764;
  reg [31:0] _RAND_1765;
  reg [63:0] _RAND_1766;
  reg [31:0] _RAND_1767;
  reg [31:0] _RAND_1768;
  reg [31:0] _RAND_1769;
  reg [63:0] _RAND_1770;
  reg [31:0] _RAND_1771;
  reg [31:0] _RAND_1772;
  reg [31:0] _RAND_1773;
  reg [63:0] _RAND_1774;
  reg [31:0] _RAND_1775;
  reg [31:0] _RAND_1776;
  reg [31:0] _RAND_1777;
  reg [63:0] _RAND_1778;
  reg [31:0] _RAND_1779;
  reg [31:0] _RAND_1780;
  reg [31:0] _RAND_1781;
  reg [63:0] _RAND_1782;
  reg [31:0] _RAND_1783;
  reg [31:0] _RAND_1784;
  reg [31:0] _RAND_1785;
  reg [63:0] _RAND_1786;
  reg [31:0] _RAND_1787;
  reg [31:0] _RAND_1788;
  reg [31:0] _RAND_1789;
  reg [63:0] _RAND_1790;
  reg [31:0] _RAND_1791;
  reg [31:0] _RAND_1792;
  reg [31:0] _RAND_1793;
  reg [63:0] _RAND_1794;
  reg [31:0] _RAND_1795;
  reg [31:0] _RAND_1796;
  reg [31:0] _RAND_1797;
  reg [63:0] _RAND_1798;
  reg [31:0] _RAND_1799;
  reg [31:0] _RAND_1800;
  reg [31:0] _RAND_1801;
  reg [63:0] _RAND_1802;
  reg [31:0] _RAND_1803;
  reg [31:0] _RAND_1804;
  reg [31:0] _RAND_1805;
  reg [63:0] _RAND_1806;
  reg [31:0] _RAND_1807;
  reg [31:0] _RAND_1808;
  reg [31:0] _RAND_1809;
  reg [63:0] _RAND_1810;
  reg [31:0] _RAND_1811;
  reg [31:0] _RAND_1812;
  reg [31:0] _RAND_1813;
  reg [63:0] _RAND_1814;
  reg [31:0] _RAND_1815;
  reg [31:0] _RAND_1816;
  reg [31:0] _RAND_1817;
  reg [63:0] _RAND_1818;
  reg [31:0] _RAND_1819;
  reg [31:0] _RAND_1820;
  reg [31:0] _RAND_1821;
  reg [63:0] _RAND_1822;
  reg [31:0] _RAND_1823;
  reg [31:0] _RAND_1824;
  reg [31:0] _RAND_1825;
  reg [63:0] _RAND_1826;
  reg [31:0] _RAND_1827;
  reg [31:0] _RAND_1828;
  reg [31:0] _RAND_1829;
  reg [63:0] _RAND_1830;
  reg [31:0] _RAND_1831;
  reg [31:0] _RAND_1832;
  reg [31:0] _RAND_1833;
  reg [63:0] _RAND_1834;
  reg [31:0] _RAND_1835;
  reg [31:0] _RAND_1836;
  reg [31:0] _RAND_1837;
  reg [63:0] _RAND_1838;
  reg [31:0] _RAND_1839;
  reg [31:0] _RAND_1840;
  reg [31:0] _RAND_1841;
  reg [63:0] _RAND_1842;
  reg [31:0] _RAND_1843;
  reg [31:0] _RAND_1844;
  reg [31:0] _RAND_1845;
  reg [63:0] _RAND_1846;
  reg [31:0] _RAND_1847;
  reg [31:0] _RAND_1848;
  reg [31:0] _RAND_1849;
  reg [63:0] _RAND_1850;
  reg [31:0] _RAND_1851;
  reg [31:0] _RAND_1852;
  reg [31:0] _RAND_1853;
  reg [63:0] _RAND_1854;
  reg [31:0] _RAND_1855;
  reg [31:0] _RAND_1856;
  reg [31:0] _RAND_1857;
  reg [63:0] _RAND_1858;
  reg [31:0] _RAND_1859;
  reg [31:0] _RAND_1860;
  reg [31:0] _RAND_1861;
  reg [63:0] _RAND_1862;
  reg [31:0] _RAND_1863;
  reg [31:0] _RAND_1864;
  reg [31:0] _RAND_1865;
  reg [63:0] _RAND_1866;
  reg [31:0] _RAND_1867;
  reg [31:0] _RAND_1868;
  reg [31:0] _RAND_1869;
  reg [63:0] _RAND_1870;
  reg [31:0] _RAND_1871;
  reg [31:0] _RAND_1872;
  reg [31:0] _RAND_1873;
  reg [63:0] _RAND_1874;
  reg [31:0] _RAND_1875;
  reg [31:0] _RAND_1876;
  reg [31:0] _RAND_1877;
  reg [63:0] _RAND_1878;
  reg [31:0] _RAND_1879;
  reg [31:0] _RAND_1880;
  reg [31:0] _RAND_1881;
  reg [63:0] _RAND_1882;
  reg [31:0] _RAND_1883;
  reg [31:0] _RAND_1884;
  reg [31:0] _RAND_1885;
  reg [63:0] _RAND_1886;
  reg [31:0] _RAND_1887;
  reg [31:0] _RAND_1888;
  reg [31:0] _RAND_1889;
  reg [63:0] _RAND_1890;
  reg [31:0] _RAND_1891;
  reg [31:0] _RAND_1892;
  reg [31:0] _RAND_1893;
  reg [63:0] _RAND_1894;
  reg [31:0] _RAND_1895;
  reg [31:0] _RAND_1896;
  reg [31:0] _RAND_1897;
  reg [63:0] _RAND_1898;
  reg [31:0] _RAND_1899;
  reg [31:0] _RAND_1900;
  reg [31:0] _RAND_1901;
  reg [63:0] _RAND_1902;
  reg [31:0] _RAND_1903;
  reg [31:0] _RAND_1904;
  reg [31:0] _RAND_1905;
  reg [63:0] _RAND_1906;
  reg [31:0] _RAND_1907;
  reg [31:0] _RAND_1908;
  reg [31:0] _RAND_1909;
  reg [63:0] _RAND_1910;
  reg [31:0] _RAND_1911;
  reg [31:0] _RAND_1912;
  reg [31:0] _RAND_1913;
  reg [63:0] _RAND_1914;
  reg [31:0] _RAND_1915;
  reg [31:0] _RAND_1916;
  reg [31:0] _RAND_1917;
  reg [63:0] _RAND_1918;
  reg [31:0] _RAND_1919;
  reg [31:0] _RAND_1920;
  reg [31:0] _RAND_1921;
  reg [63:0] _RAND_1922;
  reg [31:0] _RAND_1923;
  reg [31:0] _RAND_1924;
  reg [31:0] _RAND_1925;
  reg [63:0] _RAND_1926;
  reg [31:0] _RAND_1927;
  reg [31:0] _RAND_1928;
  reg [31:0] _RAND_1929;
  reg [63:0] _RAND_1930;
  reg [31:0] _RAND_1931;
  reg [31:0] _RAND_1932;
  reg [31:0] _RAND_1933;
  reg [63:0] _RAND_1934;
  reg [31:0] _RAND_1935;
  reg [31:0] _RAND_1936;
  reg [31:0] _RAND_1937;
  reg [63:0] _RAND_1938;
  reg [31:0] _RAND_1939;
  reg [31:0] _RAND_1940;
  reg [31:0] _RAND_1941;
  reg [63:0] _RAND_1942;
  reg [31:0] _RAND_1943;
  reg [31:0] _RAND_1944;
  reg [31:0] _RAND_1945;
  reg [63:0] _RAND_1946;
  reg [31:0] _RAND_1947;
  reg [31:0] _RAND_1948;
  reg [31:0] _RAND_1949;
  reg [63:0] _RAND_1950;
  reg [31:0] _RAND_1951;
  reg [31:0] _RAND_1952;
  reg [31:0] _RAND_1953;
  reg [63:0] _RAND_1954;
  reg [31:0] _RAND_1955;
  reg [31:0] _RAND_1956;
  reg [31:0] _RAND_1957;
  reg [63:0] _RAND_1958;
  reg [31:0] _RAND_1959;
  reg [31:0] _RAND_1960;
  reg [31:0] _RAND_1961;
  reg [63:0] _RAND_1962;
  reg [31:0] _RAND_1963;
  reg [31:0] _RAND_1964;
  reg [31:0] _RAND_1965;
  reg [63:0] _RAND_1966;
  reg [31:0] _RAND_1967;
  reg [31:0] _RAND_1968;
  reg [31:0] _RAND_1969;
  reg [63:0] _RAND_1970;
  reg [31:0] _RAND_1971;
  reg [31:0] _RAND_1972;
  reg [31:0] _RAND_1973;
  reg [63:0] _RAND_1974;
  reg [31:0] _RAND_1975;
  reg [31:0] _RAND_1976;
  reg [31:0] _RAND_1977;
  reg [63:0] _RAND_1978;
  reg [31:0] _RAND_1979;
  reg [31:0] _RAND_1980;
  reg [31:0] _RAND_1981;
  reg [63:0] _RAND_1982;
  reg [31:0] _RAND_1983;
  reg [31:0] _RAND_1984;
  reg [31:0] _RAND_1985;
  reg [63:0] _RAND_1986;
  reg [31:0] _RAND_1987;
  reg [31:0] _RAND_1988;
  reg [31:0] _RAND_1989;
  reg [63:0] _RAND_1990;
  reg [31:0] _RAND_1991;
  reg [31:0] _RAND_1992;
  reg [31:0] _RAND_1993;
  reg [63:0] _RAND_1994;
  reg [31:0] _RAND_1995;
  reg [31:0] _RAND_1996;
  reg [31:0] _RAND_1997;
  reg [63:0] _RAND_1998;
  reg [31:0] _RAND_1999;
  reg [31:0] _RAND_2000;
  reg [31:0] _RAND_2001;
  reg [63:0] _RAND_2002;
  reg [31:0] _RAND_2003;
  reg [31:0] _RAND_2004;
  reg [31:0] _RAND_2005;
  reg [63:0] _RAND_2006;
  reg [31:0] _RAND_2007;
  reg [31:0] _RAND_2008;
  reg [31:0] _RAND_2009;
  reg [63:0] _RAND_2010;
  reg [31:0] _RAND_2011;
  reg [31:0] _RAND_2012;
  reg [31:0] _RAND_2013;
  reg [63:0] _RAND_2014;
  reg [31:0] _RAND_2015;
  reg [31:0] _RAND_2016;
  reg [31:0] _RAND_2017;
  reg [63:0] _RAND_2018;
  reg [31:0] _RAND_2019;
  reg [31:0] _RAND_2020;
  reg [31:0] _RAND_2021;
  reg [63:0] _RAND_2022;
  reg [31:0] _RAND_2023;
  reg [31:0] _RAND_2024;
  reg [31:0] _RAND_2025;
  reg [63:0] _RAND_2026;
  reg [31:0] _RAND_2027;
  reg [31:0] _RAND_2028;
  reg [31:0] _RAND_2029;
  reg [63:0] _RAND_2030;
  reg [31:0] _RAND_2031;
  reg [31:0] _RAND_2032;
  reg [31:0] _RAND_2033;
  reg [63:0] _RAND_2034;
  reg [31:0] _RAND_2035;
  reg [31:0] _RAND_2036;
  reg [31:0] _RAND_2037;
  reg [63:0] _RAND_2038;
  reg [31:0] _RAND_2039;
  reg [31:0] _RAND_2040;
  reg [31:0] _RAND_2041;
  reg [63:0] _RAND_2042;
  reg [31:0] _RAND_2043;
  reg [31:0] _RAND_2044;
  reg [31:0] _RAND_2045;
  reg [63:0] _RAND_2046;
  reg [31:0] _RAND_2047;
  reg [31:0] _RAND_2048;
`endif // RANDOMIZE_REG_INIT
  reg  btb_0_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_0_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_0_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_0_bht; // @[branch_predictor.scala 30:22]
  reg  btb_1_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_1_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_1_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_1_bht; // @[branch_predictor.scala 30:22]
  reg  btb_2_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_2_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_2_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_2_bht; // @[branch_predictor.scala 30:22]
  reg  btb_3_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_3_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_3_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_3_bht; // @[branch_predictor.scala 30:22]
  reg  btb_4_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_4_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_4_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_4_bht; // @[branch_predictor.scala 30:22]
  reg  btb_5_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_5_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_5_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_5_bht; // @[branch_predictor.scala 30:22]
  reg  btb_6_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_6_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_6_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_6_bht; // @[branch_predictor.scala 30:22]
  reg  btb_7_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_7_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_7_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_7_bht; // @[branch_predictor.scala 30:22]
  reg  btb_8_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_8_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_8_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_8_bht; // @[branch_predictor.scala 30:22]
  reg  btb_9_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_9_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_9_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_9_bht; // @[branch_predictor.scala 30:22]
  reg  btb_10_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_10_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_10_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_10_bht; // @[branch_predictor.scala 30:22]
  reg  btb_11_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_11_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_11_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_11_bht; // @[branch_predictor.scala 30:22]
  reg  btb_12_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_12_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_12_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_12_bht; // @[branch_predictor.scala 30:22]
  reg  btb_13_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_13_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_13_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_13_bht; // @[branch_predictor.scala 30:22]
  reg  btb_14_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_14_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_14_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_14_bht; // @[branch_predictor.scala 30:22]
  reg  btb_15_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_15_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_15_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_15_bht; // @[branch_predictor.scala 30:22]
  reg  btb_16_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_16_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_16_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_16_bht; // @[branch_predictor.scala 30:22]
  reg  btb_17_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_17_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_17_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_17_bht; // @[branch_predictor.scala 30:22]
  reg  btb_18_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_18_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_18_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_18_bht; // @[branch_predictor.scala 30:22]
  reg  btb_19_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_19_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_19_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_19_bht; // @[branch_predictor.scala 30:22]
  reg  btb_20_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_20_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_20_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_20_bht; // @[branch_predictor.scala 30:22]
  reg  btb_21_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_21_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_21_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_21_bht; // @[branch_predictor.scala 30:22]
  reg  btb_22_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_22_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_22_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_22_bht; // @[branch_predictor.scala 30:22]
  reg  btb_23_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_23_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_23_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_23_bht; // @[branch_predictor.scala 30:22]
  reg  btb_24_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_24_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_24_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_24_bht; // @[branch_predictor.scala 30:22]
  reg  btb_25_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_25_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_25_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_25_bht; // @[branch_predictor.scala 30:22]
  reg  btb_26_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_26_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_26_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_26_bht; // @[branch_predictor.scala 30:22]
  reg  btb_27_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_27_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_27_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_27_bht; // @[branch_predictor.scala 30:22]
  reg  btb_28_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_28_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_28_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_28_bht; // @[branch_predictor.scala 30:22]
  reg  btb_29_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_29_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_29_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_29_bht; // @[branch_predictor.scala 30:22]
  reg  btb_30_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_30_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_30_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_30_bht; // @[branch_predictor.scala 30:22]
  reg  btb_31_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_31_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_31_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_31_bht; // @[branch_predictor.scala 30:22]
  reg  btb_32_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_32_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_32_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_32_bht; // @[branch_predictor.scala 30:22]
  reg  btb_33_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_33_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_33_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_33_bht; // @[branch_predictor.scala 30:22]
  reg  btb_34_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_34_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_34_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_34_bht; // @[branch_predictor.scala 30:22]
  reg  btb_35_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_35_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_35_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_35_bht; // @[branch_predictor.scala 30:22]
  reg  btb_36_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_36_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_36_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_36_bht; // @[branch_predictor.scala 30:22]
  reg  btb_37_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_37_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_37_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_37_bht; // @[branch_predictor.scala 30:22]
  reg  btb_38_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_38_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_38_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_38_bht; // @[branch_predictor.scala 30:22]
  reg  btb_39_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_39_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_39_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_39_bht; // @[branch_predictor.scala 30:22]
  reg  btb_40_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_40_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_40_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_40_bht; // @[branch_predictor.scala 30:22]
  reg  btb_41_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_41_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_41_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_41_bht; // @[branch_predictor.scala 30:22]
  reg  btb_42_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_42_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_42_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_42_bht; // @[branch_predictor.scala 30:22]
  reg  btb_43_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_43_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_43_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_43_bht; // @[branch_predictor.scala 30:22]
  reg  btb_44_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_44_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_44_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_44_bht; // @[branch_predictor.scala 30:22]
  reg  btb_45_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_45_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_45_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_45_bht; // @[branch_predictor.scala 30:22]
  reg  btb_46_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_46_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_46_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_46_bht; // @[branch_predictor.scala 30:22]
  reg  btb_47_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_47_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_47_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_47_bht; // @[branch_predictor.scala 30:22]
  reg  btb_48_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_48_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_48_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_48_bht; // @[branch_predictor.scala 30:22]
  reg  btb_49_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_49_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_49_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_49_bht; // @[branch_predictor.scala 30:22]
  reg  btb_50_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_50_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_50_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_50_bht; // @[branch_predictor.scala 30:22]
  reg  btb_51_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_51_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_51_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_51_bht; // @[branch_predictor.scala 30:22]
  reg  btb_52_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_52_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_52_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_52_bht; // @[branch_predictor.scala 30:22]
  reg  btb_53_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_53_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_53_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_53_bht; // @[branch_predictor.scala 30:22]
  reg  btb_54_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_54_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_54_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_54_bht; // @[branch_predictor.scala 30:22]
  reg  btb_55_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_55_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_55_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_55_bht; // @[branch_predictor.scala 30:22]
  reg  btb_56_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_56_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_56_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_56_bht; // @[branch_predictor.scala 30:22]
  reg  btb_57_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_57_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_57_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_57_bht; // @[branch_predictor.scala 30:22]
  reg  btb_58_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_58_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_58_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_58_bht; // @[branch_predictor.scala 30:22]
  reg  btb_59_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_59_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_59_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_59_bht; // @[branch_predictor.scala 30:22]
  reg  btb_60_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_60_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_60_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_60_bht; // @[branch_predictor.scala 30:22]
  reg  btb_61_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_61_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_61_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_61_bht; // @[branch_predictor.scala 30:22]
  reg  btb_62_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_62_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_62_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_62_bht; // @[branch_predictor.scala 30:22]
  reg  btb_63_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_63_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_63_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_63_bht; // @[branch_predictor.scala 30:22]
  reg  btb_64_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_64_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_64_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_64_bht; // @[branch_predictor.scala 30:22]
  reg  btb_65_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_65_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_65_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_65_bht; // @[branch_predictor.scala 30:22]
  reg  btb_66_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_66_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_66_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_66_bht; // @[branch_predictor.scala 30:22]
  reg  btb_67_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_67_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_67_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_67_bht; // @[branch_predictor.scala 30:22]
  reg  btb_68_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_68_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_68_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_68_bht; // @[branch_predictor.scala 30:22]
  reg  btb_69_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_69_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_69_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_69_bht; // @[branch_predictor.scala 30:22]
  reg  btb_70_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_70_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_70_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_70_bht; // @[branch_predictor.scala 30:22]
  reg  btb_71_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_71_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_71_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_71_bht; // @[branch_predictor.scala 30:22]
  reg  btb_72_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_72_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_72_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_72_bht; // @[branch_predictor.scala 30:22]
  reg  btb_73_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_73_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_73_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_73_bht; // @[branch_predictor.scala 30:22]
  reg  btb_74_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_74_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_74_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_74_bht; // @[branch_predictor.scala 30:22]
  reg  btb_75_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_75_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_75_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_75_bht; // @[branch_predictor.scala 30:22]
  reg  btb_76_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_76_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_76_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_76_bht; // @[branch_predictor.scala 30:22]
  reg  btb_77_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_77_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_77_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_77_bht; // @[branch_predictor.scala 30:22]
  reg  btb_78_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_78_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_78_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_78_bht; // @[branch_predictor.scala 30:22]
  reg  btb_79_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_79_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_79_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_79_bht; // @[branch_predictor.scala 30:22]
  reg  btb_80_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_80_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_80_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_80_bht; // @[branch_predictor.scala 30:22]
  reg  btb_81_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_81_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_81_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_81_bht; // @[branch_predictor.scala 30:22]
  reg  btb_82_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_82_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_82_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_82_bht; // @[branch_predictor.scala 30:22]
  reg  btb_83_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_83_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_83_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_83_bht; // @[branch_predictor.scala 30:22]
  reg  btb_84_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_84_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_84_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_84_bht; // @[branch_predictor.scala 30:22]
  reg  btb_85_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_85_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_85_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_85_bht; // @[branch_predictor.scala 30:22]
  reg  btb_86_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_86_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_86_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_86_bht; // @[branch_predictor.scala 30:22]
  reg  btb_87_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_87_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_87_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_87_bht; // @[branch_predictor.scala 30:22]
  reg  btb_88_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_88_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_88_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_88_bht; // @[branch_predictor.scala 30:22]
  reg  btb_89_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_89_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_89_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_89_bht; // @[branch_predictor.scala 30:22]
  reg  btb_90_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_90_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_90_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_90_bht; // @[branch_predictor.scala 30:22]
  reg  btb_91_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_91_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_91_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_91_bht; // @[branch_predictor.scala 30:22]
  reg  btb_92_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_92_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_92_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_92_bht; // @[branch_predictor.scala 30:22]
  reg  btb_93_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_93_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_93_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_93_bht; // @[branch_predictor.scala 30:22]
  reg  btb_94_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_94_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_94_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_94_bht; // @[branch_predictor.scala 30:22]
  reg  btb_95_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_95_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_95_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_95_bht; // @[branch_predictor.scala 30:22]
  reg  btb_96_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_96_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_96_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_96_bht; // @[branch_predictor.scala 30:22]
  reg  btb_97_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_97_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_97_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_97_bht; // @[branch_predictor.scala 30:22]
  reg  btb_98_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_98_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_98_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_98_bht; // @[branch_predictor.scala 30:22]
  reg  btb_99_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_99_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_99_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_99_bht; // @[branch_predictor.scala 30:22]
  reg  btb_100_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_100_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_100_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_100_bht; // @[branch_predictor.scala 30:22]
  reg  btb_101_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_101_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_101_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_101_bht; // @[branch_predictor.scala 30:22]
  reg  btb_102_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_102_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_102_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_102_bht; // @[branch_predictor.scala 30:22]
  reg  btb_103_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_103_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_103_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_103_bht; // @[branch_predictor.scala 30:22]
  reg  btb_104_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_104_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_104_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_104_bht; // @[branch_predictor.scala 30:22]
  reg  btb_105_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_105_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_105_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_105_bht; // @[branch_predictor.scala 30:22]
  reg  btb_106_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_106_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_106_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_106_bht; // @[branch_predictor.scala 30:22]
  reg  btb_107_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_107_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_107_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_107_bht; // @[branch_predictor.scala 30:22]
  reg  btb_108_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_108_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_108_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_108_bht; // @[branch_predictor.scala 30:22]
  reg  btb_109_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_109_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_109_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_109_bht; // @[branch_predictor.scala 30:22]
  reg  btb_110_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_110_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_110_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_110_bht; // @[branch_predictor.scala 30:22]
  reg  btb_111_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_111_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_111_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_111_bht; // @[branch_predictor.scala 30:22]
  reg  btb_112_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_112_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_112_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_112_bht; // @[branch_predictor.scala 30:22]
  reg  btb_113_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_113_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_113_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_113_bht; // @[branch_predictor.scala 30:22]
  reg  btb_114_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_114_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_114_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_114_bht; // @[branch_predictor.scala 30:22]
  reg  btb_115_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_115_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_115_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_115_bht; // @[branch_predictor.scala 30:22]
  reg  btb_116_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_116_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_116_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_116_bht; // @[branch_predictor.scala 30:22]
  reg  btb_117_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_117_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_117_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_117_bht; // @[branch_predictor.scala 30:22]
  reg  btb_118_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_118_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_118_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_118_bht; // @[branch_predictor.scala 30:22]
  reg  btb_119_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_119_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_119_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_119_bht; // @[branch_predictor.scala 30:22]
  reg  btb_120_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_120_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_120_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_120_bht; // @[branch_predictor.scala 30:22]
  reg  btb_121_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_121_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_121_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_121_bht; // @[branch_predictor.scala 30:22]
  reg  btb_122_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_122_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_122_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_122_bht; // @[branch_predictor.scala 30:22]
  reg  btb_123_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_123_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_123_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_123_bht; // @[branch_predictor.scala 30:22]
  reg  btb_124_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_124_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_124_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_124_bht; // @[branch_predictor.scala 30:22]
  reg  btb_125_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_125_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_125_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_125_bht; // @[branch_predictor.scala 30:22]
  reg  btb_126_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_126_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_126_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_126_bht; // @[branch_predictor.scala 30:22]
  reg  btb_127_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_127_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_127_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_127_bht; // @[branch_predictor.scala 30:22]
  reg  btb_128_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_128_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_128_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_128_bht; // @[branch_predictor.scala 30:22]
  reg  btb_129_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_129_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_129_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_129_bht; // @[branch_predictor.scala 30:22]
  reg  btb_130_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_130_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_130_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_130_bht; // @[branch_predictor.scala 30:22]
  reg  btb_131_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_131_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_131_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_131_bht; // @[branch_predictor.scala 30:22]
  reg  btb_132_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_132_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_132_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_132_bht; // @[branch_predictor.scala 30:22]
  reg  btb_133_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_133_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_133_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_133_bht; // @[branch_predictor.scala 30:22]
  reg  btb_134_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_134_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_134_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_134_bht; // @[branch_predictor.scala 30:22]
  reg  btb_135_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_135_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_135_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_135_bht; // @[branch_predictor.scala 30:22]
  reg  btb_136_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_136_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_136_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_136_bht; // @[branch_predictor.scala 30:22]
  reg  btb_137_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_137_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_137_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_137_bht; // @[branch_predictor.scala 30:22]
  reg  btb_138_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_138_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_138_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_138_bht; // @[branch_predictor.scala 30:22]
  reg  btb_139_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_139_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_139_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_139_bht; // @[branch_predictor.scala 30:22]
  reg  btb_140_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_140_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_140_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_140_bht; // @[branch_predictor.scala 30:22]
  reg  btb_141_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_141_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_141_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_141_bht; // @[branch_predictor.scala 30:22]
  reg  btb_142_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_142_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_142_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_142_bht; // @[branch_predictor.scala 30:22]
  reg  btb_143_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_143_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_143_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_143_bht; // @[branch_predictor.scala 30:22]
  reg  btb_144_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_144_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_144_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_144_bht; // @[branch_predictor.scala 30:22]
  reg  btb_145_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_145_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_145_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_145_bht; // @[branch_predictor.scala 30:22]
  reg  btb_146_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_146_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_146_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_146_bht; // @[branch_predictor.scala 30:22]
  reg  btb_147_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_147_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_147_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_147_bht; // @[branch_predictor.scala 30:22]
  reg  btb_148_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_148_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_148_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_148_bht; // @[branch_predictor.scala 30:22]
  reg  btb_149_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_149_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_149_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_149_bht; // @[branch_predictor.scala 30:22]
  reg  btb_150_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_150_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_150_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_150_bht; // @[branch_predictor.scala 30:22]
  reg  btb_151_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_151_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_151_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_151_bht; // @[branch_predictor.scala 30:22]
  reg  btb_152_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_152_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_152_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_152_bht; // @[branch_predictor.scala 30:22]
  reg  btb_153_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_153_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_153_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_153_bht; // @[branch_predictor.scala 30:22]
  reg  btb_154_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_154_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_154_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_154_bht; // @[branch_predictor.scala 30:22]
  reg  btb_155_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_155_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_155_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_155_bht; // @[branch_predictor.scala 30:22]
  reg  btb_156_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_156_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_156_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_156_bht; // @[branch_predictor.scala 30:22]
  reg  btb_157_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_157_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_157_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_157_bht; // @[branch_predictor.scala 30:22]
  reg  btb_158_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_158_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_158_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_158_bht; // @[branch_predictor.scala 30:22]
  reg  btb_159_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_159_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_159_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_159_bht; // @[branch_predictor.scala 30:22]
  reg  btb_160_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_160_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_160_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_160_bht; // @[branch_predictor.scala 30:22]
  reg  btb_161_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_161_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_161_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_161_bht; // @[branch_predictor.scala 30:22]
  reg  btb_162_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_162_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_162_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_162_bht; // @[branch_predictor.scala 30:22]
  reg  btb_163_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_163_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_163_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_163_bht; // @[branch_predictor.scala 30:22]
  reg  btb_164_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_164_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_164_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_164_bht; // @[branch_predictor.scala 30:22]
  reg  btb_165_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_165_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_165_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_165_bht; // @[branch_predictor.scala 30:22]
  reg  btb_166_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_166_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_166_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_166_bht; // @[branch_predictor.scala 30:22]
  reg  btb_167_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_167_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_167_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_167_bht; // @[branch_predictor.scala 30:22]
  reg  btb_168_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_168_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_168_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_168_bht; // @[branch_predictor.scala 30:22]
  reg  btb_169_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_169_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_169_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_169_bht; // @[branch_predictor.scala 30:22]
  reg  btb_170_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_170_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_170_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_170_bht; // @[branch_predictor.scala 30:22]
  reg  btb_171_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_171_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_171_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_171_bht; // @[branch_predictor.scala 30:22]
  reg  btb_172_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_172_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_172_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_172_bht; // @[branch_predictor.scala 30:22]
  reg  btb_173_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_173_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_173_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_173_bht; // @[branch_predictor.scala 30:22]
  reg  btb_174_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_174_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_174_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_174_bht; // @[branch_predictor.scala 30:22]
  reg  btb_175_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_175_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_175_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_175_bht; // @[branch_predictor.scala 30:22]
  reg  btb_176_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_176_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_176_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_176_bht; // @[branch_predictor.scala 30:22]
  reg  btb_177_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_177_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_177_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_177_bht; // @[branch_predictor.scala 30:22]
  reg  btb_178_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_178_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_178_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_178_bht; // @[branch_predictor.scala 30:22]
  reg  btb_179_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_179_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_179_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_179_bht; // @[branch_predictor.scala 30:22]
  reg  btb_180_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_180_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_180_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_180_bht; // @[branch_predictor.scala 30:22]
  reg  btb_181_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_181_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_181_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_181_bht; // @[branch_predictor.scala 30:22]
  reg  btb_182_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_182_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_182_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_182_bht; // @[branch_predictor.scala 30:22]
  reg  btb_183_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_183_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_183_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_183_bht; // @[branch_predictor.scala 30:22]
  reg  btb_184_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_184_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_184_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_184_bht; // @[branch_predictor.scala 30:22]
  reg  btb_185_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_185_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_185_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_185_bht; // @[branch_predictor.scala 30:22]
  reg  btb_186_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_186_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_186_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_186_bht; // @[branch_predictor.scala 30:22]
  reg  btb_187_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_187_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_187_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_187_bht; // @[branch_predictor.scala 30:22]
  reg  btb_188_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_188_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_188_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_188_bht; // @[branch_predictor.scala 30:22]
  reg  btb_189_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_189_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_189_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_189_bht; // @[branch_predictor.scala 30:22]
  reg  btb_190_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_190_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_190_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_190_bht; // @[branch_predictor.scala 30:22]
  reg  btb_191_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_191_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_191_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_191_bht; // @[branch_predictor.scala 30:22]
  reg  btb_192_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_192_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_192_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_192_bht; // @[branch_predictor.scala 30:22]
  reg  btb_193_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_193_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_193_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_193_bht; // @[branch_predictor.scala 30:22]
  reg  btb_194_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_194_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_194_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_194_bht; // @[branch_predictor.scala 30:22]
  reg  btb_195_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_195_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_195_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_195_bht; // @[branch_predictor.scala 30:22]
  reg  btb_196_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_196_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_196_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_196_bht; // @[branch_predictor.scala 30:22]
  reg  btb_197_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_197_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_197_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_197_bht; // @[branch_predictor.scala 30:22]
  reg  btb_198_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_198_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_198_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_198_bht; // @[branch_predictor.scala 30:22]
  reg  btb_199_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_199_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_199_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_199_bht; // @[branch_predictor.scala 30:22]
  reg  btb_200_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_200_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_200_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_200_bht; // @[branch_predictor.scala 30:22]
  reg  btb_201_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_201_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_201_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_201_bht; // @[branch_predictor.scala 30:22]
  reg  btb_202_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_202_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_202_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_202_bht; // @[branch_predictor.scala 30:22]
  reg  btb_203_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_203_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_203_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_203_bht; // @[branch_predictor.scala 30:22]
  reg  btb_204_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_204_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_204_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_204_bht; // @[branch_predictor.scala 30:22]
  reg  btb_205_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_205_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_205_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_205_bht; // @[branch_predictor.scala 30:22]
  reg  btb_206_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_206_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_206_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_206_bht; // @[branch_predictor.scala 30:22]
  reg  btb_207_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_207_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_207_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_207_bht; // @[branch_predictor.scala 30:22]
  reg  btb_208_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_208_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_208_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_208_bht; // @[branch_predictor.scala 30:22]
  reg  btb_209_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_209_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_209_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_209_bht; // @[branch_predictor.scala 30:22]
  reg  btb_210_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_210_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_210_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_210_bht; // @[branch_predictor.scala 30:22]
  reg  btb_211_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_211_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_211_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_211_bht; // @[branch_predictor.scala 30:22]
  reg  btb_212_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_212_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_212_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_212_bht; // @[branch_predictor.scala 30:22]
  reg  btb_213_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_213_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_213_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_213_bht; // @[branch_predictor.scala 30:22]
  reg  btb_214_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_214_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_214_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_214_bht; // @[branch_predictor.scala 30:22]
  reg  btb_215_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_215_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_215_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_215_bht; // @[branch_predictor.scala 30:22]
  reg  btb_216_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_216_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_216_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_216_bht; // @[branch_predictor.scala 30:22]
  reg  btb_217_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_217_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_217_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_217_bht; // @[branch_predictor.scala 30:22]
  reg  btb_218_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_218_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_218_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_218_bht; // @[branch_predictor.scala 30:22]
  reg  btb_219_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_219_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_219_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_219_bht; // @[branch_predictor.scala 30:22]
  reg  btb_220_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_220_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_220_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_220_bht; // @[branch_predictor.scala 30:22]
  reg  btb_221_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_221_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_221_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_221_bht; // @[branch_predictor.scala 30:22]
  reg  btb_222_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_222_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_222_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_222_bht; // @[branch_predictor.scala 30:22]
  reg  btb_223_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_223_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_223_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_223_bht; // @[branch_predictor.scala 30:22]
  reg  btb_224_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_224_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_224_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_224_bht; // @[branch_predictor.scala 30:22]
  reg  btb_225_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_225_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_225_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_225_bht; // @[branch_predictor.scala 30:22]
  reg  btb_226_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_226_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_226_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_226_bht; // @[branch_predictor.scala 30:22]
  reg  btb_227_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_227_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_227_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_227_bht; // @[branch_predictor.scala 30:22]
  reg  btb_228_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_228_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_228_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_228_bht; // @[branch_predictor.scala 30:22]
  reg  btb_229_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_229_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_229_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_229_bht; // @[branch_predictor.scala 30:22]
  reg  btb_230_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_230_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_230_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_230_bht; // @[branch_predictor.scala 30:22]
  reg  btb_231_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_231_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_231_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_231_bht; // @[branch_predictor.scala 30:22]
  reg  btb_232_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_232_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_232_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_232_bht; // @[branch_predictor.scala 30:22]
  reg  btb_233_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_233_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_233_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_233_bht; // @[branch_predictor.scala 30:22]
  reg  btb_234_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_234_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_234_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_234_bht; // @[branch_predictor.scala 30:22]
  reg  btb_235_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_235_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_235_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_235_bht; // @[branch_predictor.scala 30:22]
  reg  btb_236_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_236_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_236_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_236_bht; // @[branch_predictor.scala 30:22]
  reg  btb_237_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_237_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_237_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_237_bht; // @[branch_predictor.scala 30:22]
  reg  btb_238_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_238_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_238_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_238_bht; // @[branch_predictor.scala 30:22]
  reg  btb_239_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_239_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_239_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_239_bht; // @[branch_predictor.scala 30:22]
  reg  btb_240_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_240_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_240_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_240_bht; // @[branch_predictor.scala 30:22]
  reg  btb_241_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_241_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_241_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_241_bht; // @[branch_predictor.scala 30:22]
  reg  btb_242_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_242_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_242_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_242_bht; // @[branch_predictor.scala 30:22]
  reg  btb_243_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_243_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_243_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_243_bht; // @[branch_predictor.scala 30:22]
  reg  btb_244_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_244_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_244_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_244_bht; // @[branch_predictor.scala 30:22]
  reg  btb_245_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_245_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_245_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_245_bht; // @[branch_predictor.scala 30:22]
  reg  btb_246_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_246_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_246_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_246_bht; // @[branch_predictor.scala 30:22]
  reg  btb_247_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_247_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_247_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_247_bht; // @[branch_predictor.scala 30:22]
  reg  btb_248_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_248_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_248_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_248_bht; // @[branch_predictor.scala 30:22]
  reg  btb_249_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_249_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_249_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_249_bht; // @[branch_predictor.scala 30:22]
  reg  btb_250_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_250_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_250_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_250_bht; // @[branch_predictor.scala 30:22]
  reg  btb_251_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_251_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_251_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_251_bht; // @[branch_predictor.scala 30:22]
  reg  btb_252_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_252_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_252_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_252_bht; // @[branch_predictor.scala 30:22]
  reg  btb_253_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_253_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_253_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_253_bht; // @[branch_predictor.scala 30:22]
  reg  btb_254_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_254_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_254_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_254_bht; // @[branch_predictor.scala 30:22]
  reg  btb_255_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_255_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_255_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_255_bht; // @[branch_predictor.scala 30:22]
  reg  btb_256_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_256_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_256_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_256_bht; // @[branch_predictor.scala 30:22]
  reg  btb_257_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_257_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_257_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_257_bht; // @[branch_predictor.scala 30:22]
  reg  btb_258_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_258_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_258_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_258_bht; // @[branch_predictor.scala 30:22]
  reg  btb_259_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_259_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_259_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_259_bht; // @[branch_predictor.scala 30:22]
  reg  btb_260_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_260_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_260_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_260_bht; // @[branch_predictor.scala 30:22]
  reg  btb_261_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_261_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_261_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_261_bht; // @[branch_predictor.scala 30:22]
  reg  btb_262_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_262_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_262_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_262_bht; // @[branch_predictor.scala 30:22]
  reg  btb_263_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_263_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_263_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_263_bht; // @[branch_predictor.scala 30:22]
  reg  btb_264_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_264_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_264_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_264_bht; // @[branch_predictor.scala 30:22]
  reg  btb_265_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_265_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_265_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_265_bht; // @[branch_predictor.scala 30:22]
  reg  btb_266_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_266_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_266_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_266_bht; // @[branch_predictor.scala 30:22]
  reg  btb_267_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_267_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_267_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_267_bht; // @[branch_predictor.scala 30:22]
  reg  btb_268_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_268_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_268_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_268_bht; // @[branch_predictor.scala 30:22]
  reg  btb_269_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_269_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_269_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_269_bht; // @[branch_predictor.scala 30:22]
  reg  btb_270_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_270_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_270_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_270_bht; // @[branch_predictor.scala 30:22]
  reg  btb_271_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_271_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_271_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_271_bht; // @[branch_predictor.scala 30:22]
  reg  btb_272_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_272_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_272_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_272_bht; // @[branch_predictor.scala 30:22]
  reg  btb_273_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_273_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_273_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_273_bht; // @[branch_predictor.scala 30:22]
  reg  btb_274_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_274_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_274_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_274_bht; // @[branch_predictor.scala 30:22]
  reg  btb_275_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_275_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_275_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_275_bht; // @[branch_predictor.scala 30:22]
  reg  btb_276_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_276_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_276_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_276_bht; // @[branch_predictor.scala 30:22]
  reg  btb_277_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_277_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_277_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_277_bht; // @[branch_predictor.scala 30:22]
  reg  btb_278_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_278_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_278_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_278_bht; // @[branch_predictor.scala 30:22]
  reg  btb_279_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_279_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_279_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_279_bht; // @[branch_predictor.scala 30:22]
  reg  btb_280_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_280_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_280_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_280_bht; // @[branch_predictor.scala 30:22]
  reg  btb_281_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_281_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_281_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_281_bht; // @[branch_predictor.scala 30:22]
  reg  btb_282_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_282_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_282_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_282_bht; // @[branch_predictor.scala 30:22]
  reg  btb_283_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_283_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_283_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_283_bht; // @[branch_predictor.scala 30:22]
  reg  btb_284_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_284_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_284_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_284_bht; // @[branch_predictor.scala 30:22]
  reg  btb_285_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_285_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_285_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_285_bht; // @[branch_predictor.scala 30:22]
  reg  btb_286_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_286_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_286_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_286_bht; // @[branch_predictor.scala 30:22]
  reg  btb_287_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_287_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_287_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_287_bht; // @[branch_predictor.scala 30:22]
  reg  btb_288_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_288_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_288_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_288_bht; // @[branch_predictor.scala 30:22]
  reg  btb_289_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_289_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_289_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_289_bht; // @[branch_predictor.scala 30:22]
  reg  btb_290_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_290_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_290_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_290_bht; // @[branch_predictor.scala 30:22]
  reg  btb_291_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_291_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_291_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_291_bht; // @[branch_predictor.scala 30:22]
  reg  btb_292_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_292_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_292_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_292_bht; // @[branch_predictor.scala 30:22]
  reg  btb_293_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_293_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_293_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_293_bht; // @[branch_predictor.scala 30:22]
  reg  btb_294_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_294_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_294_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_294_bht; // @[branch_predictor.scala 30:22]
  reg  btb_295_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_295_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_295_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_295_bht; // @[branch_predictor.scala 30:22]
  reg  btb_296_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_296_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_296_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_296_bht; // @[branch_predictor.scala 30:22]
  reg  btb_297_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_297_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_297_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_297_bht; // @[branch_predictor.scala 30:22]
  reg  btb_298_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_298_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_298_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_298_bht; // @[branch_predictor.scala 30:22]
  reg  btb_299_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_299_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_299_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_299_bht; // @[branch_predictor.scala 30:22]
  reg  btb_300_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_300_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_300_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_300_bht; // @[branch_predictor.scala 30:22]
  reg  btb_301_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_301_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_301_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_301_bht; // @[branch_predictor.scala 30:22]
  reg  btb_302_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_302_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_302_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_302_bht; // @[branch_predictor.scala 30:22]
  reg  btb_303_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_303_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_303_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_303_bht; // @[branch_predictor.scala 30:22]
  reg  btb_304_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_304_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_304_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_304_bht; // @[branch_predictor.scala 30:22]
  reg  btb_305_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_305_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_305_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_305_bht; // @[branch_predictor.scala 30:22]
  reg  btb_306_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_306_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_306_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_306_bht; // @[branch_predictor.scala 30:22]
  reg  btb_307_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_307_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_307_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_307_bht; // @[branch_predictor.scala 30:22]
  reg  btb_308_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_308_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_308_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_308_bht; // @[branch_predictor.scala 30:22]
  reg  btb_309_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_309_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_309_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_309_bht; // @[branch_predictor.scala 30:22]
  reg  btb_310_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_310_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_310_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_310_bht; // @[branch_predictor.scala 30:22]
  reg  btb_311_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_311_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_311_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_311_bht; // @[branch_predictor.scala 30:22]
  reg  btb_312_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_312_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_312_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_312_bht; // @[branch_predictor.scala 30:22]
  reg  btb_313_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_313_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_313_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_313_bht; // @[branch_predictor.scala 30:22]
  reg  btb_314_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_314_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_314_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_314_bht; // @[branch_predictor.scala 30:22]
  reg  btb_315_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_315_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_315_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_315_bht; // @[branch_predictor.scala 30:22]
  reg  btb_316_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_316_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_316_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_316_bht; // @[branch_predictor.scala 30:22]
  reg  btb_317_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_317_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_317_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_317_bht; // @[branch_predictor.scala 30:22]
  reg  btb_318_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_318_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_318_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_318_bht; // @[branch_predictor.scala 30:22]
  reg  btb_319_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_319_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_319_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_319_bht; // @[branch_predictor.scala 30:22]
  reg  btb_320_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_320_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_320_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_320_bht; // @[branch_predictor.scala 30:22]
  reg  btb_321_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_321_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_321_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_321_bht; // @[branch_predictor.scala 30:22]
  reg  btb_322_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_322_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_322_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_322_bht; // @[branch_predictor.scala 30:22]
  reg  btb_323_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_323_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_323_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_323_bht; // @[branch_predictor.scala 30:22]
  reg  btb_324_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_324_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_324_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_324_bht; // @[branch_predictor.scala 30:22]
  reg  btb_325_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_325_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_325_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_325_bht; // @[branch_predictor.scala 30:22]
  reg  btb_326_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_326_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_326_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_326_bht; // @[branch_predictor.scala 30:22]
  reg  btb_327_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_327_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_327_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_327_bht; // @[branch_predictor.scala 30:22]
  reg  btb_328_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_328_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_328_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_328_bht; // @[branch_predictor.scala 30:22]
  reg  btb_329_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_329_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_329_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_329_bht; // @[branch_predictor.scala 30:22]
  reg  btb_330_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_330_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_330_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_330_bht; // @[branch_predictor.scala 30:22]
  reg  btb_331_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_331_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_331_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_331_bht; // @[branch_predictor.scala 30:22]
  reg  btb_332_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_332_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_332_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_332_bht; // @[branch_predictor.scala 30:22]
  reg  btb_333_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_333_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_333_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_333_bht; // @[branch_predictor.scala 30:22]
  reg  btb_334_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_334_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_334_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_334_bht; // @[branch_predictor.scala 30:22]
  reg  btb_335_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_335_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_335_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_335_bht; // @[branch_predictor.scala 30:22]
  reg  btb_336_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_336_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_336_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_336_bht; // @[branch_predictor.scala 30:22]
  reg  btb_337_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_337_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_337_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_337_bht; // @[branch_predictor.scala 30:22]
  reg  btb_338_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_338_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_338_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_338_bht; // @[branch_predictor.scala 30:22]
  reg  btb_339_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_339_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_339_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_339_bht; // @[branch_predictor.scala 30:22]
  reg  btb_340_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_340_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_340_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_340_bht; // @[branch_predictor.scala 30:22]
  reg  btb_341_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_341_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_341_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_341_bht; // @[branch_predictor.scala 30:22]
  reg  btb_342_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_342_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_342_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_342_bht; // @[branch_predictor.scala 30:22]
  reg  btb_343_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_343_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_343_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_343_bht; // @[branch_predictor.scala 30:22]
  reg  btb_344_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_344_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_344_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_344_bht; // @[branch_predictor.scala 30:22]
  reg  btb_345_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_345_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_345_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_345_bht; // @[branch_predictor.scala 30:22]
  reg  btb_346_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_346_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_346_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_346_bht; // @[branch_predictor.scala 30:22]
  reg  btb_347_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_347_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_347_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_347_bht; // @[branch_predictor.scala 30:22]
  reg  btb_348_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_348_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_348_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_348_bht; // @[branch_predictor.scala 30:22]
  reg  btb_349_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_349_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_349_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_349_bht; // @[branch_predictor.scala 30:22]
  reg  btb_350_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_350_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_350_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_350_bht; // @[branch_predictor.scala 30:22]
  reg  btb_351_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_351_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_351_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_351_bht; // @[branch_predictor.scala 30:22]
  reg  btb_352_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_352_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_352_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_352_bht; // @[branch_predictor.scala 30:22]
  reg  btb_353_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_353_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_353_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_353_bht; // @[branch_predictor.scala 30:22]
  reg  btb_354_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_354_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_354_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_354_bht; // @[branch_predictor.scala 30:22]
  reg  btb_355_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_355_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_355_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_355_bht; // @[branch_predictor.scala 30:22]
  reg  btb_356_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_356_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_356_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_356_bht; // @[branch_predictor.scala 30:22]
  reg  btb_357_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_357_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_357_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_357_bht; // @[branch_predictor.scala 30:22]
  reg  btb_358_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_358_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_358_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_358_bht; // @[branch_predictor.scala 30:22]
  reg  btb_359_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_359_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_359_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_359_bht; // @[branch_predictor.scala 30:22]
  reg  btb_360_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_360_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_360_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_360_bht; // @[branch_predictor.scala 30:22]
  reg  btb_361_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_361_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_361_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_361_bht; // @[branch_predictor.scala 30:22]
  reg  btb_362_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_362_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_362_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_362_bht; // @[branch_predictor.scala 30:22]
  reg  btb_363_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_363_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_363_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_363_bht; // @[branch_predictor.scala 30:22]
  reg  btb_364_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_364_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_364_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_364_bht; // @[branch_predictor.scala 30:22]
  reg  btb_365_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_365_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_365_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_365_bht; // @[branch_predictor.scala 30:22]
  reg  btb_366_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_366_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_366_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_366_bht; // @[branch_predictor.scala 30:22]
  reg  btb_367_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_367_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_367_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_367_bht; // @[branch_predictor.scala 30:22]
  reg  btb_368_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_368_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_368_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_368_bht; // @[branch_predictor.scala 30:22]
  reg  btb_369_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_369_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_369_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_369_bht; // @[branch_predictor.scala 30:22]
  reg  btb_370_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_370_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_370_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_370_bht; // @[branch_predictor.scala 30:22]
  reg  btb_371_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_371_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_371_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_371_bht; // @[branch_predictor.scala 30:22]
  reg  btb_372_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_372_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_372_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_372_bht; // @[branch_predictor.scala 30:22]
  reg  btb_373_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_373_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_373_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_373_bht; // @[branch_predictor.scala 30:22]
  reg  btb_374_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_374_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_374_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_374_bht; // @[branch_predictor.scala 30:22]
  reg  btb_375_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_375_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_375_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_375_bht; // @[branch_predictor.scala 30:22]
  reg  btb_376_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_376_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_376_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_376_bht; // @[branch_predictor.scala 30:22]
  reg  btb_377_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_377_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_377_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_377_bht; // @[branch_predictor.scala 30:22]
  reg  btb_378_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_378_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_378_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_378_bht; // @[branch_predictor.scala 30:22]
  reg  btb_379_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_379_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_379_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_379_bht; // @[branch_predictor.scala 30:22]
  reg  btb_380_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_380_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_380_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_380_bht; // @[branch_predictor.scala 30:22]
  reg  btb_381_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_381_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_381_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_381_bht; // @[branch_predictor.scala 30:22]
  reg  btb_382_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_382_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_382_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_382_bht; // @[branch_predictor.scala 30:22]
  reg  btb_383_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_383_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_383_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_383_bht; // @[branch_predictor.scala 30:22]
  reg  btb_384_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_384_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_384_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_384_bht; // @[branch_predictor.scala 30:22]
  reg  btb_385_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_385_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_385_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_385_bht; // @[branch_predictor.scala 30:22]
  reg  btb_386_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_386_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_386_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_386_bht; // @[branch_predictor.scala 30:22]
  reg  btb_387_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_387_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_387_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_387_bht; // @[branch_predictor.scala 30:22]
  reg  btb_388_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_388_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_388_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_388_bht; // @[branch_predictor.scala 30:22]
  reg  btb_389_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_389_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_389_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_389_bht; // @[branch_predictor.scala 30:22]
  reg  btb_390_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_390_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_390_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_390_bht; // @[branch_predictor.scala 30:22]
  reg  btb_391_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_391_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_391_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_391_bht; // @[branch_predictor.scala 30:22]
  reg  btb_392_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_392_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_392_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_392_bht; // @[branch_predictor.scala 30:22]
  reg  btb_393_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_393_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_393_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_393_bht; // @[branch_predictor.scala 30:22]
  reg  btb_394_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_394_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_394_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_394_bht; // @[branch_predictor.scala 30:22]
  reg  btb_395_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_395_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_395_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_395_bht; // @[branch_predictor.scala 30:22]
  reg  btb_396_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_396_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_396_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_396_bht; // @[branch_predictor.scala 30:22]
  reg  btb_397_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_397_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_397_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_397_bht; // @[branch_predictor.scala 30:22]
  reg  btb_398_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_398_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_398_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_398_bht; // @[branch_predictor.scala 30:22]
  reg  btb_399_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_399_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_399_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_399_bht; // @[branch_predictor.scala 30:22]
  reg  btb_400_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_400_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_400_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_400_bht; // @[branch_predictor.scala 30:22]
  reg  btb_401_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_401_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_401_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_401_bht; // @[branch_predictor.scala 30:22]
  reg  btb_402_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_402_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_402_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_402_bht; // @[branch_predictor.scala 30:22]
  reg  btb_403_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_403_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_403_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_403_bht; // @[branch_predictor.scala 30:22]
  reg  btb_404_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_404_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_404_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_404_bht; // @[branch_predictor.scala 30:22]
  reg  btb_405_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_405_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_405_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_405_bht; // @[branch_predictor.scala 30:22]
  reg  btb_406_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_406_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_406_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_406_bht; // @[branch_predictor.scala 30:22]
  reg  btb_407_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_407_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_407_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_407_bht; // @[branch_predictor.scala 30:22]
  reg  btb_408_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_408_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_408_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_408_bht; // @[branch_predictor.scala 30:22]
  reg  btb_409_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_409_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_409_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_409_bht; // @[branch_predictor.scala 30:22]
  reg  btb_410_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_410_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_410_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_410_bht; // @[branch_predictor.scala 30:22]
  reg  btb_411_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_411_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_411_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_411_bht; // @[branch_predictor.scala 30:22]
  reg  btb_412_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_412_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_412_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_412_bht; // @[branch_predictor.scala 30:22]
  reg  btb_413_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_413_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_413_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_413_bht; // @[branch_predictor.scala 30:22]
  reg  btb_414_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_414_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_414_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_414_bht; // @[branch_predictor.scala 30:22]
  reg  btb_415_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_415_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_415_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_415_bht; // @[branch_predictor.scala 30:22]
  reg  btb_416_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_416_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_416_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_416_bht; // @[branch_predictor.scala 30:22]
  reg  btb_417_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_417_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_417_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_417_bht; // @[branch_predictor.scala 30:22]
  reg  btb_418_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_418_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_418_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_418_bht; // @[branch_predictor.scala 30:22]
  reg  btb_419_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_419_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_419_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_419_bht; // @[branch_predictor.scala 30:22]
  reg  btb_420_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_420_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_420_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_420_bht; // @[branch_predictor.scala 30:22]
  reg  btb_421_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_421_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_421_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_421_bht; // @[branch_predictor.scala 30:22]
  reg  btb_422_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_422_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_422_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_422_bht; // @[branch_predictor.scala 30:22]
  reg  btb_423_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_423_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_423_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_423_bht; // @[branch_predictor.scala 30:22]
  reg  btb_424_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_424_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_424_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_424_bht; // @[branch_predictor.scala 30:22]
  reg  btb_425_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_425_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_425_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_425_bht; // @[branch_predictor.scala 30:22]
  reg  btb_426_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_426_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_426_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_426_bht; // @[branch_predictor.scala 30:22]
  reg  btb_427_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_427_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_427_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_427_bht; // @[branch_predictor.scala 30:22]
  reg  btb_428_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_428_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_428_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_428_bht; // @[branch_predictor.scala 30:22]
  reg  btb_429_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_429_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_429_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_429_bht; // @[branch_predictor.scala 30:22]
  reg  btb_430_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_430_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_430_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_430_bht; // @[branch_predictor.scala 30:22]
  reg  btb_431_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_431_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_431_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_431_bht; // @[branch_predictor.scala 30:22]
  reg  btb_432_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_432_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_432_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_432_bht; // @[branch_predictor.scala 30:22]
  reg  btb_433_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_433_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_433_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_433_bht; // @[branch_predictor.scala 30:22]
  reg  btb_434_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_434_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_434_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_434_bht; // @[branch_predictor.scala 30:22]
  reg  btb_435_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_435_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_435_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_435_bht; // @[branch_predictor.scala 30:22]
  reg  btb_436_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_436_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_436_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_436_bht; // @[branch_predictor.scala 30:22]
  reg  btb_437_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_437_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_437_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_437_bht; // @[branch_predictor.scala 30:22]
  reg  btb_438_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_438_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_438_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_438_bht; // @[branch_predictor.scala 30:22]
  reg  btb_439_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_439_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_439_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_439_bht; // @[branch_predictor.scala 30:22]
  reg  btb_440_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_440_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_440_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_440_bht; // @[branch_predictor.scala 30:22]
  reg  btb_441_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_441_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_441_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_441_bht; // @[branch_predictor.scala 30:22]
  reg  btb_442_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_442_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_442_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_442_bht; // @[branch_predictor.scala 30:22]
  reg  btb_443_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_443_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_443_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_443_bht; // @[branch_predictor.scala 30:22]
  reg  btb_444_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_444_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_444_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_444_bht; // @[branch_predictor.scala 30:22]
  reg  btb_445_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_445_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_445_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_445_bht; // @[branch_predictor.scala 30:22]
  reg  btb_446_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_446_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_446_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_446_bht; // @[branch_predictor.scala 30:22]
  reg  btb_447_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_447_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_447_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_447_bht; // @[branch_predictor.scala 30:22]
  reg  btb_448_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_448_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_448_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_448_bht; // @[branch_predictor.scala 30:22]
  reg  btb_449_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_449_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_449_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_449_bht; // @[branch_predictor.scala 30:22]
  reg  btb_450_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_450_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_450_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_450_bht; // @[branch_predictor.scala 30:22]
  reg  btb_451_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_451_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_451_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_451_bht; // @[branch_predictor.scala 30:22]
  reg  btb_452_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_452_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_452_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_452_bht; // @[branch_predictor.scala 30:22]
  reg  btb_453_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_453_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_453_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_453_bht; // @[branch_predictor.scala 30:22]
  reg  btb_454_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_454_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_454_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_454_bht; // @[branch_predictor.scala 30:22]
  reg  btb_455_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_455_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_455_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_455_bht; // @[branch_predictor.scala 30:22]
  reg  btb_456_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_456_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_456_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_456_bht; // @[branch_predictor.scala 30:22]
  reg  btb_457_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_457_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_457_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_457_bht; // @[branch_predictor.scala 30:22]
  reg  btb_458_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_458_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_458_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_458_bht; // @[branch_predictor.scala 30:22]
  reg  btb_459_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_459_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_459_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_459_bht; // @[branch_predictor.scala 30:22]
  reg  btb_460_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_460_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_460_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_460_bht; // @[branch_predictor.scala 30:22]
  reg  btb_461_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_461_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_461_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_461_bht; // @[branch_predictor.scala 30:22]
  reg  btb_462_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_462_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_462_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_462_bht; // @[branch_predictor.scala 30:22]
  reg  btb_463_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_463_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_463_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_463_bht; // @[branch_predictor.scala 30:22]
  reg  btb_464_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_464_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_464_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_464_bht; // @[branch_predictor.scala 30:22]
  reg  btb_465_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_465_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_465_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_465_bht; // @[branch_predictor.scala 30:22]
  reg  btb_466_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_466_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_466_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_466_bht; // @[branch_predictor.scala 30:22]
  reg  btb_467_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_467_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_467_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_467_bht; // @[branch_predictor.scala 30:22]
  reg  btb_468_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_468_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_468_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_468_bht; // @[branch_predictor.scala 30:22]
  reg  btb_469_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_469_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_469_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_469_bht; // @[branch_predictor.scala 30:22]
  reg  btb_470_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_470_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_470_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_470_bht; // @[branch_predictor.scala 30:22]
  reg  btb_471_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_471_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_471_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_471_bht; // @[branch_predictor.scala 30:22]
  reg  btb_472_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_472_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_472_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_472_bht; // @[branch_predictor.scala 30:22]
  reg  btb_473_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_473_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_473_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_473_bht; // @[branch_predictor.scala 30:22]
  reg  btb_474_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_474_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_474_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_474_bht; // @[branch_predictor.scala 30:22]
  reg  btb_475_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_475_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_475_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_475_bht; // @[branch_predictor.scala 30:22]
  reg  btb_476_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_476_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_476_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_476_bht; // @[branch_predictor.scala 30:22]
  reg  btb_477_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_477_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_477_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_477_bht; // @[branch_predictor.scala 30:22]
  reg  btb_478_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_478_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_478_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_478_bht; // @[branch_predictor.scala 30:22]
  reg  btb_479_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_479_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_479_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_479_bht; // @[branch_predictor.scala 30:22]
  reg  btb_480_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_480_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_480_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_480_bht; // @[branch_predictor.scala 30:22]
  reg  btb_481_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_481_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_481_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_481_bht; // @[branch_predictor.scala 30:22]
  reg  btb_482_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_482_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_482_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_482_bht; // @[branch_predictor.scala 30:22]
  reg  btb_483_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_483_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_483_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_483_bht; // @[branch_predictor.scala 30:22]
  reg  btb_484_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_484_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_484_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_484_bht; // @[branch_predictor.scala 30:22]
  reg  btb_485_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_485_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_485_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_485_bht; // @[branch_predictor.scala 30:22]
  reg  btb_486_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_486_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_486_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_486_bht; // @[branch_predictor.scala 30:22]
  reg  btb_487_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_487_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_487_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_487_bht; // @[branch_predictor.scala 30:22]
  reg  btb_488_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_488_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_488_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_488_bht; // @[branch_predictor.scala 30:22]
  reg  btb_489_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_489_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_489_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_489_bht; // @[branch_predictor.scala 30:22]
  reg  btb_490_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_490_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_490_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_490_bht; // @[branch_predictor.scala 30:22]
  reg  btb_491_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_491_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_491_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_491_bht; // @[branch_predictor.scala 30:22]
  reg  btb_492_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_492_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_492_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_492_bht; // @[branch_predictor.scala 30:22]
  reg  btb_493_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_493_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_493_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_493_bht; // @[branch_predictor.scala 30:22]
  reg  btb_494_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_494_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_494_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_494_bht; // @[branch_predictor.scala 30:22]
  reg  btb_495_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_495_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_495_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_495_bht; // @[branch_predictor.scala 30:22]
  reg  btb_496_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_496_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_496_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_496_bht; // @[branch_predictor.scala 30:22]
  reg  btb_497_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_497_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_497_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_497_bht; // @[branch_predictor.scala 30:22]
  reg  btb_498_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_498_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_498_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_498_bht; // @[branch_predictor.scala 30:22]
  reg  btb_499_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_499_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_499_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_499_bht; // @[branch_predictor.scala 30:22]
  reg  btb_500_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_500_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_500_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_500_bht; // @[branch_predictor.scala 30:22]
  reg  btb_501_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_501_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_501_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_501_bht; // @[branch_predictor.scala 30:22]
  reg  btb_502_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_502_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_502_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_502_bht; // @[branch_predictor.scala 30:22]
  reg  btb_503_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_503_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_503_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_503_bht; // @[branch_predictor.scala 30:22]
  reg  btb_504_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_504_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_504_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_504_bht; // @[branch_predictor.scala 30:22]
  reg  btb_505_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_505_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_505_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_505_bht; // @[branch_predictor.scala 30:22]
  reg  btb_506_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_506_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_506_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_506_bht; // @[branch_predictor.scala 30:22]
  reg  btb_507_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_507_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_507_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_507_bht; // @[branch_predictor.scala 30:22]
  reg  btb_508_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_508_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_508_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_508_bht; // @[branch_predictor.scala 30:22]
  reg  btb_509_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_509_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_509_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_509_bht; // @[branch_predictor.scala 30:22]
  reg  btb_510_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_510_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_510_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_510_bht; // @[branch_predictor.scala 30:22]
  reg  btb_511_valid; // @[branch_predictor.scala 30:22]
  reg [9:0] btb_511_tag; // @[branch_predictor.scala 30:22]
  reg [63:0] btb_511_target_address; // @[branch_predictor.scala 30:22]
  reg [1:0] btb_511_bht; // @[branch_predictor.scala 30:22]
  reg [8:0] btb_victim_ptr; // @[branch_predictor.scala 32:33]
  wire  _GEN_0 = btb_0_tag == io_i_addr[12:3] & btb_0_valid; // @[branch_predictor.scala 34:36 40:45 41:44]
  wire [63:0] _GEN_1 = btb_0_tag == io_i_addr[12:3] ? btb_0_target_address : 64'h0; // @[branch_predictor.scala 35:37 40:45 42:45]
  wire  _GEN_4 = btb_0_tag == io_i_addr[12:3] & ~btb_0_bht[1]; // @[branch_predictor.scala 38:36 40:45 45:44]
  wire  _GEN_5 = btb_1_tag == io_i_addr[12:3] ? btb_1_valid : _GEN_0; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_6 = btb_1_tag == io_i_addr[12:3] ? btb_1_target_address : _GEN_1; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_9 = btb_1_tag == io_i_addr[12:3] ? ~btb_1_bht[1] : _GEN_4; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_10 = btb_2_tag == io_i_addr[12:3] ? btb_2_valid : _GEN_5; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_11 = btb_2_tag == io_i_addr[12:3] ? btb_2_target_address : _GEN_6; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_14 = btb_2_tag == io_i_addr[12:3] ? ~btb_2_bht[1] : _GEN_9; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_15 = btb_3_tag == io_i_addr[12:3] ? btb_3_valid : _GEN_10; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_16 = btb_3_tag == io_i_addr[12:3] ? btb_3_target_address : _GEN_11; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_19 = btb_3_tag == io_i_addr[12:3] ? ~btb_3_bht[1] : _GEN_14; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_20 = btb_4_tag == io_i_addr[12:3] ? btb_4_valid : _GEN_15; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_21 = btb_4_tag == io_i_addr[12:3] ? btb_4_target_address : _GEN_16; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_24 = btb_4_tag == io_i_addr[12:3] ? ~btb_4_bht[1] : _GEN_19; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_25 = btb_5_tag == io_i_addr[12:3] ? btb_5_valid : _GEN_20; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_26 = btb_5_tag == io_i_addr[12:3] ? btb_5_target_address : _GEN_21; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_29 = btb_5_tag == io_i_addr[12:3] ? ~btb_5_bht[1] : _GEN_24; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_30 = btb_6_tag == io_i_addr[12:3] ? btb_6_valid : _GEN_25; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_31 = btb_6_tag == io_i_addr[12:3] ? btb_6_target_address : _GEN_26; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_34 = btb_6_tag == io_i_addr[12:3] ? ~btb_6_bht[1] : _GEN_29; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_35 = btb_7_tag == io_i_addr[12:3] ? btb_7_valid : _GEN_30; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_36 = btb_7_tag == io_i_addr[12:3] ? btb_7_target_address : _GEN_31; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_39 = btb_7_tag == io_i_addr[12:3] ? ~btb_7_bht[1] : _GEN_34; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_40 = btb_8_tag == io_i_addr[12:3] ? btb_8_valid : _GEN_35; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_41 = btb_8_tag == io_i_addr[12:3] ? btb_8_target_address : _GEN_36; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_44 = btb_8_tag == io_i_addr[12:3] ? ~btb_8_bht[1] : _GEN_39; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_45 = btb_9_tag == io_i_addr[12:3] ? btb_9_valid : _GEN_40; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_46 = btb_9_tag == io_i_addr[12:3] ? btb_9_target_address : _GEN_41; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_49 = btb_9_tag == io_i_addr[12:3] ? ~btb_9_bht[1] : _GEN_44; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_50 = btb_10_tag == io_i_addr[12:3] ? btb_10_valid : _GEN_45; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_51 = btb_10_tag == io_i_addr[12:3] ? btb_10_target_address : _GEN_46; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_54 = btb_10_tag == io_i_addr[12:3] ? ~btb_10_bht[1] : _GEN_49; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_55 = btb_11_tag == io_i_addr[12:3] ? btb_11_valid : _GEN_50; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_56 = btb_11_tag == io_i_addr[12:3] ? btb_11_target_address : _GEN_51; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_59 = btb_11_tag == io_i_addr[12:3] ? ~btb_11_bht[1] : _GEN_54; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_60 = btb_12_tag == io_i_addr[12:3] ? btb_12_valid : _GEN_55; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_61 = btb_12_tag == io_i_addr[12:3] ? btb_12_target_address : _GEN_56; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_64 = btb_12_tag == io_i_addr[12:3] ? ~btb_12_bht[1] : _GEN_59; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_65 = btb_13_tag == io_i_addr[12:3] ? btb_13_valid : _GEN_60; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_66 = btb_13_tag == io_i_addr[12:3] ? btb_13_target_address : _GEN_61; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_69 = btb_13_tag == io_i_addr[12:3] ? ~btb_13_bht[1] : _GEN_64; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_70 = btb_14_tag == io_i_addr[12:3] ? btb_14_valid : _GEN_65; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_71 = btb_14_tag == io_i_addr[12:3] ? btb_14_target_address : _GEN_66; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_74 = btb_14_tag == io_i_addr[12:3] ? ~btb_14_bht[1] : _GEN_69; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_75 = btb_15_tag == io_i_addr[12:3] ? btb_15_valid : _GEN_70; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_76 = btb_15_tag == io_i_addr[12:3] ? btb_15_target_address : _GEN_71; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_79 = btb_15_tag == io_i_addr[12:3] ? ~btb_15_bht[1] : _GEN_74; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_80 = btb_16_tag == io_i_addr[12:3] ? btb_16_valid : _GEN_75; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_81 = btb_16_tag == io_i_addr[12:3] ? btb_16_target_address : _GEN_76; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_84 = btb_16_tag == io_i_addr[12:3] ? ~btb_16_bht[1] : _GEN_79; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_85 = btb_17_tag == io_i_addr[12:3] ? btb_17_valid : _GEN_80; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_86 = btb_17_tag == io_i_addr[12:3] ? btb_17_target_address : _GEN_81; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_89 = btb_17_tag == io_i_addr[12:3] ? ~btb_17_bht[1] : _GEN_84; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_90 = btb_18_tag == io_i_addr[12:3] ? btb_18_valid : _GEN_85; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_91 = btb_18_tag == io_i_addr[12:3] ? btb_18_target_address : _GEN_86; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_94 = btb_18_tag == io_i_addr[12:3] ? ~btb_18_bht[1] : _GEN_89; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_95 = btb_19_tag == io_i_addr[12:3] ? btb_19_valid : _GEN_90; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_96 = btb_19_tag == io_i_addr[12:3] ? btb_19_target_address : _GEN_91; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_99 = btb_19_tag == io_i_addr[12:3] ? ~btb_19_bht[1] : _GEN_94; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_100 = btb_20_tag == io_i_addr[12:3] ? btb_20_valid : _GEN_95; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_101 = btb_20_tag == io_i_addr[12:3] ? btb_20_target_address : _GEN_96; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_104 = btb_20_tag == io_i_addr[12:3] ? ~btb_20_bht[1] : _GEN_99; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_105 = btb_21_tag == io_i_addr[12:3] ? btb_21_valid : _GEN_100; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_106 = btb_21_tag == io_i_addr[12:3] ? btb_21_target_address : _GEN_101; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_109 = btb_21_tag == io_i_addr[12:3] ? ~btb_21_bht[1] : _GEN_104; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_110 = btb_22_tag == io_i_addr[12:3] ? btb_22_valid : _GEN_105; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_111 = btb_22_tag == io_i_addr[12:3] ? btb_22_target_address : _GEN_106; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_114 = btb_22_tag == io_i_addr[12:3] ? ~btb_22_bht[1] : _GEN_109; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_115 = btb_23_tag == io_i_addr[12:3] ? btb_23_valid : _GEN_110; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_116 = btb_23_tag == io_i_addr[12:3] ? btb_23_target_address : _GEN_111; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_119 = btb_23_tag == io_i_addr[12:3] ? ~btb_23_bht[1] : _GEN_114; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_120 = btb_24_tag == io_i_addr[12:3] ? btb_24_valid : _GEN_115; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_121 = btb_24_tag == io_i_addr[12:3] ? btb_24_target_address : _GEN_116; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_124 = btb_24_tag == io_i_addr[12:3] ? ~btb_24_bht[1] : _GEN_119; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_125 = btb_25_tag == io_i_addr[12:3] ? btb_25_valid : _GEN_120; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_126 = btb_25_tag == io_i_addr[12:3] ? btb_25_target_address : _GEN_121; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_129 = btb_25_tag == io_i_addr[12:3] ? ~btb_25_bht[1] : _GEN_124; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_130 = btb_26_tag == io_i_addr[12:3] ? btb_26_valid : _GEN_125; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_131 = btb_26_tag == io_i_addr[12:3] ? btb_26_target_address : _GEN_126; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_134 = btb_26_tag == io_i_addr[12:3] ? ~btb_26_bht[1] : _GEN_129; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_135 = btb_27_tag == io_i_addr[12:3] ? btb_27_valid : _GEN_130; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_136 = btb_27_tag == io_i_addr[12:3] ? btb_27_target_address : _GEN_131; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_139 = btb_27_tag == io_i_addr[12:3] ? ~btb_27_bht[1] : _GEN_134; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_140 = btb_28_tag == io_i_addr[12:3] ? btb_28_valid : _GEN_135; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_141 = btb_28_tag == io_i_addr[12:3] ? btb_28_target_address : _GEN_136; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_144 = btb_28_tag == io_i_addr[12:3] ? ~btb_28_bht[1] : _GEN_139; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_145 = btb_29_tag == io_i_addr[12:3] ? btb_29_valid : _GEN_140; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_146 = btb_29_tag == io_i_addr[12:3] ? btb_29_target_address : _GEN_141; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_149 = btb_29_tag == io_i_addr[12:3] ? ~btb_29_bht[1] : _GEN_144; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_150 = btb_30_tag == io_i_addr[12:3] ? btb_30_valid : _GEN_145; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_151 = btb_30_tag == io_i_addr[12:3] ? btb_30_target_address : _GEN_146; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_154 = btb_30_tag == io_i_addr[12:3] ? ~btb_30_bht[1] : _GEN_149; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_155 = btb_31_tag == io_i_addr[12:3] ? btb_31_valid : _GEN_150; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_156 = btb_31_tag == io_i_addr[12:3] ? btb_31_target_address : _GEN_151; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_159 = btb_31_tag == io_i_addr[12:3] ? ~btb_31_bht[1] : _GEN_154; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_160 = btb_32_tag == io_i_addr[12:3] ? btb_32_valid : _GEN_155; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_161 = btb_32_tag == io_i_addr[12:3] ? btb_32_target_address : _GEN_156; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_164 = btb_32_tag == io_i_addr[12:3] ? ~btb_32_bht[1] : _GEN_159; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_165 = btb_33_tag == io_i_addr[12:3] ? btb_33_valid : _GEN_160; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_166 = btb_33_tag == io_i_addr[12:3] ? btb_33_target_address : _GEN_161; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_169 = btb_33_tag == io_i_addr[12:3] ? ~btb_33_bht[1] : _GEN_164; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_170 = btb_34_tag == io_i_addr[12:3] ? btb_34_valid : _GEN_165; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_171 = btb_34_tag == io_i_addr[12:3] ? btb_34_target_address : _GEN_166; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_174 = btb_34_tag == io_i_addr[12:3] ? ~btb_34_bht[1] : _GEN_169; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_175 = btb_35_tag == io_i_addr[12:3] ? btb_35_valid : _GEN_170; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_176 = btb_35_tag == io_i_addr[12:3] ? btb_35_target_address : _GEN_171; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_179 = btb_35_tag == io_i_addr[12:3] ? ~btb_35_bht[1] : _GEN_174; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_180 = btb_36_tag == io_i_addr[12:3] ? btb_36_valid : _GEN_175; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_181 = btb_36_tag == io_i_addr[12:3] ? btb_36_target_address : _GEN_176; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_184 = btb_36_tag == io_i_addr[12:3] ? ~btb_36_bht[1] : _GEN_179; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_185 = btb_37_tag == io_i_addr[12:3] ? btb_37_valid : _GEN_180; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_186 = btb_37_tag == io_i_addr[12:3] ? btb_37_target_address : _GEN_181; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_189 = btb_37_tag == io_i_addr[12:3] ? ~btb_37_bht[1] : _GEN_184; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_190 = btb_38_tag == io_i_addr[12:3] ? btb_38_valid : _GEN_185; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_191 = btb_38_tag == io_i_addr[12:3] ? btb_38_target_address : _GEN_186; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_194 = btb_38_tag == io_i_addr[12:3] ? ~btb_38_bht[1] : _GEN_189; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_195 = btb_39_tag == io_i_addr[12:3] ? btb_39_valid : _GEN_190; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_196 = btb_39_tag == io_i_addr[12:3] ? btb_39_target_address : _GEN_191; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_199 = btb_39_tag == io_i_addr[12:3] ? ~btb_39_bht[1] : _GEN_194; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_200 = btb_40_tag == io_i_addr[12:3] ? btb_40_valid : _GEN_195; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_201 = btb_40_tag == io_i_addr[12:3] ? btb_40_target_address : _GEN_196; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_204 = btb_40_tag == io_i_addr[12:3] ? ~btb_40_bht[1] : _GEN_199; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_205 = btb_41_tag == io_i_addr[12:3] ? btb_41_valid : _GEN_200; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_206 = btb_41_tag == io_i_addr[12:3] ? btb_41_target_address : _GEN_201; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_209 = btb_41_tag == io_i_addr[12:3] ? ~btb_41_bht[1] : _GEN_204; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_210 = btb_42_tag == io_i_addr[12:3] ? btb_42_valid : _GEN_205; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_211 = btb_42_tag == io_i_addr[12:3] ? btb_42_target_address : _GEN_206; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_214 = btb_42_tag == io_i_addr[12:3] ? ~btb_42_bht[1] : _GEN_209; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_215 = btb_43_tag == io_i_addr[12:3] ? btb_43_valid : _GEN_210; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_216 = btb_43_tag == io_i_addr[12:3] ? btb_43_target_address : _GEN_211; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_219 = btb_43_tag == io_i_addr[12:3] ? ~btb_43_bht[1] : _GEN_214; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_220 = btb_44_tag == io_i_addr[12:3] ? btb_44_valid : _GEN_215; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_221 = btb_44_tag == io_i_addr[12:3] ? btb_44_target_address : _GEN_216; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_224 = btb_44_tag == io_i_addr[12:3] ? ~btb_44_bht[1] : _GEN_219; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_225 = btb_45_tag == io_i_addr[12:3] ? btb_45_valid : _GEN_220; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_226 = btb_45_tag == io_i_addr[12:3] ? btb_45_target_address : _GEN_221; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_229 = btb_45_tag == io_i_addr[12:3] ? ~btb_45_bht[1] : _GEN_224; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_230 = btb_46_tag == io_i_addr[12:3] ? btb_46_valid : _GEN_225; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_231 = btb_46_tag == io_i_addr[12:3] ? btb_46_target_address : _GEN_226; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_234 = btb_46_tag == io_i_addr[12:3] ? ~btb_46_bht[1] : _GEN_229; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_235 = btb_47_tag == io_i_addr[12:3] ? btb_47_valid : _GEN_230; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_236 = btb_47_tag == io_i_addr[12:3] ? btb_47_target_address : _GEN_231; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_239 = btb_47_tag == io_i_addr[12:3] ? ~btb_47_bht[1] : _GEN_234; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_240 = btb_48_tag == io_i_addr[12:3] ? btb_48_valid : _GEN_235; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_241 = btb_48_tag == io_i_addr[12:3] ? btb_48_target_address : _GEN_236; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_244 = btb_48_tag == io_i_addr[12:3] ? ~btb_48_bht[1] : _GEN_239; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_245 = btb_49_tag == io_i_addr[12:3] ? btb_49_valid : _GEN_240; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_246 = btb_49_tag == io_i_addr[12:3] ? btb_49_target_address : _GEN_241; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_249 = btb_49_tag == io_i_addr[12:3] ? ~btb_49_bht[1] : _GEN_244; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_250 = btb_50_tag == io_i_addr[12:3] ? btb_50_valid : _GEN_245; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_251 = btb_50_tag == io_i_addr[12:3] ? btb_50_target_address : _GEN_246; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_254 = btb_50_tag == io_i_addr[12:3] ? ~btb_50_bht[1] : _GEN_249; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_255 = btb_51_tag == io_i_addr[12:3] ? btb_51_valid : _GEN_250; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_256 = btb_51_tag == io_i_addr[12:3] ? btb_51_target_address : _GEN_251; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_259 = btb_51_tag == io_i_addr[12:3] ? ~btb_51_bht[1] : _GEN_254; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_260 = btb_52_tag == io_i_addr[12:3] ? btb_52_valid : _GEN_255; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_261 = btb_52_tag == io_i_addr[12:3] ? btb_52_target_address : _GEN_256; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_264 = btb_52_tag == io_i_addr[12:3] ? ~btb_52_bht[1] : _GEN_259; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_265 = btb_53_tag == io_i_addr[12:3] ? btb_53_valid : _GEN_260; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_266 = btb_53_tag == io_i_addr[12:3] ? btb_53_target_address : _GEN_261; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_269 = btb_53_tag == io_i_addr[12:3] ? ~btb_53_bht[1] : _GEN_264; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_270 = btb_54_tag == io_i_addr[12:3] ? btb_54_valid : _GEN_265; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_271 = btb_54_tag == io_i_addr[12:3] ? btb_54_target_address : _GEN_266; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_274 = btb_54_tag == io_i_addr[12:3] ? ~btb_54_bht[1] : _GEN_269; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_275 = btb_55_tag == io_i_addr[12:3] ? btb_55_valid : _GEN_270; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_276 = btb_55_tag == io_i_addr[12:3] ? btb_55_target_address : _GEN_271; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_279 = btb_55_tag == io_i_addr[12:3] ? ~btb_55_bht[1] : _GEN_274; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_280 = btb_56_tag == io_i_addr[12:3] ? btb_56_valid : _GEN_275; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_281 = btb_56_tag == io_i_addr[12:3] ? btb_56_target_address : _GEN_276; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_284 = btb_56_tag == io_i_addr[12:3] ? ~btb_56_bht[1] : _GEN_279; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_285 = btb_57_tag == io_i_addr[12:3] ? btb_57_valid : _GEN_280; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_286 = btb_57_tag == io_i_addr[12:3] ? btb_57_target_address : _GEN_281; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_289 = btb_57_tag == io_i_addr[12:3] ? ~btb_57_bht[1] : _GEN_284; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_290 = btb_58_tag == io_i_addr[12:3] ? btb_58_valid : _GEN_285; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_291 = btb_58_tag == io_i_addr[12:3] ? btb_58_target_address : _GEN_286; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_294 = btb_58_tag == io_i_addr[12:3] ? ~btb_58_bht[1] : _GEN_289; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_295 = btb_59_tag == io_i_addr[12:3] ? btb_59_valid : _GEN_290; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_296 = btb_59_tag == io_i_addr[12:3] ? btb_59_target_address : _GEN_291; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_299 = btb_59_tag == io_i_addr[12:3] ? ~btb_59_bht[1] : _GEN_294; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_300 = btb_60_tag == io_i_addr[12:3] ? btb_60_valid : _GEN_295; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_301 = btb_60_tag == io_i_addr[12:3] ? btb_60_target_address : _GEN_296; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_304 = btb_60_tag == io_i_addr[12:3] ? ~btb_60_bht[1] : _GEN_299; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_305 = btb_61_tag == io_i_addr[12:3] ? btb_61_valid : _GEN_300; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_306 = btb_61_tag == io_i_addr[12:3] ? btb_61_target_address : _GEN_301; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_309 = btb_61_tag == io_i_addr[12:3] ? ~btb_61_bht[1] : _GEN_304; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_310 = btb_62_tag == io_i_addr[12:3] ? btb_62_valid : _GEN_305; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_311 = btb_62_tag == io_i_addr[12:3] ? btb_62_target_address : _GEN_306; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_314 = btb_62_tag == io_i_addr[12:3] ? ~btb_62_bht[1] : _GEN_309; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_315 = btb_63_tag == io_i_addr[12:3] ? btb_63_valid : _GEN_310; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_316 = btb_63_tag == io_i_addr[12:3] ? btb_63_target_address : _GEN_311; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_319 = btb_63_tag == io_i_addr[12:3] ? ~btb_63_bht[1] : _GEN_314; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_320 = btb_64_tag == io_i_addr[12:3] ? btb_64_valid : _GEN_315; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_321 = btb_64_tag == io_i_addr[12:3] ? btb_64_target_address : _GEN_316; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_324 = btb_64_tag == io_i_addr[12:3] ? ~btb_64_bht[1] : _GEN_319; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_325 = btb_65_tag == io_i_addr[12:3] ? btb_65_valid : _GEN_320; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_326 = btb_65_tag == io_i_addr[12:3] ? btb_65_target_address : _GEN_321; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_329 = btb_65_tag == io_i_addr[12:3] ? ~btb_65_bht[1] : _GEN_324; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_330 = btb_66_tag == io_i_addr[12:3] ? btb_66_valid : _GEN_325; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_331 = btb_66_tag == io_i_addr[12:3] ? btb_66_target_address : _GEN_326; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_334 = btb_66_tag == io_i_addr[12:3] ? ~btb_66_bht[1] : _GEN_329; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_335 = btb_67_tag == io_i_addr[12:3] ? btb_67_valid : _GEN_330; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_336 = btb_67_tag == io_i_addr[12:3] ? btb_67_target_address : _GEN_331; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_339 = btb_67_tag == io_i_addr[12:3] ? ~btb_67_bht[1] : _GEN_334; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_340 = btb_68_tag == io_i_addr[12:3] ? btb_68_valid : _GEN_335; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_341 = btb_68_tag == io_i_addr[12:3] ? btb_68_target_address : _GEN_336; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_344 = btb_68_tag == io_i_addr[12:3] ? ~btb_68_bht[1] : _GEN_339; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_345 = btb_69_tag == io_i_addr[12:3] ? btb_69_valid : _GEN_340; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_346 = btb_69_tag == io_i_addr[12:3] ? btb_69_target_address : _GEN_341; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_349 = btb_69_tag == io_i_addr[12:3] ? ~btb_69_bht[1] : _GEN_344; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_350 = btb_70_tag == io_i_addr[12:3] ? btb_70_valid : _GEN_345; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_351 = btb_70_tag == io_i_addr[12:3] ? btb_70_target_address : _GEN_346; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_354 = btb_70_tag == io_i_addr[12:3] ? ~btb_70_bht[1] : _GEN_349; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_355 = btb_71_tag == io_i_addr[12:3] ? btb_71_valid : _GEN_350; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_356 = btb_71_tag == io_i_addr[12:3] ? btb_71_target_address : _GEN_351; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_359 = btb_71_tag == io_i_addr[12:3] ? ~btb_71_bht[1] : _GEN_354; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_360 = btb_72_tag == io_i_addr[12:3] ? btb_72_valid : _GEN_355; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_361 = btb_72_tag == io_i_addr[12:3] ? btb_72_target_address : _GEN_356; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_364 = btb_72_tag == io_i_addr[12:3] ? ~btb_72_bht[1] : _GEN_359; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_365 = btb_73_tag == io_i_addr[12:3] ? btb_73_valid : _GEN_360; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_366 = btb_73_tag == io_i_addr[12:3] ? btb_73_target_address : _GEN_361; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_369 = btb_73_tag == io_i_addr[12:3] ? ~btb_73_bht[1] : _GEN_364; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_370 = btb_74_tag == io_i_addr[12:3] ? btb_74_valid : _GEN_365; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_371 = btb_74_tag == io_i_addr[12:3] ? btb_74_target_address : _GEN_366; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_374 = btb_74_tag == io_i_addr[12:3] ? ~btb_74_bht[1] : _GEN_369; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_375 = btb_75_tag == io_i_addr[12:3] ? btb_75_valid : _GEN_370; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_376 = btb_75_tag == io_i_addr[12:3] ? btb_75_target_address : _GEN_371; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_379 = btb_75_tag == io_i_addr[12:3] ? ~btb_75_bht[1] : _GEN_374; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_380 = btb_76_tag == io_i_addr[12:3] ? btb_76_valid : _GEN_375; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_381 = btb_76_tag == io_i_addr[12:3] ? btb_76_target_address : _GEN_376; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_384 = btb_76_tag == io_i_addr[12:3] ? ~btb_76_bht[1] : _GEN_379; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_385 = btb_77_tag == io_i_addr[12:3] ? btb_77_valid : _GEN_380; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_386 = btb_77_tag == io_i_addr[12:3] ? btb_77_target_address : _GEN_381; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_389 = btb_77_tag == io_i_addr[12:3] ? ~btb_77_bht[1] : _GEN_384; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_390 = btb_78_tag == io_i_addr[12:3] ? btb_78_valid : _GEN_385; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_391 = btb_78_tag == io_i_addr[12:3] ? btb_78_target_address : _GEN_386; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_394 = btb_78_tag == io_i_addr[12:3] ? ~btb_78_bht[1] : _GEN_389; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_395 = btb_79_tag == io_i_addr[12:3] ? btb_79_valid : _GEN_390; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_396 = btb_79_tag == io_i_addr[12:3] ? btb_79_target_address : _GEN_391; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_399 = btb_79_tag == io_i_addr[12:3] ? ~btb_79_bht[1] : _GEN_394; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_400 = btb_80_tag == io_i_addr[12:3] ? btb_80_valid : _GEN_395; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_401 = btb_80_tag == io_i_addr[12:3] ? btb_80_target_address : _GEN_396; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_404 = btb_80_tag == io_i_addr[12:3] ? ~btb_80_bht[1] : _GEN_399; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_405 = btb_81_tag == io_i_addr[12:3] ? btb_81_valid : _GEN_400; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_406 = btb_81_tag == io_i_addr[12:3] ? btb_81_target_address : _GEN_401; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_409 = btb_81_tag == io_i_addr[12:3] ? ~btb_81_bht[1] : _GEN_404; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_410 = btb_82_tag == io_i_addr[12:3] ? btb_82_valid : _GEN_405; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_411 = btb_82_tag == io_i_addr[12:3] ? btb_82_target_address : _GEN_406; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_414 = btb_82_tag == io_i_addr[12:3] ? ~btb_82_bht[1] : _GEN_409; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_415 = btb_83_tag == io_i_addr[12:3] ? btb_83_valid : _GEN_410; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_416 = btb_83_tag == io_i_addr[12:3] ? btb_83_target_address : _GEN_411; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_419 = btb_83_tag == io_i_addr[12:3] ? ~btb_83_bht[1] : _GEN_414; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_420 = btb_84_tag == io_i_addr[12:3] ? btb_84_valid : _GEN_415; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_421 = btb_84_tag == io_i_addr[12:3] ? btb_84_target_address : _GEN_416; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_424 = btb_84_tag == io_i_addr[12:3] ? ~btb_84_bht[1] : _GEN_419; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_425 = btb_85_tag == io_i_addr[12:3] ? btb_85_valid : _GEN_420; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_426 = btb_85_tag == io_i_addr[12:3] ? btb_85_target_address : _GEN_421; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_429 = btb_85_tag == io_i_addr[12:3] ? ~btb_85_bht[1] : _GEN_424; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_430 = btb_86_tag == io_i_addr[12:3] ? btb_86_valid : _GEN_425; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_431 = btb_86_tag == io_i_addr[12:3] ? btb_86_target_address : _GEN_426; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_434 = btb_86_tag == io_i_addr[12:3] ? ~btb_86_bht[1] : _GEN_429; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_435 = btb_87_tag == io_i_addr[12:3] ? btb_87_valid : _GEN_430; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_436 = btb_87_tag == io_i_addr[12:3] ? btb_87_target_address : _GEN_431; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_439 = btb_87_tag == io_i_addr[12:3] ? ~btb_87_bht[1] : _GEN_434; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_440 = btb_88_tag == io_i_addr[12:3] ? btb_88_valid : _GEN_435; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_441 = btb_88_tag == io_i_addr[12:3] ? btb_88_target_address : _GEN_436; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_444 = btb_88_tag == io_i_addr[12:3] ? ~btb_88_bht[1] : _GEN_439; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_445 = btb_89_tag == io_i_addr[12:3] ? btb_89_valid : _GEN_440; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_446 = btb_89_tag == io_i_addr[12:3] ? btb_89_target_address : _GEN_441; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_449 = btb_89_tag == io_i_addr[12:3] ? ~btb_89_bht[1] : _GEN_444; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_450 = btb_90_tag == io_i_addr[12:3] ? btb_90_valid : _GEN_445; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_451 = btb_90_tag == io_i_addr[12:3] ? btb_90_target_address : _GEN_446; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_454 = btb_90_tag == io_i_addr[12:3] ? ~btb_90_bht[1] : _GEN_449; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_455 = btb_91_tag == io_i_addr[12:3] ? btb_91_valid : _GEN_450; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_456 = btb_91_tag == io_i_addr[12:3] ? btb_91_target_address : _GEN_451; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_459 = btb_91_tag == io_i_addr[12:3] ? ~btb_91_bht[1] : _GEN_454; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_460 = btb_92_tag == io_i_addr[12:3] ? btb_92_valid : _GEN_455; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_461 = btb_92_tag == io_i_addr[12:3] ? btb_92_target_address : _GEN_456; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_464 = btb_92_tag == io_i_addr[12:3] ? ~btb_92_bht[1] : _GEN_459; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_465 = btb_93_tag == io_i_addr[12:3] ? btb_93_valid : _GEN_460; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_466 = btb_93_tag == io_i_addr[12:3] ? btb_93_target_address : _GEN_461; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_469 = btb_93_tag == io_i_addr[12:3] ? ~btb_93_bht[1] : _GEN_464; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_470 = btb_94_tag == io_i_addr[12:3] ? btb_94_valid : _GEN_465; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_471 = btb_94_tag == io_i_addr[12:3] ? btb_94_target_address : _GEN_466; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_474 = btb_94_tag == io_i_addr[12:3] ? ~btb_94_bht[1] : _GEN_469; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_475 = btb_95_tag == io_i_addr[12:3] ? btb_95_valid : _GEN_470; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_476 = btb_95_tag == io_i_addr[12:3] ? btb_95_target_address : _GEN_471; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_479 = btb_95_tag == io_i_addr[12:3] ? ~btb_95_bht[1] : _GEN_474; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_480 = btb_96_tag == io_i_addr[12:3] ? btb_96_valid : _GEN_475; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_481 = btb_96_tag == io_i_addr[12:3] ? btb_96_target_address : _GEN_476; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_484 = btb_96_tag == io_i_addr[12:3] ? ~btb_96_bht[1] : _GEN_479; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_485 = btb_97_tag == io_i_addr[12:3] ? btb_97_valid : _GEN_480; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_486 = btb_97_tag == io_i_addr[12:3] ? btb_97_target_address : _GEN_481; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_489 = btb_97_tag == io_i_addr[12:3] ? ~btb_97_bht[1] : _GEN_484; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_490 = btb_98_tag == io_i_addr[12:3] ? btb_98_valid : _GEN_485; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_491 = btb_98_tag == io_i_addr[12:3] ? btb_98_target_address : _GEN_486; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_494 = btb_98_tag == io_i_addr[12:3] ? ~btb_98_bht[1] : _GEN_489; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_495 = btb_99_tag == io_i_addr[12:3] ? btb_99_valid : _GEN_490; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_496 = btb_99_tag == io_i_addr[12:3] ? btb_99_target_address : _GEN_491; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_499 = btb_99_tag == io_i_addr[12:3] ? ~btb_99_bht[1] : _GEN_494; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_500 = btb_100_tag == io_i_addr[12:3] ? btb_100_valid : _GEN_495; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_501 = btb_100_tag == io_i_addr[12:3] ? btb_100_target_address : _GEN_496; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_504 = btb_100_tag == io_i_addr[12:3] ? ~btb_100_bht[1] : _GEN_499; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_505 = btb_101_tag == io_i_addr[12:3] ? btb_101_valid : _GEN_500; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_506 = btb_101_tag == io_i_addr[12:3] ? btb_101_target_address : _GEN_501; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_509 = btb_101_tag == io_i_addr[12:3] ? ~btb_101_bht[1] : _GEN_504; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_510 = btb_102_tag == io_i_addr[12:3] ? btb_102_valid : _GEN_505; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_511 = btb_102_tag == io_i_addr[12:3] ? btb_102_target_address : _GEN_506; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_514 = btb_102_tag == io_i_addr[12:3] ? ~btb_102_bht[1] : _GEN_509; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_515 = btb_103_tag == io_i_addr[12:3] ? btb_103_valid : _GEN_510; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_516 = btb_103_tag == io_i_addr[12:3] ? btb_103_target_address : _GEN_511; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_519 = btb_103_tag == io_i_addr[12:3] ? ~btb_103_bht[1] : _GEN_514; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_520 = btb_104_tag == io_i_addr[12:3] ? btb_104_valid : _GEN_515; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_521 = btb_104_tag == io_i_addr[12:3] ? btb_104_target_address : _GEN_516; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_524 = btb_104_tag == io_i_addr[12:3] ? ~btb_104_bht[1] : _GEN_519; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_525 = btb_105_tag == io_i_addr[12:3] ? btb_105_valid : _GEN_520; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_526 = btb_105_tag == io_i_addr[12:3] ? btb_105_target_address : _GEN_521; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_529 = btb_105_tag == io_i_addr[12:3] ? ~btb_105_bht[1] : _GEN_524; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_530 = btb_106_tag == io_i_addr[12:3] ? btb_106_valid : _GEN_525; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_531 = btb_106_tag == io_i_addr[12:3] ? btb_106_target_address : _GEN_526; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_534 = btb_106_tag == io_i_addr[12:3] ? ~btb_106_bht[1] : _GEN_529; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_535 = btb_107_tag == io_i_addr[12:3] ? btb_107_valid : _GEN_530; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_536 = btb_107_tag == io_i_addr[12:3] ? btb_107_target_address : _GEN_531; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_539 = btb_107_tag == io_i_addr[12:3] ? ~btb_107_bht[1] : _GEN_534; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_540 = btb_108_tag == io_i_addr[12:3] ? btb_108_valid : _GEN_535; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_541 = btb_108_tag == io_i_addr[12:3] ? btb_108_target_address : _GEN_536; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_544 = btb_108_tag == io_i_addr[12:3] ? ~btb_108_bht[1] : _GEN_539; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_545 = btb_109_tag == io_i_addr[12:3] ? btb_109_valid : _GEN_540; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_546 = btb_109_tag == io_i_addr[12:3] ? btb_109_target_address : _GEN_541; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_549 = btb_109_tag == io_i_addr[12:3] ? ~btb_109_bht[1] : _GEN_544; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_550 = btb_110_tag == io_i_addr[12:3] ? btb_110_valid : _GEN_545; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_551 = btb_110_tag == io_i_addr[12:3] ? btb_110_target_address : _GEN_546; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_554 = btb_110_tag == io_i_addr[12:3] ? ~btb_110_bht[1] : _GEN_549; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_555 = btb_111_tag == io_i_addr[12:3] ? btb_111_valid : _GEN_550; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_556 = btb_111_tag == io_i_addr[12:3] ? btb_111_target_address : _GEN_551; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_559 = btb_111_tag == io_i_addr[12:3] ? ~btb_111_bht[1] : _GEN_554; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_560 = btb_112_tag == io_i_addr[12:3] ? btb_112_valid : _GEN_555; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_561 = btb_112_tag == io_i_addr[12:3] ? btb_112_target_address : _GEN_556; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_564 = btb_112_tag == io_i_addr[12:3] ? ~btb_112_bht[1] : _GEN_559; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_565 = btb_113_tag == io_i_addr[12:3] ? btb_113_valid : _GEN_560; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_566 = btb_113_tag == io_i_addr[12:3] ? btb_113_target_address : _GEN_561; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_569 = btb_113_tag == io_i_addr[12:3] ? ~btb_113_bht[1] : _GEN_564; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_570 = btb_114_tag == io_i_addr[12:3] ? btb_114_valid : _GEN_565; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_571 = btb_114_tag == io_i_addr[12:3] ? btb_114_target_address : _GEN_566; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_574 = btb_114_tag == io_i_addr[12:3] ? ~btb_114_bht[1] : _GEN_569; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_575 = btb_115_tag == io_i_addr[12:3] ? btb_115_valid : _GEN_570; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_576 = btb_115_tag == io_i_addr[12:3] ? btb_115_target_address : _GEN_571; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_579 = btb_115_tag == io_i_addr[12:3] ? ~btb_115_bht[1] : _GEN_574; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_580 = btb_116_tag == io_i_addr[12:3] ? btb_116_valid : _GEN_575; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_581 = btb_116_tag == io_i_addr[12:3] ? btb_116_target_address : _GEN_576; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_584 = btb_116_tag == io_i_addr[12:3] ? ~btb_116_bht[1] : _GEN_579; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_585 = btb_117_tag == io_i_addr[12:3] ? btb_117_valid : _GEN_580; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_586 = btb_117_tag == io_i_addr[12:3] ? btb_117_target_address : _GEN_581; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_589 = btb_117_tag == io_i_addr[12:3] ? ~btb_117_bht[1] : _GEN_584; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_590 = btb_118_tag == io_i_addr[12:3] ? btb_118_valid : _GEN_585; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_591 = btb_118_tag == io_i_addr[12:3] ? btb_118_target_address : _GEN_586; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_594 = btb_118_tag == io_i_addr[12:3] ? ~btb_118_bht[1] : _GEN_589; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_595 = btb_119_tag == io_i_addr[12:3] ? btb_119_valid : _GEN_590; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_596 = btb_119_tag == io_i_addr[12:3] ? btb_119_target_address : _GEN_591; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_599 = btb_119_tag == io_i_addr[12:3] ? ~btb_119_bht[1] : _GEN_594; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_600 = btb_120_tag == io_i_addr[12:3] ? btb_120_valid : _GEN_595; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_601 = btb_120_tag == io_i_addr[12:3] ? btb_120_target_address : _GEN_596; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_604 = btb_120_tag == io_i_addr[12:3] ? ~btb_120_bht[1] : _GEN_599; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_605 = btb_121_tag == io_i_addr[12:3] ? btb_121_valid : _GEN_600; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_606 = btb_121_tag == io_i_addr[12:3] ? btb_121_target_address : _GEN_601; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_609 = btb_121_tag == io_i_addr[12:3] ? ~btb_121_bht[1] : _GEN_604; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_610 = btb_122_tag == io_i_addr[12:3] ? btb_122_valid : _GEN_605; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_611 = btb_122_tag == io_i_addr[12:3] ? btb_122_target_address : _GEN_606; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_614 = btb_122_tag == io_i_addr[12:3] ? ~btb_122_bht[1] : _GEN_609; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_615 = btb_123_tag == io_i_addr[12:3] ? btb_123_valid : _GEN_610; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_616 = btb_123_tag == io_i_addr[12:3] ? btb_123_target_address : _GEN_611; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_619 = btb_123_tag == io_i_addr[12:3] ? ~btb_123_bht[1] : _GEN_614; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_620 = btb_124_tag == io_i_addr[12:3] ? btb_124_valid : _GEN_615; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_621 = btb_124_tag == io_i_addr[12:3] ? btb_124_target_address : _GEN_616; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_624 = btb_124_tag == io_i_addr[12:3] ? ~btb_124_bht[1] : _GEN_619; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_625 = btb_125_tag == io_i_addr[12:3] ? btb_125_valid : _GEN_620; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_626 = btb_125_tag == io_i_addr[12:3] ? btb_125_target_address : _GEN_621; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_629 = btb_125_tag == io_i_addr[12:3] ? ~btb_125_bht[1] : _GEN_624; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_630 = btb_126_tag == io_i_addr[12:3] ? btb_126_valid : _GEN_625; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_631 = btb_126_tag == io_i_addr[12:3] ? btb_126_target_address : _GEN_626; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_634 = btb_126_tag == io_i_addr[12:3] ? ~btb_126_bht[1] : _GEN_629; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_635 = btb_127_tag == io_i_addr[12:3] ? btb_127_valid : _GEN_630; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_636 = btb_127_tag == io_i_addr[12:3] ? btb_127_target_address : _GEN_631; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_639 = btb_127_tag == io_i_addr[12:3] ? ~btb_127_bht[1] : _GEN_634; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_640 = btb_128_tag == io_i_addr[12:3] ? btb_128_valid : _GEN_635; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_641 = btb_128_tag == io_i_addr[12:3] ? btb_128_target_address : _GEN_636; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_644 = btb_128_tag == io_i_addr[12:3] ? ~btb_128_bht[1] : _GEN_639; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_645 = btb_129_tag == io_i_addr[12:3] ? btb_129_valid : _GEN_640; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_646 = btb_129_tag == io_i_addr[12:3] ? btb_129_target_address : _GEN_641; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_649 = btb_129_tag == io_i_addr[12:3] ? ~btb_129_bht[1] : _GEN_644; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_650 = btb_130_tag == io_i_addr[12:3] ? btb_130_valid : _GEN_645; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_651 = btb_130_tag == io_i_addr[12:3] ? btb_130_target_address : _GEN_646; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_654 = btb_130_tag == io_i_addr[12:3] ? ~btb_130_bht[1] : _GEN_649; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_655 = btb_131_tag == io_i_addr[12:3] ? btb_131_valid : _GEN_650; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_656 = btb_131_tag == io_i_addr[12:3] ? btb_131_target_address : _GEN_651; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_659 = btb_131_tag == io_i_addr[12:3] ? ~btb_131_bht[1] : _GEN_654; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_660 = btb_132_tag == io_i_addr[12:3] ? btb_132_valid : _GEN_655; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_661 = btb_132_tag == io_i_addr[12:3] ? btb_132_target_address : _GEN_656; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_664 = btb_132_tag == io_i_addr[12:3] ? ~btb_132_bht[1] : _GEN_659; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_665 = btb_133_tag == io_i_addr[12:3] ? btb_133_valid : _GEN_660; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_666 = btb_133_tag == io_i_addr[12:3] ? btb_133_target_address : _GEN_661; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_669 = btb_133_tag == io_i_addr[12:3] ? ~btb_133_bht[1] : _GEN_664; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_670 = btb_134_tag == io_i_addr[12:3] ? btb_134_valid : _GEN_665; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_671 = btb_134_tag == io_i_addr[12:3] ? btb_134_target_address : _GEN_666; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_674 = btb_134_tag == io_i_addr[12:3] ? ~btb_134_bht[1] : _GEN_669; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_675 = btb_135_tag == io_i_addr[12:3] ? btb_135_valid : _GEN_670; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_676 = btb_135_tag == io_i_addr[12:3] ? btb_135_target_address : _GEN_671; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_679 = btb_135_tag == io_i_addr[12:3] ? ~btb_135_bht[1] : _GEN_674; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_680 = btb_136_tag == io_i_addr[12:3] ? btb_136_valid : _GEN_675; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_681 = btb_136_tag == io_i_addr[12:3] ? btb_136_target_address : _GEN_676; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_684 = btb_136_tag == io_i_addr[12:3] ? ~btb_136_bht[1] : _GEN_679; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_685 = btb_137_tag == io_i_addr[12:3] ? btb_137_valid : _GEN_680; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_686 = btb_137_tag == io_i_addr[12:3] ? btb_137_target_address : _GEN_681; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_689 = btb_137_tag == io_i_addr[12:3] ? ~btb_137_bht[1] : _GEN_684; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_690 = btb_138_tag == io_i_addr[12:3] ? btb_138_valid : _GEN_685; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_691 = btb_138_tag == io_i_addr[12:3] ? btb_138_target_address : _GEN_686; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_694 = btb_138_tag == io_i_addr[12:3] ? ~btb_138_bht[1] : _GEN_689; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_695 = btb_139_tag == io_i_addr[12:3] ? btb_139_valid : _GEN_690; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_696 = btb_139_tag == io_i_addr[12:3] ? btb_139_target_address : _GEN_691; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_699 = btb_139_tag == io_i_addr[12:3] ? ~btb_139_bht[1] : _GEN_694; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_700 = btb_140_tag == io_i_addr[12:3] ? btb_140_valid : _GEN_695; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_701 = btb_140_tag == io_i_addr[12:3] ? btb_140_target_address : _GEN_696; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_704 = btb_140_tag == io_i_addr[12:3] ? ~btb_140_bht[1] : _GEN_699; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_705 = btb_141_tag == io_i_addr[12:3] ? btb_141_valid : _GEN_700; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_706 = btb_141_tag == io_i_addr[12:3] ? btb_141_target_address : _GEN_701; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_709 = btb_141_tag == io_i_addr[12:3] ? ~btb_141_bht[1] : _GEN_704; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_710 = btb_142_tag == io_i_addr[12:3] ? btb_142_valid : _GEN_705; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_711 = btb_142_tag == io_i_addr[12:3] ? btb_142_target_address : _GEN_706; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_714 = btb_142_tag == io_i_addr[12:3] ? ~btb_142_bht[1] : _GEN_709; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_715 = btb_143_tag == io_i_addr[12:3] ? btb_143_valid : _GEN_710; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_716 = btb_143_tag == io_i_addr[12:3] ? btb_143_target_address : _GEN_711; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_719 = btb_143_tag == io_i_addr[12:3] ? ~btb_143_bht[1] : _GEN_714; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_720 = btb_144_tag == io_i_addr[12:3] ? btb_144_valid : _GEN_715; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_721 = btb_144_tag == io_i_addr[12:3] ? btb_144_target_address : _GEN_716; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_724 = btb_144_tag == io_i_addr[12:3] ? ~btb_144_bht[1] : _GEN_719; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_725 = btb_145_tag == io_i_addr[12:3] ? btb_145_valid : _GEN_720; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_726 = btb_145_tag == io_i_addr[12:3] ? btb_145_target_address : _GEN_721; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_729 = btb_145_tag == io_i_addr[12:3] ? ~btb_145_bht[1] : _GEN_724; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_730 = btb_146_tag == io_i_addr[12:3] ? btb_146_valid : _GEN_725; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_731 = btb_146_tag == io_i_addr[12:3] ? btb_146_target_address : _GEN_726; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_734 = btb_146_tag == io_i_addr[12:3] ? ~btb_146_bht[1] : _GEN_729; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_735 = btb_147_tag == io_i_addr[12:3] ? btb_147_valid : _GEN_730; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_736 = btb_147_tag == io_i_addr[12:3] ? btb_147_target_address : _GEN_731; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_739 = btb_147_tag == io_i_addr[12:3] ? ~btb_147_bht[1] : _GEN_734; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_740 = btb_148_tag == io_i_addr[12:3] ? btb_148_valid : _GEN_735; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_741 = btb_148_tag == io_i_addr[12:3] ? btb_148_target_address : _GEN_736; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_744 = btb_148_tag == io_i_addr[12:3] ? ~btb_148_bht[1] : _GEN_739; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_745 = btb_149_tag == io_i_addr[12:3] ? btb_149_valid : _GEN_740; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_746 = btb_149_tag == io_i_addr[12:3] ? btb_149_target_address : _GEN_741; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_749 = btb_149_tag == io_i_addr[12:3] ? ~btb_149_bht[1] : _GEN_744; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_750 = btb_150_tag == io_i_addr[12:3] ? btb_150_valid : _GEN_745; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_751 = btb_150_tag == io_i_addr[12:3] ? btb_150_target_address : _GEN_746; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_754 = btb_150_tag == io_i_addr[12:3] ? ~btb_150_bht[1] : _GEN_749; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_755 = btb_151_tag == io_i_addr[12:3] ? btb_151_valid : _GEN_750; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_756 = btb_151_tag == io_i_addr[12:3] ? btb_151_target_address : _GEN_751; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_759 = btb_151_tag == io_i_addr[12:3] ? ~btb_151_bht[1] : _GEN_754; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_760 = btb_152_tag == io_i_addr[12:3] ? btb_152_valid : _GEN_755; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_761 = btb_152_tag == io_i_addr[12:3] ? btb_152_target_address : _GEN_756; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_764 = btb_152_tag == io_i_addr[12:3] ? ~btb_152_bht[1] : _GEN_759; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_765 = btb_153_tag == io_i_addr[12:3] ? btb_153_valid : _GEN_760; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_766 = btb_153_tag == io_i_addr[12:3] ? btb_153_target_address : _GEN_761; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_769 = btb_153_tag == io_i_addr[12:3] ? ~btb_153_bht[1] : _GEN_764; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_770 = btb_154_tag == io_i_addr[12:3] ? btb_154_valid : _GEN_765; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_771 = btb_154_tag == io_i_addr[12:3] ? btb_154_target_address : _GEN_766; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_774 = btb_154_tag == io_i_addr[12:3] ? ~btb_154_bht[1] : _GEN_769; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_775 = btb_155_tag == io_i_addr[12:3] ? btb_155_valid : _GEN_770; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_776 = btb_155_tag == io_i_addr[12:3] ? btb_155_target_address : _GEN_771; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_779 = btb_155_tag == io_i_addr[12:3] ? ~btb_155_bht[1] : _GEN_774; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_780 = btb_156_tag == io_i_addr[12:3] ? btb_156_valid : _GEN_775; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_781 = btb_156_tag == io_i_addr[12:3] ? btb_156_target_address : _GEN_776; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_784 = btb_156_tag == io_i_addr[12:3] ? ~btb_156_bht[1] : _GEN_779; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_785 = btb_157_tag == io_i_addr[12:3] ? btb_157_valid : _GEN_780; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_786 = btb_157_tag == io_i_addr[12:3] ? btb_157_target_address : _GEN_781; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_789 = btb_157_tag == io_i_addr[12:3] ? ~btb_157_bht[1] : _GEN_784; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_790 = btb_158_tag == io_i_addr[12:3] ? btb_158_valid : _GEN_785; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_791 = btb_158_tag == io_i_addr[12:3] ? btb_158_target_address : _GEN_786; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_794 = btb_158_tag == io_i_addr[12:3] ? ~btb_158_bht[1] : _GEN_789; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_795 = btb_159_tag == io_i_addr[12:3] ? btb_159_valid : _GEN_790; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_796 = btb_159_tag == io_i_addr[12:3] ? btb_159_target_address : _GEN_791; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_799 = btb_159_tag == io_i_addr[12:3] ? ~btb_159_bht[1] : _GEN_794; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_800 = btb_160_tag == io_i_addr[12:3] ? btb_160_valid : _GEN_795; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_801 = btb_160_tag == io_i_addr[12:3] ? btb_160_target_address : _GEN_796; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_804 = btb_160_tag == io_i_addr[12:3] ? ~btb_160_bht[1] : _GEN_799; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_805 = btb_161_tag == io_i_addr[12:3] ? btb_161_valid : _GEN_800; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_806 = btb_161_tag == io_i_addr[12:3] ? btb_161_target_address : _GEN_801; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_809 = btb_161_tag == io_i_addr[12:3] ? ~btb_161_bht[1] : _GEN_804; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_810 = btb_162_tag == io_i_addr[12:3] ? btb_162_valid : _GEN_805; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_811 = btb_162_tag == io_i_addr[12:3] ? btb_162_target_address : _GEN_806; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_814 = btb_162_tag == io_i_addr[12:3] ? ~btb_162_bht[1] : _GEN_809; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_815 = btb_163_tag == io_i_addr[12:3] ? btb_163_valid : _GEN_810; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_816 = btb_163_tag == io_i_addr[12:3] ? btb_163_target_address : _GEN_811; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_819 = btb_163_tag == io_i_addr[12:3] ? ~btb_163_bht[1] : _GEN_814; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_820 = btb_164_tag == io_i_addr[12:3] ? btb_164_valid : _GEN_815; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_821 = btb_164_tag == io_i_addr[12:3] ? btb_164_target_address : _GEN_816; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_824 = btb_164_tag == io_i_addr[12:3] ? ~btb_164_bht[1] : _GEN_819; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_825 = btb_165_tag == io_i_addr[12:3] ? btb_165_valid : _GEN_820; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_826 = btb_165_tag == io_i_addr[12:3] ? btb_165_target_address : _GEN_821; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_829 = btb_165_tag == io_i_addr[12:3] ? ~btb_165_bht[1] : _GEN_824; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_830 = btb_166_tag == io_i_addr[12:3] ? btb_166_valid : _GEN_825; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_831 = btb_166_tag == io_i_addr[12:3] ? btb_166_target_address : _GEN_826; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_834 = btb_166_tag == io_i_addr[12:3] ? ~btb_166_bht[1] : _GEN_829; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_835 = btb_167_tag == io_i_addr[12:3] ? btb_167_valid : _GEN_830; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_836 = btb_167_tag == io_i_addr[12:3] ? btb_167_target_address : _GEN_831; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_839 = btb_167_tag == io_i_addr[12:3] ? ~btb_167_bht[1] : _GEN_834; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_840 = btb_168_tag == io_i_addr[12:3] ? btb_168_valid : _GEN_835; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_841 = btb_168_tag == io_i_addr[12:3] ? btb_168_target_address : _GEN_836; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_844 = btb_168_tag == io_i_addr[12:3] ? ~btb_168_bht[1] : _GEN_839; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_845 = btb_169_tag == io_i_addr[12:3] ? btb_169_valid : _GEN_840; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_846 = btb_169_tag == io_i_addr[12:3] ? btb_169_target_address : _GEN_841; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_849 = btb_169_tag == io_i_addr[12:3] ? ~btb_169_bht[1] : _GEN_844; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_850 = btb_170_tag == io_i_addr[12:3] ? btb_170_valid : _GEN_845; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_851 = btb_170_tag == io_i_addr[12:3] ? btb_170_target_address : _GEN_846; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_854 = btb_170_tag == io_i_addr[12:3] ? ~btb_170_bht[1] : _GEN_849; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_855 = btb_171_tag == io_i_addr[12:3] ? btb_171_valid : _GEN_850; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_856 = btb_171_tag == io_i_addr[12:3] ? btb_171_target_address : _GEN_851; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_859 = btb_171_tag == io_i_addr[12:3] ? ~btb_171_bht[1] : _GEN_854; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_860 = btb_172_tag == io_i_addr[12:3] ? btb_172_valid : _GEN_855; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_861 = btb_172_tag == io_i_addr[12:3] ? btb_172_target_address : _GEN_856; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_864 = btb_172_tag == io_i_addr[12:3] ? ~btb_172_bht[1] : _GEN_859; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_865 = btb_173_tag == io_i_addr[12:3] ? btb_173_valid : _GEN_860; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_866 = btb_173_tag == io_i_addr[12:3] ? btb_173_target_address : _GEN_861; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_869 = btb_173_tag == io_i_addr[12:3] ? ~btb_173_bht[1] : _GEN_864; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_870 = btb_174_tag == io_i_addr[12:3] ? btb_174_valid : _GEN_865; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_871 = btb_174_tag == io_i_addr[12:3] ? btb_174_target_address : _GEN_866; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_874 = btb_174_tag == io_i_addr[12:3] ? ~btb_174_bht[1] : _GEN_869; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_875 = btb_175_tag == io_i_addr[12:3] ? btb_175_valid : _GEN_870; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_876 = btb_175_tag == io_i_addr[12:3] ? btb_175_target_address : _GEN_871; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_879 = btb_175_tag == io_i_addr[12:3] ? ~btb_175_bht[1] : _GEN_874; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_880 = btb_176_tag == io_i_addr[12:3] ? btb_176_valid : _GEN_875; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_881 = btb_176_tag == io_i_addr[12:3] ? btb_176_target_address : _GEN_876; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_884 = btb_176_tag == io_i_addr[12:3] ? ~btb_176_bht[1] : _GEN_879; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_885 = btb_177_tag == io_i_addr[12:3] ? btb_177_valid : _GEN_880; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_886 = btb_177_tag == io_i_addr[12:3] ? btb_177_target_address : _GEN_881; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_889 = btb_177_tag == io_i_addr[12:3] ? ~btb_177_bht[1] : _GEN_884; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_890 = btb_178_tag == io_i_addr[12:3] ? btb_178_valid : _GEN_885; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_891 = btb_178_tag == io_i_addr[12:3] ? btb_178_target_address : _GEN_886; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_894 = btb_178_tag == io_i_addr[12:3] ? ~btb_178_bht[1] : _GEN_889; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_895 = btb_179_tag == io_i_addr[12:3] ? btb_179_valid : _GEN_890; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_896 = btb_179_tag == io_i_addr[12:3] ? btb_179_target_address : _GEN_891; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_899 = btb_179_tag == io_i_addr[12:3] ? ~btb_179_bht[1] : _GEN_894; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_900 = btb_180_tag == io_i_addr[12:3] ? btb_180_valid : _GEN_895; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_901 = btb_180_tag == io_i_addr[12:3] ? btb_180_target_address : _GEN_896; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_904 = btb_180_tag == io_i_addr[12:3] ? ~btb_180_bht[1] : _GEN_899; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_905 = btb_181_tag == io_i_addr[12:3] ? btb_181_valid : _GEN_900; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_906 = btb_181_tag == io_i_addr[12:3] ? btb_181_target_address : _GEN_901; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_909 = btb_181_tag == io_i_addr[12:3] ? ~btb_181_bht[1] : _GEN_904; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_910 = btb_182_tag == io_i_addr[12:3] ? btb_182_valid : _GEN_905; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_911 = btb_182_tag == io_i_addr[12:3] ? btb_182_target_address : _GEN_906; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_914 = btb_182_tag == io_i_addr[12:3] ? ~btb_182_bht[1] : _GEN_909; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_915 = btb_183_tag == io_i_addr[12:3] ? btb_183_valid : _GEN_910; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_916 = btb_183_tag == io_i_addr[12:3] ? btb_183_target_address : _GEN_911; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_919 = btb_183_tag == io_i_addr[12:3] ? ~btb_183_bht[1] : _GEN_914; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_920 = btb_184_tag == io_i_addr[12:3] ? btb_184_valid : _GEN_915; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_921 = btb_184_tag == io_i_addr[12:3] ? btb_184_target_address : _GEN_916; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_924 = btb_184_tag == io_i_addr[12:3] ? ~btb_184_bht[1] : _GEN_919; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_925 = btb_185_tag == io_i_addr[12:3] ? btb_185_valid : _GEN_920; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_926 = btb_185_tag == io_i_addr[12:3] ? btb_185_target_address : _GEN_921; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_929 = btb_185_tag == io_i_addr[12:3] ? ~btb_185_bht[1] : _GEN_924; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_930 = btb_186_tag == io_i_addr[12:3] ? btb_186_valid : _GEN_925; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_931 = btb_186_tag == io_i_addr[12:3] ? btb_186_target_address : _GEN_926; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_934 = btb_186_tag == io_i_addr[12:3] ? ~btb_186_bht[1] : _GEN_929; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_935 = btb_187_tag == io_i_addr[12:3] ? btb_187_valid : _GEN_930; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_936 = btb_187_tag == io_i_addr[12:3] ? btb_187_target_address : _GEN_931; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_939 = btb_187_tag == io_i_addr[12:3] ? ~btb_187_bht[1] : _GEN_934; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_940 = btb_188_tag == io_i_addr[12:3] ? btb_188_valid : _GEN_935; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_941 = btb_188_tag == io_i_addr[12:3] ? btb_188_target_address : _GEN_936; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_944 = btb_188_tag == io_i_addr[12:3] ? ~btb_188_bht[1] : _GEN_939; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_945 = btb_189_tag == io_i_addr[12:3] ? btb_189_valid : _GEN_940; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_946 = btb_189_tag == io_i_addr[12:3] ? btb_189_target_address : _GEN_941; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_949 = btb_189_tag == io_i_addr[12:3] ? ~btb_189_bht[1] : _GEN_944; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_950 = btb_190_tag == io_i_addr[12:3] ? btb_190_valid : _GEN_945; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_951 = btb_190_tag == io_i_addr[12:3] ? btb_190_target_address : _GEN_946; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_954 = btb_190_tag == io_i_addr[12:3] ? ~btb_190_bht[1] : _GEN_949; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_955 = btb_191_tag == io_i_addr[12:3] ? btb_191_valid : _GEN_950; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_956 = btb_191_tag == io_i_addr[12:3] ? btb_191_target_address : _GEN_951; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_959 = btb_191_tag == io_i_addr[12:3] ? ~btb_191_bht[1] : _GEN_954; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_960 = btb_192_tag == io_i_addr[12:3] ? btb_192_valid : _GEN_955; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_961 = btb_192_tag == io_i_addr[12:3] ? btb_192_target_address : _GEN_956; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_964 = btb_192_tag == io_i_addr[12:3] ? ~btb_192_bht[1] : _GEN_959; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_965 = btb_193_tag == io_i_addr[12:3] ? btb_193_valid : _GEN_960; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_966 = btb_193_tag == io_i_addr[12:3] ? btb_193_target_address : _GEN_961; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_969 = btb_193_tag == io_i_addr[12:3] ? ~btb_193_bht[1] : _GEN_964; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_970 = btb_194_tag == io_i_addr[12:3] ? btb_194_valid : _GEN_965; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_971 = btb_194_tag == io_i_addr[12:3] ? btb_194_target_address : _GEN_966; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_974 = btb_194_tag == io_i_addr[12:3] ? ~btb_194_bht[1] : _GEN_969; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_975 = btb_195_tag == io_i_addr[12:3] ? btb_195_valid : _GEN_970; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_976 = btb_195_tag == io_i_addr[12:3] ? btb_195_target_address : _GEN_971; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_979 = btb_195_tag == io_i_addr[12:3] ? ~btb_195_bht[1] : _GEN_974; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_980 = btb_196_tag == io_i_addr[12:3] ? btb_196_valid : _GEN_975; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_981 = btb_196_tag == io_i_addr[12:3] ? btb_196_target_address : _GEN_976; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_984 = btb_196_tag == io_i_addr[12:3] ? ~btb_196_bht[1] : _GEN_979; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_985 = btb_197_tag == io_i_addr[12:3] ? btb_197_valid : _GEN_980; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_986 = btb_197_tag == io_i_addr[12:3] ? btb_197_target_address : _GEN_981; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_989 = btb_197_tag == io_i_addr[12:3] ? ~btb_197_bht[1] : _GEN_984; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_990 = btb_198_tag == io_i_addr[12:3] ? btb_198_valid : _GEN_985; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_991 = btb_198_tag == io_i_addr[12:3] ? btb_198_target_address : _GEN_986; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_994 = btb_198_tag == io_i_addr[12:3] ? ~btb_198_bht[1] : _GEN_989; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_995 = btb_199_tag == io_i_addr[12:3] ? btb_199_valid : _GEN_990; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_996 = btb_199_tag == io_i_addr[12:3] ? btb_199_target_address : _GEN_991; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_999 = btb_199_tag == io_i_addr[12:3] ? ~btb_199_bht[1] : _GEN_994; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1000 = btb_200_tag == io_i_addr[12:3] ? btb_200_valid : _GEN_995; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1001 = btb_200_tag == io_i_addr[12:3] ? btb_200_target_address : _GEN_996; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1004 = btb_200_tag == io_i_addr[12:3] ? ~btb_200_bht[1] : _GEN_999; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1005 = btb_201_tag == io_i_addr[12:3] ? btb_201_valid : _GEN_1000; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1006 = btb_201_tag == io_i_addr[12:3] ? btb_201_target_address : _GEN_1001; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1009 = btb_201_tag == io_i_addr[12:3] ? ~btb_201_bht[1] : _GEN_1004; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1010 = btb_202_tag == io_i_addr[12:3] ? btb_202_valid : _GEN_1005; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1011 = btb_202_tag == io_i_addr[12:3] ? btb_202_target_address : _GEN_1006; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1014 = btb_202_tag == io_i_addr[12:3] ? ~btb_202_bht[1] : _GEN_1009; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1015 = btb_203_tag == io_i_addr[12:3] ? btb_203_valid : _GEN_1010; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1016 = btb_203_tag == io_i_addr[12:3] ? btb_203_target_address : _GEN_1011; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1019 = btb_203_tag == io_i_addr[12:3] ? ~btb_203_bht[1] : _GEN_1014; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1020 = btb_204_tag == io_i_addr[12:3] ? btb_204_valid : _GEN_1015; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1021 = btb_204_tag == io_i_addr[12:3] ? btb_204_target_address : _GEN_1016; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1024 = btb_204_tag == io_i_addr[12:3] ? ~btb_204_bht[1] : _GEN_1019; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1025 = btb_205_tag == io_i_addr[12:3] ? btb_205_valid : _GEN_1020; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1026 = btb_205_tag == io_i_addr[12:3] ? btb_205_target_address : _GEN_1021; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1029 = btb_205_tag == io_i_addr[12:3] ? ~btb_205_bht[1] : _GEN_1024; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1030 = btb_206_tag == io_i_addr[12:3] ? btb_206_valid : _GEN_1025; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1031 = btb_206_tag == io_i_addr[12:3] ? btb_206_target_address : _GEN_1026; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1034 = btb_206_tag == io_i_addr[12:3] ? ~btb_206_bht[1] : _GEN_1029; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1035 = btb_207_tag == io_i_addr[12:3] ? btb_207_valid : _GEN_1030; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1036 = btb_207_tag == io_i_addr[12:3] ? btb_207_target_address : _GEN_1031; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1039 = btb_207_tag == io_i_addr[12:3] ? ~btb_207_bht[1] : _GEN_1034; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1040 = btb_208_tag == io_i_addr[12:3] ? btb_208_valid : _GEN_1035; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1041 = btb_208_tag == io_i_addr[12:3] ? btb_208_target_address : _GEN_1036; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1044 = btb_208_tag == io_i_addr[12:3] ? ~btb_208_bht[1] : _GEN_1039; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1045 = btb_209_tag == io_i_addr[12:3] ? btb_209_valid : _GEN_1040; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1046 = btb_209_tag == io_i_addr[12:3] ? btb_209_target_address : _GEN_1041; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1049 = btb_209_tag == io_i_addr[12:3] ? ~btb_209_bht[1] : _GEN_1044; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1050 = btb_210_tag == io_i_addr[12:3] ? btb_210_valid : _GEN_1045; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1051 = btb_210_tag == io_i_addr[12:3] ? btb_210_target_address : _GEN_1046; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1054 = btb_210_tag == io_i_addr[12:3] ? ~btb_210_bht[1] : _GEN_1049; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1055 = btb_211_tag == io_i_addr[12:3] ? btb_211_valid : _GEN_1050; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1056 = btb_211_tag == io_i_addr[12:3] ? btb_211_target_address : _GEN_1051; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1059 = btb_211_tag == io_i_addr[12:3] ? ~btb_211_bht[1] : _GEN_1054; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1060 = btb_212_tag == io_i_addr[12:3] ? btb_212_valid : _GEN_1055; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1061 = btb_212_tag == io_i_addr[12:3] ? btb_212_target_address : _GEN_1056; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1064 = btb_212_tag == io_i_addr[12:3] ? ~btb_212_bht[1] : _GEN_1059; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1065 = btb_213_tag == io_i_addr[12:3] ? btb_213_valid : _GEN_1060; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1066 = btb_213_tag == io_i_addr[12:3] ? btb_213_target_address : _GEN_1061; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1069 = btb_213_tag == io_i_addr[12:3] ? ~btb_213_bht[1] : _GEN_1064; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1070 = btb_214_tag == io_i_addr[12:3] ? btb_214_valid : _GEN_1065; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1071 = btb_214_tag == io_i_addr[12:3] ? btb_214_target_address : _GEN_1066; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1074 = btb_214_tag == io_i_addr[12:3] ? ~btb_214_bht[1] : _GEN_1069; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1075 = btb_215_tag == io_i_addr[12:3] ? btb_215_valid : _GEN_1070; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1076 = btb_215_tag == io_i_addr[12:3] ? btb_215_target_address : _GEN_1071; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1079 = btb_215_tag == io_i_addr[12:3] ? ~btb_215_bht[1] : _GEN_1074; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1080 = btb_216_tag == io_i_addr[12:3] ? btb_216_valid : _GEN_1075; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1081 = btb_216_tag == io_i_addr[12:3] ? btb_216_target_address : _GEN_1076; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1084 = btb_216_tag == io_i_addr[12:3] ? ~btb_216_bht[1] : _GEN_1079; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1085 = btb_217_tag == io_i_addr[12:3] ? btb_217_valid : _GEN_1080; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1086 = btb_217_tag == io_i_addr[12:3] ? btb_217_target_address : _GEN_1081; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1089 = btb_217_tag == io_i_addr[12:3] ? ~btb_217_bht[1] : _GEN_1084; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1090 = btb_218_tag == io_i_addr[12:3] ? btb_218_valid : _GEN_1085; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1091 = btb_218_tag == io_i_addr[12:3] ? btb_218_target_address : _GEN_1086; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1094 = btb_218_tag == io_i_addr[12:3] ? ~btb_218_bht[1] : _GEN_1089; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1095 = btb_219_tag == io_i_addr[12:3] ? btb_219_valid : _GEN_1090; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1096 = btb_219_tag == io_i_addr[12:3] ? btb_219_target_address : _GEN_1091; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1099 = btb_219_tag == io_i_addr[12:3] ? ~btb_219_bht[1] : _GEN_1094; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1100 = btb_220_tag == io_i_addr[12:3] ? btb_220_valid : _GEN_1095; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1101 = btb_220_tag == io_i_addr[12:3] ? btb_220_target_address : _GEN_1096; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1104 = btb_220_tag == io_i_addr[12:3] ? ~btb_220_bht[1] : _GEN_1099; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1105 = btb_221_tag == io_i_addr[12:3] ? btb_221_valid : _GEN_1100; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1106 = btb_221_tag == io_i_addr[12:3] ? btb_221_target_address : _GEN_1101; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1109 = btb_221_tag == io_i_addr[12:3] ? ~btb_221_bht[1] : _GEN_1104; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1110 = btb_222_tag == io_i_addr[12:3] ? btb_222_valid : _GEN_1105; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1111 = btb_222_tag == io_i_addr[12:3] ? btb_222_target_address : _GEN_1106; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1114 = btb_222_tag == io_i_addr[12:3] ? ~btb_222_bht[1] : _GEN_1109; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1115 = btb_223_tag == io_i_addr[12:3] ? btb_223_valid : _GEN_1110; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1116 = btb_223_tag == io_i_addr[12:3] ? btb_223_target_address : _GEN_1111; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1119 = btb_223_tag == io_i_addr[12:3] ? ~btb_223_bht[1] : _GEN_1114; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1120 = btb_224_tag == io_i_addr[12:3] ? btb_224_valid : _GEN_1115; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1121 = btb_224_tag == io_i_addr[12:3] ? btb_224_target_address : _GEN_1116; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1124 = btb_224_tag == io_i_addr[12:3] ? ~btb_224_bht[1] : _GEN_1119; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1125 = btb_225_tag == io_i_addr[12:3] ? btb_225_valid : _GEN_1120; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1126 = btb_225_tag == io_i_addr[12:3] ? btb_225_target_address : _GEN_1121; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1129 = btb_225_tag == io_i_addr[12:3] ? ~btb_225_bht[1] : _GEN_1124; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1130 = btb_226_tag == io_i_addr[12:3] ? btb_226_valid : _GEN_1125; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1131 = btb_226_tag == io_i_addr[12:3] ? btb_226_target_address : _GEN_1126; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1134 = btb_226_tag == io_i_addr[12:3] ? ~btb_226_bht[1] : _GEN_1129; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1135 = btb_227_tag == io_i_addr[12:3] ? btb_227_valid : _GEN_1130; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1136 = btb_227_tag == io_i_addr[12:3] ? btb_227_target_address : _GEN_1131; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1139 = btb_227_tag == io_i_addr[12:3] ? ~btb_227_bht[1] : _GEN_1134; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1140 = btb_228_tag == io_i_addr[12:3] ? btb_228_valid : _GEN_1135; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1141 = btb_228_tag == io_i_addr[12:3] ? btb_228_target_address : _GEN_1136; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1144 = btb_228_tag == io_i_addr[12:3] ? ~btb_228_bht[1] : _GEN_1139; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1145 = btb_229_tag == io_i_addr[12:3] ? btb_229_valid : _GEN_1140; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1146 = btb_229_tag == io_i_addr[12:3] ? btb_229_target_address : _GEN_1141; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1149 = btb_229_tag == io_i_addr[12:3] ? ~btb_229_bht[1] : _GEN_1144; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1150 = btb_230_tag == io_i_addr[12:3] ? btb_230_valid : _GEN_1145; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1151 = btb_230_tag == io_i_addr[12:3] ? btb_230_target_address : _GEN_1146; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1154 = btb_230_tag == io_i_addr[12:3] ? ~btb_230_bht[1] : _GEN_1149; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1155 = btb_231_tag == io_i_addr[12:3] ? btb_231_valid : _GEN_1150; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1156 = btb_231_tag == io_i_addr[12:3] ? btb_231_target_address : _GEN_1151; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1159 = btb_231_tag == io_i_addr[12:3] ? ~btb_231_bht[1] : _GEN_1154; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1160 = btb_232_tag == io_i_addr[12:3] ? btb_232_valid : _GEN_1155; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1161 = btb_232_tag == io_i_addr[12:3] ? btb_232_target_address : _GEN_1156; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1164 = btb_232_tag == io_i_addr[12:3] ? ~btb_232_bht[1] : _GEN_1159; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1165 = btb_233_tag == io_i_addr[12:3] ? btb_233_valid : _GEN_1160; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1166 = btb_233_tag == io_i_addr[12:3] ? btb_233_target_address : _GEN_1161; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1169 = btb_233_tag == io_i_addr[12:3] ? ~btb_233_bht[1] : _GEN_1164; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1170 = btb_234_tag == io_i_addr[12:3] ? btb_234_valid : _GEN_1165; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1171 = btb_234_tag == io_i_addr[12:3] ? btb_234_target_address : _GEN_1166; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1174 = btb_234_tag == io_i_addr[12:3] ? ~btb_234_bht[1] : _GEN_1169; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1175 = btb_235_tag == io_i_addr[12:3] ? btb_235_valid : _GEN_1170; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1176 = btb_235_tag == io_i_addr[12:3] ? btb_235_target_address : _GEN_1171; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1179 = btb_235_tag == io_i_addr[12:3] ? ~btb_235_bht[1] : _GEN_1174; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1180 = btb_236_tag == io_i_addr[12:3] ? btb_236_valid : _GEN_1175; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1181 = btb_236_tag == io_i_addr[12:3] ? btb_236_target_address : _GEN_1176; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1184 = btb_236_tag == io_i_addr[12:3] ? ~btb_236_bht[1] : _GEN_1179; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1185 = btb_237_tag == io_i_addr[12:3] ? btb_237_valid : _GEN_1180; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1186 = btb_237_tag == io_i_addr[12:3] ? btb_237_target_address : _GEN_1181; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1189 = btb_237_tag == io_i_addr[12:3] ? ~btb_237_bht[1] : _GEN_1184; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1190 = btb_238_tag == io_i_addr[12:3] ? btb_238_valid : _GEN_1185; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1191 = btb_238_tag == io_i_addr[12:3] ? btb_238_target_address : _GEN_1186; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1194 = btb_238_tag == io_i_addr[12:3] ? ~btb_238_bht[1] : _GEN_1189; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1195 = btb_239_tag == io_i_addr[12:3] ? btb_239_valid : _GEN_1190; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1196 = btb_239_tag == io_i_addr[12:3] ? btb_239_target_address : _GEN_1191; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1199 = btb_239_tag == io_i_addr[12:3] ? ~btb_239_bht[1] : _GEN_1194; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1200 = btb_240_tag == io_i_addr[12:3] ? btb_240_valid : _GEN_1195; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1201 = btb_240_tag == io_i_addr[12:3] ? btb_240_target_address : _GEN_1196; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1204 = btb_240_tag == io_i_addr[12:3] ? ~btb_240_bht[1] : _GEN_1199; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1205 = btb_241_tag == io_i_addr[12:3] ? btb_241_valid : _GEN_1200; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1206 = btb_241_tag == io_i_addr[12:3] ? btb_241_target_address : _GEN_1201; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1209 = btb_241_tag == io_i_addr[12:3] ? ~btb_241_bht[1] : _GEN_1204; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1210 = btb_242_tag == io_i_addr[12:3] ? btb_242_valid : _GEN_1205; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1211 = btb_242_tag == io_i_addr[12:3] ? btb_242_target_address : _GEN_1206; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1214 = btb_242_tag == io_i_addr[12:3] ? ~btb_242_bht[1] : _GEN_1209; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1215 = btb_243_tag == io_i_addr[12:3] ? btb_243_valid : _GEN_1210; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1216 = btb_243_tag == io_i_addr[12:3] ? btb_243_target_address : _GEN_1211; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1219 = btb_243_tag == io_i_addr[12:3] ? ~btb_243_bht[1] : _GEN_1214; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1220 = btb_244_tag == io_i_addr[12:3] ? btb_244_valid : _GEN_1215; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1221 = btb_244_tag == io_i_addr[12:3] ? btb_244_target_address : _GEN_1216; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1224 = btb_244_tag == io_i_addr[12:3] ? ~btb_244_bht[1] : _GEN_1219; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1225 = btb_245_tag == io_i_addr[12:3] ? btb_245_valid : _GEN_1220; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1226 = btb_245_tag == io_i_addr[12:3] ? btb_245_target_address : _GEN_1221; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1229 = btb_245_tag == io_i_addr[12:3] ? ~btb_245_bht[1] : _GEN_1224; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1230 = btb_246_tag == io_i_addr[12:3] ? btb_246_valid : _GEN_1225; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1231 = btb_246_tag == io_i_addr[12:3] ? btb_246_target_address : _GEN_1226; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1234 = btb_246_tag == io_i_addr[12:3] ? ~btb_246_bht[1] : _GEN_1229; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1235 = btb_247_tag == io_i_addr[12:3] ? btb_247_valid : _GEN_1230; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1236 = btb_247_tag == io_i_addr[12:3] ? btb_247_target_address : _GEN_1231; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1239 = btb_247_tag == io_i_addr[12:3] ? ~btb_247_bht[1] : _GEN_1234; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1240 = btb_248_tag == io_i_addr[12:3] ? btb_248_valid : _GEN_1235; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1241 = btb_248_tag == io_i_addr[12:3] ? btb_248_target_address : _GEN_1236; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1244 = btb_248_tag == io_i_addr[12:3] ? ~btb_248_bht[1] : _GEN_1239; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1245 = btb_249_tag == io_i_addr[12:3] ? btb_249_valid : _GEN_1240; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1246 = btb_249_tag == io_i_addr[12:3] ? btb_249_target_address : _GEN_1241; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1249 = btb_249_tag == io_i_addr[12:3] ? ~btb_249_bht[1] : _GEN_1244; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1250 = btb_250_tag == io_i_addr[12:3] ? btb_250_valid : _GEN_1245; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1251 = btb_250_tag == io_i_addr[12:3] ? btb_250_target_address : _GEN_1246; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1254 = btb_250_tag == io_i_addr[12:3] ? ~btb_250_bht[1] : _GEN_1249; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1255 = btb_251_tag == io_i_addr[12:3] ? btb_251_valid : _GEN_1250; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1256 = btb_251_tag == io_i_addr[12:3] ? btb_251_target_address : _GEN_1251; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1259 = btb_251_tag == io_i_addr[12:3] ? ~btb_251_bht[1] : _GEN_1254; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1260 = btb_252_tag == io_i_addr[12:3] ? btb_252_valid : _GEN_1255; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1261 = btb_252_tag == io_i_addr[12:3] ? btb_252_target_address : _GEN_1256; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1264 = btb_252_tag == io_i_addr[12:3] ? ~btb_252_bht[1] : _GEN_1259; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1265 = btb_253_tag == io_i_addr[12:3] ? btb_253_valid : _GEN_1260; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1266 = btb_253_tag == io_i_addr[12:3] ? btb_253_target_address : _GEN_1261; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1269 = btb_253_tag == io_i_addr[12:3] ? ~btb_253_bht[1] : _GEN_1264; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1270 = btb_254_tag == io_i_addr[12:3] ? btb_254_valid : _GEN_1265; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1271 = btb_254_tag == io_i_addr[12:3] ? btb_254_target_address : _GEN_1266; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1274 = btb_254_tag == io_i_addr[12:3] ? ~btb_254_bht[1] : _GEN_1269; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1275 = btb_255_tag == io_i_addr[12:3] ? btb_255_valid : _GEN_1270; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1276 = btb_255_tag == io_i_addr[12:3] ? btb_255_target_address : _GEN_1271; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1279 = btb_255_tag == io_i_addr[12:3] ? ~btb_255_bht[1] : _GEN_1274; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1280 = btb_256_tag == io_i_addr[12:3] ? btb_256_valid : _GEN_1275; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1281 = btb_256_tag == io_i_addr[12:3] ? btb_256_target_address : _GEN_1276; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1284 = btb_256_tag == io_i_addr[12:3] ? ~btb_256_bht[1] : _GEN_1279; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1285 = btb_257_tag == io_i_addr[12:3] ? btb_257_valid : _GEN_1280; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1286 = btb_257_tag == io_i_addr[12:3] ? btb_257_target_address : _GEN_1281; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1289 = btb_257_tag == io_i_addr[12:3] ? ~btb_257_bht[1] : _GEN_1284; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1290 = btb_258_tag == io_i_addr[12:3] ? btb_258_valid : _GEN_1285; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1291 = btb_258_tag == io_i_addr[12:3] ? btb_258_target_address : _GEN_1286; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1294 = btb_258_tag == io_i_addr[12:3] ? ~btb_258_bht[1] : _GEN_1289; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1295 = btb_259_tag == io_i_addr[12:3] ? btb_259_valid : _GEN_1290; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1296 = btb_259_tag == io_i_addr[12:3] ? btb_259_target_address : _GEN_1291; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1299 = btb_259_tag == io_i_addr[12:3] ? ~btb_259_bht[1] : _GEN_1294; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1300 = btb_260_tag == io_i_addr[12:3] ? btb_260_valid : _GEN_1295; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1301 = btb_260_tag == io_i_addr[12:3] ? btb_260_target_address : _GEN_1296; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1304 = btb_260_tag == io_i_addr[12:3] ? ~btb_260_bht[1] : _GEN_1299; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1305 = btb_261_tag == io_i_addr[12:3] ? btb_261_valid : _GEN_1300; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1306 = btb_261_tag == io_i_addr[12:3] ? btb_261_target_address : _GEN_1301; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1309 = btb_261_tag == io_i_addr[12:3] ? ~btb_261_bht[1] : _GEN_1304; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1310 = btb_262_tag == io_i_addr[12:3] ? btb_262_valid : _GEN_1305; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1311 = btb_262_tag == io_i_addr[12:3] ? btb_262_target_address : _GEN_1306; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1314 = btb_262_tag == io_i_addr[12:3] ? ~btb_262_bht[1] : _GEN_1309; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1315 = btb_263_tag == io_i_addr[12:3] ? btb_263_valid : _GEN_1310; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1316 = btb_263_tag == io_i_addr[12:3] ? btb_263_target_address : _GEN_1311; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1319 = btb_263_tag == io_i_addr[12:3] ? ~btb_263_bht[1] : _GEN_1314; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1320 = btb_264_tag == io_i_addr[12:3] ? btb_264_valid : _GEN_1315; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1321 = btb_264_tag == io_i_addr[12:3] ? btb_264_target_address : _GEN_1316; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1324 = btb_264_tag == io_i_addr[12:3] ? ~btb_264_bht[1] : _GEN_1319; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1325 = btb_265_tag == io_i_addr[12:3] ? btb_265_valid : _GEN_1320; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1326 = btb_265_tag == io_i_addr[12:3] ? btb_265_target_address : _GEN_1321; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1329 = btb_265_tag == io_i_addr[12:3] ? ~btb_265_bht[1] : _GEN_1324; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1330 = btb_266_tag == io_i_addr[12:3] ? btb_266_valid : _GEN_1325; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1331 = btb_266_tag == io_i_addr[12:3] ? btb_266_target_address : _GEN_1326; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1334 = btb_266_tag == io_i_addr[12:3] ? ~btb_266_bht[1] : _GEN_1329; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1335 = btb_267_tag == io_i_addr[12:3] ? btb_267_valid : _GEN_1330; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1336 = btb_267_tag == io_i_addr[12:3] ? btb_267_target_address : _GEN_1331; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1339 = btb_267_tag == io_i_addr[12:3] ? ~btb_267_bht[1] : _GEN_1334; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1340 = btb_268_tag == io_i_addr[12:3] ? btb_268_valid : _GEN_1335; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1341 = btb_268_tag == io_i_addr[12:3] ? btb_268_target_address : _GEN_1336; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1344 = btb_268_tag == io_i_addr[12:3] ? ~btb_268_bht[1] : _GEN_1339; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1345 = btb_269_tag == io_i_addr[12:3] ? btb_269_valid : _GEN_1340; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1346 = btb_269_tag == io_i_addr[12:3] ? btb_269_target_address : _GEN_1341; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1349 = btb_269_tag == io_i_addr[12:3] ? ~btb_269_bht[1] : _GEN_1344; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1350 = btb_270_tag == io_i_addr[12:3] ? btb_270_valid : _GEN_1345; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1351 = btb_270_tag == io_i_addr[12:3] ? btb_270_target_address : _GEN_1346; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1354 = btb_270_tag == io_i_addr[12:3] ? ~btb_270_bht[1] : _GEN_1349; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1355 = btb_271_tag == io_i_addr[12:3] ? btb_271_valid : _GEN_1350; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1356 = btb_271_tag == io_i_addr[12:3] ? btb_271_target_address : _GEN_1351; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1359 = btb_271_tag == io_i_addr[12:3] ? ~btb_271_bht[1] : _GEN_1354; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1360 = btb_272_tag == io_i_addr[12:3] ? btb_272_valid : _GEN_1355; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1361 = btb_272_tag == io_i_addr[12:3] ? btb_272_target_address : _GEN_1356; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1364 = btb_272_tag == io_i_addr[12:3] ? ~btb_272_bht[1] : _GEN_1359; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1365 = btb_273_tag == io_i_addr[12:3] ? btb_273_valid : _GEN_1360; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1366 = btb_273_tag == io_i_addr[12:3] ? btb_273_target_address : _GEN_1361; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1369 = btb_273_tag == io_i_addr[12:3] ? ~btb_273_bht[1] : _GEN_1364; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1370 = btb_274_tag == io_i_addr[12:3] ? btb_274_valid : _GEN_1365; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1371 = btb_274_tag == io_i_addr[12:3] ? btb_274_target_address : _GEN_1366; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1374 = btb_274_tag == io_i_addr[12:3] ? ~btb_274_bht[1] : _GEN_1369; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1375 = btb_275_tag == io_i_addr[12:3] ? btb_275_valid : _GEN_1370; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1376 = btb_275_tag == io_i_addr[12:3] ? btb_275_target_address : _GEN_1371; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1379 = btb_275_tag == io_i_addr[12:3] ? ~btb_275_bht[1] : _GEN_1374; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1380 = btb_276_tag == io_i_addr[12:3] ? btb_276_valid : _GEN_1375; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1381 = btb_276_tag == io_i_addr[12:3] ? btb_276_target_address : _GEN_1376; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1384 = btb_276_tag == io_i_addr[12:3] ? ~btb_276_bht[1] : _GEN_1379; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1385 = btb_277_tag == io_i_addr[12:3] ? btb_277_valid : _GEN_1380; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1386 = btb_277_tag == io_i_addr[12:3] ? btb_277_target_address : _GEN_1381; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1389 = btb_277_tag == io_i_addr[12:3] ? ~btb_277_bht[1] : _GEN_1384; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1390 = btb_278_tag == io_i_addr[12:3] ? btb_278_valid : _GEN_1385; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1391 = btb_278_tag == io_i_addr[12:3] ? btb_278_target_address : _GEN_1386; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1394 = btb_278_tag == io_i_addr[12:3] ? ~btb_278_bht[1] : _GEN_1389; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1395 = btb_279_tag == io_i_addr[12:3] ? btb_279_valid : _GEN_1390; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1396 = btb_279_tag == io_i_addr[12:3] ? btb_279_target_address : _GEN_1391; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1399 = btb_279_tag == io_i_addr[12:3] ? ~btb_279_bht[1] : _GEN_1394; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1400 = btb_280_tag == io_i_addr[12:3] ? btb_280_valid : _GEN_1395; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1401 = btb_280_tag == io_i_addr[12:3] ? btb_280_target_address : _GEN_1396; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1404 = btb_280_tag == io_i_addr[12:3] ? ~btb_280_bht[1] : _GEN_1399; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1405 = btb_281_tag == io_i_addr[12:3] ? btb_281_valid : _GEN_1400; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1406 = btb_281_tag == io_i_addr[12:3] ? btb_281_target_address : _GEN_1401; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1409 = btb_281_tag == io_i_addr[12:3] ? ~btb_281_bht[1] : _GEN_1404; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1410 = btb_282_tag == io_i_addr[12:3] ? btb_282_valid : _GEN_1405; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1411 = btb_282_tag == io_i_addr[12:3] ? btb_282_target_address : _GEN_1406; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1414 = btb_282_tag == io_i_addr[12:3] ? ~btb_282_bht[1] : _GEN_1409; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1415 = btb_283_tag == io_i_addr[12:3] ? btb_283_valid : _GEN_1410; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1416 = btb_283_tag == io_i_addr[12:3] ? btb_283_target_address : _GEN_1411; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1419 = btb_283_tag == io_i_addr[12:3] ? ~btb_283_bht[1] : _GEN_1414; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1420 = btb_284_tag == io_i_addr[12:3] ? btb_284_valid : _GEN_1415; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1421 = btb_284_tag == io_i_addr[12:3] ? btb_284_target_address : _GEN_1416; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1424 = btb_284_tag == io_i_addr[12:3] ? ~btb_284_bht[1] : _GEN_1419; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1425 = btb_285_tag == io_i_addr[12:3] ? btb_285_valid : _GEN_1420; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1426 = btb_285_tag == io_i_addr[12:3] ? btb_285_target_address : _GEN_1421; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1429 = btb_285_tag == io_i_addr[12:3] ? ~btb_285_bht[1] : _GEN_1424; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1430 = btb_286_tag == io_i_addr[12:3] ? btb_286_valid : _GEN_1425; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1431 = btb_286_tag == io_i_addr[12:3] ? btb_286_target_address : _GEN_1426; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1434 = btb_286_tag == io_i_addr[12:3] ? ~btb_286_bht[1] : _GEN_1429; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1435 = btb_287_tag == io_i_addr[12:3] ? btb_287_valid : _GEN_1430; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1436 = btb_287_tag == io_i_addr[12:3] ? btb_287_target_address : _GEN_1431; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1439 = btb_287_tag == io_i_addr[12:3] ? ~btb_287_bht[1] : _GEN_1434; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1440 = btb_288_tag == io_i_addr[12:3] ? btb_288_valid : _GEN_1435; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1441 = btb_288_tag == io_i_addr[12:3] ? btb_288_target_address : _GEN_1436; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1444 = btb_288_tag == io_i_addr[12:3] ? ~btb_288_bht[1] : _GEN_1439; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1445 = btb_289_tag == io_i_addr[12:3] ? btb_289_valid : _GEN_1440; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1446 = btb_289_tag == io_i_addr[12:3] ? btb_289_target_address : _GEN_1441; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1449 = btb_289_tag == io_i_addr[12:3] ? ~btb_289_bht[1] : _GEN_1444; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1450 = btb_290_tag == io_i_addr[12:3] ? btb_290_valid : _GEN_1445; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1451 = btb_290_tag == io_i_addr[12:3] ? btb_290_target_address : _GEN_1446; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1454 = btb_290_tag == io_i_addr[12:3] ? ~btb_290_bht[1] : _GEN_1449; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1455 = btb_291_tag == io_i_addr[12:3] ? btb_291_valid : _GEN_1450; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1456 = btb_291_tag == io_i_addr[12:3] ? btb_291_target_address : _GEN_1451; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1459 = btb_291_tag == io_i_addr[12:3] ? ~btb_291_bht[1] : _GEN_1454; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1460 = btb_292_tag == io_i_addr[12:3] ? btb_292_valid : _GEN_1455; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1461 = btb_292_tag == io_i_addr[12:3] ? btb_292_target_address : _GEN_1456; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1464 = btb_292_tag == io_i_addr[12:3] ? ~btb_292_bht[1] : _GEN_1459; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1465 = btb_293_tag == io_i_addr[12:3] ? btb_293_valid : _GEN_1460; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1466 = btb_293_tag == io_i_addr[12:3] ? btb_293_target_address : _GEN_1461; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1469 = btb_293_tag == io_i_addr[12:3] ? ~btb_293_bht[1] : _GEN_1464; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1470 = btb_294_tag == io_i_addr[12:3] ? btb_294_valid : _GEN_1465; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1471 = btb_294_tag == io_i_addr[12:3] ? btb_294_target_address : _GEN_1466; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1474 = btb_294_tag == io_i_addr[12:3] ? ~btb_294_bht[1] : _GEN_1469; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1475 = btb_295_tag == io_i_addr[12:3] ? btb_295_valid : _GEN_1470; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1476 = btb_295_tag == io_i_addr[12:3] ? btb_295_target_address : _GEN_1471; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1479 = btb_295_tag == io_i_addr[12:3] ? ~btb_295_bht[1] : _GEN_1474; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1480 = btb_296_tag == io_i_addr[12:3] ? btb_296_valid : _GEN_1475; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1481 = btb_296_tag == io_i_addr[12:3] ? btb_296_target_address : _GEN_1476; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1484 = btb_296_tag == io_i_addr[12:3] ? ~btb_296_bht[1] : _GEN_1479; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1485 = btb_297_tag == io_i_addr[12:3] ? btb_297_valid : _GEN_1480; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1486 = btb_297_tag == io_i_addr[12:3] ? btb_297_target_address : _GEN_1481; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1489 = btb_297_tag == io_i_addr[12:3] ? ~btb_297_bht[1] : _GEN_1484; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1490 = btb_298_tag == io_i_addr[12:3] ? btb_298_valid : _GEN_1485; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1491 = btb_298_tag == io_i_addr[12:3] ? btb_298_target_address : _GEN_1486; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1494 = btb_298_tag == io_i_addr[12:3] ? ~btb_298_bht[1] : _GEN_1489; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1495 = btb_299_tag == io_i_addr[12:3] ? btb_299_valid : _GEN_1490; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1496 = btb_299_tag == io_i_addr[12:3] ? btb_299_target_address : _GEN_1491; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1499 = btb_299_tag == io_i_addr[12:3] ? ~btb_299_bht[1] : _GEN_1494; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1500 = btb_300_tag == io_i_addr[12:3] ? btb_300_valid : _GEN_1495; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1501 = btb_300_tag == io_i_addr[12:3] ? btb_300_target_address : _GEN_1496; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1504 = btb_300_tag == io_i_addr[12:3] ? ~btb_300_bht[1] : _GEN_1499; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1505 = btb_301_tag == io_i_addr[12:3] ? btb_301_valid : _GEN_1500; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1506 = btb_301_tag == io_i_addr[12:3] ? btb_301_target_address : _GEN_1501; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1509 = btb_301_tag == io_i_addr[12:3] ? ~btb_301_bht[1] : _GEN_1504; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1510 = btb_302_tag == io_i_addr[12:3] ? btb_302_valid : _GEN_1505; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1511 = btb_302_tag == io_i_addr[12:3] ? btb_302_target_address : _GEN_1506; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1514 = btb_302_tag == io_i_addr[12:3] ? ~btb_302_bht[1] : _GEN_1509; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1515 = btb_303_tag == io_i_addr[12:3] ? btb_303_valid : _GEN_1510; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1516 = btb_303_tag == io_i_addr[12:3] ? btb_303_target_address : _GEN_1511; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1519 = btb_303_tag == io_i_addr[12:3] ? ~btb_303_bht[1] : _GEN_1514; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1520 = btb_304_tag == io_i_addr[12:3] ? btb_304_valid : _GEN_1515; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1521 = btb_304_tag == io_i_addr[12:3] ? btb_304_target_address : _GEN_1516; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1524 = btb_304_tag == io_i_addr[12:3] ? ~btb_304_bht[1] : _GEN_1519; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1525 = btb_305_tag == io_i_addr[12:3] ? btb_305_valid : _GEN_1520; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1526 = btb_305_tag == io_i_addr[12:3] ? btb_305_target_address : _GEN_1521; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1529 = btb_305_tag == io_i_addr[12:3] ? ~btb_305_bht[1] : _GEN_1524; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1530 = btb_306_tag == io_i_addr[12:3] ? btb_306_valid : _GEN_1525; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1531 = btb_306_tag == io_i_addr[12:3] ? btb_306_target_address : _GEN_1526; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1534 = btb_306_tag == io_i_addr[12:3] ? ~btb_306_bht[1] : _GEN_1529; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1535 = btb_307_tag == io_i_addr[12:3] ? btb_307_valid : _GEN_1530; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1536 = btb_307_tag == io_i_addr[12:3] ? btb_307_target_address : _GEN_1531; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1539 = btb_307_tag == io_i_addr[12:3] ? ~btb_307_bht[1] : _GEN_1534; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1540 = btb_308_tag == io_i_addr[12:3] ? btb_308_valid : _GEN_1535; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1541 = btb_308_tag == io_i_addr[12:3] ? btb_308_target_address : _GEN_1536; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1544 = btb_308_tag == io_i_addr[12:3] ? ~btb_308_bht[1] : _GEN_1539; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1545 = btb_309_tag == io_i_addr[12:3] ? btb_309_valid : _GEN_1540; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1546 = btb_309_tag == io_i_addr[12:3] ? btb_309_target_address : _GEN_1541; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1549 = btb_309_tag == io_i_addr[12:3] ? ~btb_309_bht[1] : _GEN_1544; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1550 = btb_310_tag == io_i_addr[12:3] ? btb_310_valid : _GEN_1545; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1551 = btb_310_tag == io_i_addr[12:3] ? btb_310_target_address : _GEN_1546; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1554 = btb_310_tag == io_i_addr[12:3] ? ~btb_310_bht[1] : _GEN_1549; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1555 = btb_311_tag == io_i_addr[12:3] ? btb_311_valid : _GEN_1550; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1556 = btb_311_tag == io_i_addr[12:3] ? btb_311_target_address : _GEN_1551; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1559 = btb_311_tag == io_i_addr[12:3] ? ~btb_311_bht[1] : _GEN_1554; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1560 = btb_312_tag == io_i_addr[12:3] ? btb_312_valid : _GEN_1555; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1561 = btb_312_tag == io_i_addr[12:3] ? btb_312_target_address : _GEN_1556; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1564 = btb_312_tag == io_i_addr[12:3] ? ~btb_312_bht[1] : _GEN_1559; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1565 = btb_313_tag == io_i_addr[12:3] ? btb_313_valid : _GEN_1560; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1566 = btb_313_tag == io_i_addr[12:3] ? btb_313_target_address : _GEN_1561; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1569 = btb_313_tag == io_i_addr[12:3] ? ~btb_313_bht[1] : _GEN_1564; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1570 = btb_314_tag == io_i_addr[12:3] ? btb_314_valid : _GEN_1565; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1571 = btb_314_tag == io_i_addr[12:3] ? btb_314_target_address : _GEN_1566; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1574 = btb_314_tag == io_i_addr[12:3] ? ~btb_314_bht[1] : _GEN_1569; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1575 = btb_315_tag == io_i_addr[12:3] ? btb_315_valid : _GEN_1570; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1576 = btb_315_tag == io_i_addr[12:3] ? btb_315_target_address : _GEN_1571; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1579 = btb_315_tag == io_i_addr[12:3] ? ~btb_315_bht[1] : _GEN_1574; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1580 = btb_316_tag == io_i_addr[12:3] ? btb_316_valid : _GEN_1575; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1581 = btb_316_tag == io_i_addr[12:3] ? btb_316_target_address : _GEN_1576; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1584 = btb_316_tag == io_i_addr[12:3] ? ~btb_316_bht[1] : _GEN_1579; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1585 = btb_317_tag == io_i_addr[12:3] ? btb_317_valid : _GEN_1580; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1586 = btb_317_tag == io_i_addr[12:3] ? btb_317_target_address : _GEN_1581; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1589 = btb_317_tag == io_i_addr[12:3] ? ~btb_317_bht[1] : _GEN_1584; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1590 = btb_318_tag == io_i_addr[12:3] ? btb_318_valid : _GEN_1585; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1591 = btb_318_tag == io_i_addr[12:3] ? btb_318_target_address : _GEN_1586; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1594 = btb_318_tag == io_i_addr[12:3] ? ~btb_318_bht[1] : _GEN_1589; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1595 = btb_319_tag == io_i_addr[12:3] ? btb_319_valid : _GEN_1590; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1596 = btb_319_tag == io_i_addr[12:3] ? btb_319_target_address : _GEN_1591; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1599 = btb_319_tag == io_i_addr[12:3] ? ~btb_319_bht[1] : _GEN_1594; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1600 = btb_320_tag == io_i_addr[12:3] ? btb_320_valid : _GEN_1595; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1601 = btb_320_tag == io_i_addr[12:3] ? btb_320_target_address : _GEN_1596; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1604 = btb_320_tag == io_i_addr[12:3] ? ~btb_320_bht[1] : _GEN_1599; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1605 = btb_321_tag == io_i_addr[12:3] ? btb_321_valid : _GEN_1600; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1606 = btb_321_tag == io_i_addr[12:3] ? btb_321_target_address : _GEN_1601; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1609 = btb_321_tag == io_i_addr[12:3] ? ~btb_321_bht[1] : _GEN_1604; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1610 = btb_322_tag == io_i_addr[12:3] ? btb_322_valid : _GEN_1605; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1611 = btb_322_tag == io_i_addr[12:3] ? btb_322_target_address : _GEN_1606; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1614 = btb_322_tag == io_i_addr[12:3] ? ~btb_322_bht[1] : _GEN_1609; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1615 = btb_323_tag == io_i_addr[12:3] ? btb_323_valid : _GEN_1610; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1616 = btb_323_tag == io_i_addr[12:3] ? btb_323_target_address : _GEN_1611; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1619 = btb_323_tag == io_i_addr[12:3] ? ~btb_323_bht[1] : _GEN_1614; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1620 = btb_324_tag == io_i_addr[12:3] ? btb_324_valid : _GEN_1615; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1621 = btb_324_tag == io_i_addr[12:3] ? btb_324_target_address : _GEN_1616; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1624 = btb_324_tag == io_i_addr[12:3] ? ~btb_324_bht[1] : _GEN_1619; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1625 = btb_325_tag == io_i_addr[12:3] ? btb_325_valid : _GEN_1620; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1626 = btb_325_tag == io_i_addr[12:3] ? btb_325_target_address : _GEN_1621; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1629 = btb_325_tag == io_i_addr[12:3] ? ~btb_325_bht[1] : _GEN_1624; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1630 = btb_326_tag == io_i_addr[12:3] ? btb_326_valid : _GEN_1625; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1631 = btb_326_tag == io_i_addr[12:3] ? btb_326_target_address : _GEN_1626; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1634 = btb_326_tag == io_i_addr[12:3] ? ~btb_326_bht[1] : _GEN_1629; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1635 = btb_327_tag == io_i_addr[12:3] ? btb_327_valid : _GEN_1630; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1636 = btb_327_tag == io_i_addr[12:3] ? btb_327_target_address : _GEN_1631; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1639 = btb_327_tag == io_i_addr[12:3] ? ~btb_327_bht[1] : _GEN_1634; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1640 = btb_328_tag == io_i_addr[12:3] ? btb_328_valid : _GEN_1635; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1641 = btb_328_tag == io_i_addr[12:3] ? btb_328_target_address : _GEN_1636; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1644 = btb_328_tag == io_i_addr[12:3] ? ~btb_328_bht[1] : _GEN_1639; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1645 = btb_329_tag == io_i_addr[12:3] ? btb_329_valid : _GEN_1640; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1646 = btb_329_tag == io_i_addr[12:3] ? btb_329_target_address : _GEN_1641; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1649 = btb_329_tag == io_i_addr[12:3] ? ~btb_329_bht[1] : _GEN_1644; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1650 = btb_330_tag == io_i_addr[12:3] ? btb_330_valid : _GEN_1645; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1651 = btb_330_tag == io_i_addr[12:3] ? btb_330_target_address : _GEN_1646; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1654 = btb_330_tag == io_i_addr[12:3] ? ~btb_330_bht[1] : _GEN_1649; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1655 = btb_331_tag == io_i_addr[12:3] ? btb_331_valid : _GEN_1650; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1656 = btb_331_tag == io_i_addr[12:3] ? btb_331_target_address : _GEN_1651; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1659 = btb_331_tag == io_i_addr[12:3] ? ~btb_331_bht[1] : _GEN_1654; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1660 = btb_332_tag == io_i_addr[12:3] ? btb_332_valid : _GEN_1655; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1661 = btb_332_tag == io_i_addr[12:3] ? btb_332_target_address : _GEN_1656; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1664 = btb_332_tag == io_i_addr[12:3] ? ~btb_332_bht[1] : _GEN_1659; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1665 = btb_333_tag == io_i_addr[12:3] ? btb_333_valid : _GEN_1660; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1666 = btb_333_tag == io_i_addr[12:3] ? btb_333_target_address : _GEN_1661; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1669 = btb_333_tag == io_i_addr[12:3] ? ~btb_333_bht[1] : _GEN_1664; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1670 = btb_334_tag == io_i_addr[12:3] ? btb_334_valid : _GEN_1665; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1671 = btb_334_tag == io_i_addr[12:3] ? btb_334_target_address : _GEN_1666; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1674 = btb_334_tag == io_i_addr[12:3] ? ~btb_334_bht[1] : _GEN_1669; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1675 = btb_335_tag == io_i_addr[12:3] ? btb_335_valid : _GEN_1670; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1676 = btb_335_tag == io_i_addr[12:3] ? btb_335_target_address : _GEN_1671; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1679 = btb_335_tag == io_i_addr[12:3] ? ~btb_335_bht[1] : _GEN_1674; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1680 = btb_336_tag == io_i_addr[12:3] ? btb_336_valid : _GEN_1675; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1681 = btb_336_tag == io_i_addr[12:3] ? btb_336_target_address : _GEN_1676; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1684 = btb_336_tag == io_i_addr[12:3] ? ~btb_336_bht[1] : _GEN_1679; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1685 = btb_337_tag == io_i_addr[12:3] ? btb_337_valid : _GEN_1680; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1686 = btb_337_tag == io_i_addr[12:3] ? btb_337_target_address : _GEN_1681; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1689 = btb_337_tag == io_i_addr[12:3] ? ~btb_337_bht[1] : _GEN_1684; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1690 = btb_338_tag == io_i_addr[12:3] ? btb_338_valid : _GEN_1685; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1691 = btb_338_tag == io_i_addr[12:3] ? btb_338_target_address : _GEN_1686; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1694 = btb_338_tag == io_i_addr[12:3] ? ~btb_338_bht[1] : _GEN_1689; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1695 = btb_339_tag == io_i_addr[12:3] ? btb_339_valid : _GEN_1690; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1696 = btb_339_tag == io_i_addr[12:3] ? btb_339_target_address : _GEN_1691; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1699 = btb_339_tag == io_i_addr[12:3] ? ~btb_339_bht[1] : _GEN_1694; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1700 = btb_340_tag == io_i_addr[12:3] ? btb_340_valid : _GEN_1695; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1701 = btb_340_tag == io_i_addr[12:3] ? btb_340_target_address : _GEN_1696; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1704 = btb_340_tag == io_i_addr[12:3] ? ~btb_340_bht[1] : _GEN_1699; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1705 = btb_341_tag == io_i_addr[12:3] ? btb_341_valid : _GEN_1700; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1706 = btb_341_tag == io_i_addr[12:3] ? btb_341_target_address : _GEN_1701; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1709 = btb_341_tag == io_i_addr[12:3] ? ~btb_341_bht[1] : _GEN_1704; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1710 = btb_342_tag == io_i_addr[12:3] ? btb_342_valid : _GEN_1705; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1711 = btb_342_tag == io_i_addr[12:3] ? btb_342_target_address : _GEN_1706; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1714 = btb_342_tag == io_i_addr[12:3] ? ~btb_342_bht[1] : _GEN_1709; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1715 = btb_343_tag == io_i_addr[12:3] ? btb_343_valid : _GEN_1710; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1716 = btb_343_tag == io_i_addr[12:3] ? btb_343_target_address : _GEN_1711; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1719 = btb_343_tag == io_i_addr[12:3] ? ~btb_343_bht[1] : _GEN_1714; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1720 = btb_344_tag == io_i_addr[12:3] ? btb_344_valid : _GEN_1715; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1721 = btb_344_tag == io_i_addr[12:3] ? btb_344_target_address : _GEN_1716; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1724 = btb_344_tag == io_i_addr[12:3] ? ~btb_344_bht[1] : _GEN_1719; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1725 = btb_345_tag == io_i_addr[12:3] ? btb_345_valid : _GEN_1720; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1726 = btb_345_tag == io_i_addr[12:3] ? btb_345_target_address : _GEN_1721; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1729 = btb_345_tag == io_i_addr[12:3] ? ~btb_345_bht[1] : _GEN_1724; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1730 = btb_346_tag == io_i_addr[12:3] ? btb_346_valid : _GEN_1725; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1731 = btb_346_tag == io_i_addr[12:3] ? btb_346_target_address : _GEN_1726; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1734 = btb_346_tag == io_i_addr[12:3] ? ~btb_346_bht[1] : _GEN_1729; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1735 = btb_347_tag == io_i_addr[12:3] ? btb_347_valid : _GEN_1730; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1736 = btb_347_tag == io_i_addr[12:3] ? btb_347_target_address : _GEN_1731; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1739 = btb_347_tag == io_i_addr[12:3] ? ~btb_347_bht[1] : _GEN_1734; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1740 = btb_348_tag == io_i_addr[12:3] ? btb_348_valid : _GEN_1735; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1741 = btb_348_tag == io_i_addr[12:3] ? btb_348_target_address : _GEN_1736; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1744 = btb_348_tag == io_i_addr[12:3] ? ~btb_348_bht[1] : _GEN_1739; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1745 = btb_349_tag == io_i_addr[12:3] ? btb_349_valid : _GEN_1740; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1746 = btb_349_tag == io_i_addr[12:3] ? btb_349_target_address : _GEN_1741; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1749 = btb_349_tag == io_i_addr[12:3] ? ~btb_349_bht[1] : _GEN_1744; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1750 = btb_350_tag == io_i_addr[12:3] ? btb_350_valid : _GEN_1745; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1751 = btb_350_tag == io_i_addr[12:3] ? btb_350_target_address : _GEN_1746; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1754 = btb_350_tag == io_i_addr[12:3] ? ~btb_350_bht[1] : _GEN_1749; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1755 = btb_351_tag == io_i_addr[12:3] ? btb_351_valid : _GEN_1750; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1756 = btb_351_tag == io_i_addr[12:3] ? btb_351_target_address : _GEN_1751; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1759 = btb_351_tag == io_i_addr[12:3] ? ~btb_351_bht[1] : _GEN_1754; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1760 = btb_352_tag == io_i_addr[12:3] ? btb_352_valid : _GEN_1755; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1761 = btb_352_tag == io_i_addr[12:3] ? btb_352_target_address : _GEN_1756; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1764 = btb_352_tag == io_i_addr[12:3] ? ~btb_352_bht[1] : _GEN_1759; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1765 = btb_353_tag == io_i_addr[12:3] ? btb_353_valid : _GEN_1760; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1766 = btb_353_tag == io_i_addr[12:3] ? btb_353_target_address : _GEN_1761; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1769 = btb_353_tag == io_i_addr[12:3] ? ~btb_353_bht[1] : _GEN_1764; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1770 = btb_354_tag == io_i_addr[12:3] ? btb_354_valid : _GEN_1765; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1771 = btb_354_tag == io_i_addr[12:3] ? btb_354_target_address : _GEN_1766; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1774 = btb_354_tag == io_i_addr[12:3] ? ~btb_354_bht[1] : _GEN_1769; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1775 = btb_355_tag == io_i_addr[12:3] ? btb_355_valid : _GEN_1770; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1776 = btb_355_tag == io_i_addr[12:3] ? btb_355_target_address : _GEN_1771; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1779 = btb_355_tag == io_i_addr[12:3] ? ~btb_355_bht[1] : _GEN_1774; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1780 = btb_356_tag == io_i_addr[12:3] ? btb_356_valid : _GEN_1775; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1781 = btb_356_tag == io_i_addr[12:3] ? btb_356_target_address : _GEN_1776; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1784 = btb_356_tag == io_i_addr[12:3] ? ~btb_356_bht[1] : _GEN_1779; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1785 = btb_357_tag == io_i_addr[12:3] ? btb_357_valid : _GEN_1780; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1786 = btb_357_tag == io_i_addr[12:3] ? btb_357_target_address : _GEN_1781; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1789 = btb_357_tag == io_i_addr[12:3] ? ~btb_357_bht[1] : _GEN_1784; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1790 = btb_358_tag == io_i_addr[12:3] ? btb_358_valid : _GEN_1785; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1791 = btb_358_tag == io_i_addr[12:3] ? btb_358_target_address : _GEN_1786; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1794 = btb_358_tag == io_i_addr[12:3] ? ~btb_358_bht[1] : _GEN_1789; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1795 = btb_359_tag == io_i_addr[12:3] ? btb_359_valid : _GEN_1790; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1796 = btb_359_tag == io_i_addr[12:3] ? btb_359_target_address : _GEN_1791; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1799 = btb_359_tag == io_i_addr[12:3] ? ~btb_359_bht[1] : _GEN_1794; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1800 = btb_360_tag == io_i_addr[12:3] ? btb_360_valid : _GEN_1795; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1801 = btb_360_tag == io_i_addr[12:3] ? btb_360_target_address : _GEN_1796; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1804 = btb_360_tag == io_i_addr[12:3] ? ~btb_360_bht[1] : _GEN_1799; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1805 = btb_361_tag == io_i_addr[12:3] ? btb_361_valid : _GEN_1800; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1806 = btb_361_tag == io_i_addr[12:3] ? btb_361_target_address : _GEN_1801; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1809 = btb_361_tag == io_i_addr[12:3] ? ~btb_361_bht[1] : _GEN_1804; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1810 = btb_362_tag == io_i_addr[12:3] ? btb_362_valid : _GEN_1805; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1811 = btb_362_tag == io_i_addr[12:3] ? btb_362_target_address : _GEN_1806; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1814 = btb_362_tag == io_i_addr[12:3] ? ~btb_362_bht[1] : _GEN_1809; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1815 = btb_363_tag == io_i_addr[12:3] ? btb_363_valid : _GEN_1810; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1816 = btb_363_tag == io_i_addr[12:3] ? btb_363_target_address : _GEN_1811; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1819 = btb_363_tag == io_i_addr[12:3] ? ~btb_363_bht[1] : _GEN_1814; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1820 = btb_364_tag == io_i_addr[12:3] ? btb_364_valid : _GEN_1815; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1821 = btb_364_tag == io_i_addr[12:3] ? btb_364_target_address : _GEN_1816; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1824 = btb_364_tag == io_i_addr[12:3] ? ~btb_364_bht[1] : _GEN_1819; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1825 = btb_365_tag == io_i_addr[12:3] ? btb_365_valid : _GEN_1820; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1826 = btb_365_tag == io_i_addr[12:3] ? btb_365_target_address : _GEN_1821; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1829 = btb_365_tag == io_i_addr[12:3] ? ~btb_365_bht[1] : _GEN_1824; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1830 = btb_366_tag == io_i_addr[12:3] ? btb_366_valid : _GEN_1825; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1831 = btb_366_tag == io_i_addr[12:3] ? btb_366_target_address : _GEN_1826; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1834 = btb_366_tag == io_i_addr[12:3] ? ~btb_366_bht[1] : _GEN_1829; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1835 = btb_367_tag == io_i_addr[12:3] ? btb_367_valid : _GEN_1830; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1836 = btb_367_tag == io_i_addr[12:3] ? btb_367_target_address : _GEN_1831; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1839 = btb_367_tag == io_i_addr[12:3] ? ~btb_367_bht[1] : _GEN_1834; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1840 = btb_368_tag == io_i_addr[12:3] ? btb_368_valid : _GEN_1835; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1841 = btb_368_tag == io_i_addr[12:3] ? btb_368_target_address : _GEN_1836; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1844 = btb_368_tag == io_i_addr[12:3] ? ~btb_368_bht[1] : _GEN_1839; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1845 = btb_369_tag == io_i_addr[12:3] ? btb_369_valid : _GEN_1840; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1846 = btb_369_tag == io_i_addr[12:3] ? btb_369_target_address : _GEN_1841; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1849 = btb_369_tag == io_i_addr[12:3] ? ~btb_369_bht[1] : _GEN_1844; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1850 = btb_370_tag == io_i_addr[12:3] ? btb_370_valid : _GEN_1845; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1851 = btb_370_tag == io_i_addr[12:3] ? btb_370_target_address : _GEN_1846; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1854 = btb_370_tag == io_i_addr[12:3] ? ~btb_370_bht[1] : _GEN_1849; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1855 = btb_371_tag == io_i_addr[12:3] ? btb_371_valid : _GEN_1850; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1856 = btb_371_tag == io_i_addr[12:3] ? btb_371_target_address : _GEN_1851; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1859 = btb_371_tag == io_i_addr[12:3] ? ~btb_371_bht[1] : _GEN_1854; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1860 = btb_372_tag == io_i_addr[12:3] ? btb_372_valid : _GEN_1855; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1861 = btb_372_tag == io_i_addr[12:3] ? btb_372_target_address : _GEN_1856; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1864 = btb_372_tag == io_i_addr[12:3] ? ~btb_372_bht[1] : _GEN_1859; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1865 = btb_373_tag == io_i_addr[12:3] ? btb_373_valid : _GEN_1860; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1866 = btb_373_tag == io_i_addr[12:3] ? btb_373_target_address : _GEN_1861; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1869 = btb_373_tag == io_i_addr[12:3] ? ~btb_373_bht[1] : _GEN_1864; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1870 = btb_374_tag == io_i_addr[12:3] ? btb_374_valid : _GEN_1865; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1871 = btb_374_tag == io_i_addr[12:3] ? btb_374_target_address : _GEN_1866; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1874 = btb_374_tag == io_i_addr[12:3] ? ~btb_374_bht[1] : _GEN_1869; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1875 = btb_375_tag == io_i_addr[12:3] ? btb_375_valid : _GEN_1870; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1876 = btb_375_tag == io_i_addr[12:3] ? btb_375_target_address : _GEN_1871; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1879 = btb_375_tag == io_i_addr[12:3] ? ~btb_375_bht[1] : _GEN_1874; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1880 = btb_376_tag == io_i_addr[12:3] ? btb_376_valid : _GEN_1875; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1881 = btb_376_tag == io_i_addr[12:3] ? btb_376_target_address : _GEN_1876; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1884 = btb_376_tag == io_i_addr[12:3] ? ~btb_376_bht[1] : _GEN_1879; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1885 = btb_377_tag == io_i_addr[12:3] ? btb_377_valid : _GEN_1880; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1886 = btb_377_tag == io_i_addr[12:3] ? btb_377_target_address : _GEN_1881; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1889 = btb_377_tag == io_i_addr[12:3] ? ~btb_377_bht[1] : _GEN_1884; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1890 = btb_378_tag == io_i_addr[12:3] ? btb_378_valid : _GEN_1885; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1891 = btb_378_tag == io_i_addr[12:3] ? btb_378_target_address : _GEN_1886; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1894 = btb_378_tag == io_i_addr[12:3] ? ~btb_378_bht[1] : _GEN_1889; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1895 = btb_379_tag == io_i_addr[12:3] ? btb_379_valid : _GEN_1890; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1896 = btb_379_tag == io_i_addr[12:3] ? btb_379_target_address : _GEN_1891; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1899 = btb_379_tag == io_i_addr[12:3] ? ~btb_379_bht[1] : _GEN_1894; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1900 = btb_380_tag == io_i_addr[12:3] ? btb_380_valid : _GEN_1895; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1901 = btb_380_tag == io_i_addr[12:3] ? btb_380_target_address : _GEN_1896; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1904 = btb_380_tag == io_i_addr[12:3] ? ~btb_380_bht[1] : _GEN_1899; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1905 = btb_381_tag == io_i_addr[12:3] ? btb_381_valid : _GEN_1900; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1906 = btb_381_tag == io_i_addr[12:3] ? btb_381_target_address : _GEN_1901; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1909 = btb_381_tag == io_i_addr[12:3] ? ~btb_381_bht[1] : _GEN_1904; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1910 = btb_382_tag == io_i_addr[12:3] ? btb_382_valid : _GEN_1905; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1911 = btb_382_tag == io_i_addr[12:3] ? btb_382_target_address : _GEN_1906; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1914 = btb_382_tag == io_i_addr[12:3] ? ~btb_382_bht[1] : _GEN_1909; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1915 = btb_383_tag == io_i_addr[12:3] ? btb_383_valid : _GEN_1910; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1916 = btb_383_tag == io_i_addr[12:3] ? btb_383_target_address : _GEN_1911; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1919 = btb_383_tag == io_i_addr[12:3] ? ~btb_383_bht[1] : _GEN_1914; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1920 = btb_384_tag == io_i_addr[12:3] ? btb_384_valid : _GEN_1915; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1921 = btb_384_tag == io_i_addr[12:3] ? btb_384_target_address : _GEN_1916; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1924 = btb_384_tag == io_i_addr[12:3] ? ~btb_384_bht[1] : _GEN_1919; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1925 = btb_385_tag == io_i_addr[12:3] ? btb_385_valid : _GEN_1920; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1926 = btb_385_tag == io_i_addr[12:3] ? btb_385_target_address : _GEN_1921; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1929 = btb_385_tag == io_i_addr[12:3] ? ~btb_385_bht[1] : _GEN_1924; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1930 = btb_386_tag == io_i_addr[12:3] ? btb_386_valid : _GEN_1925; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1931 = btb_386_tag == io_i_addr[12:3] ? btb_386_target_address : _GEN_1926; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1934 = btb_386_tag == io_i_addr[12:3] ? ~btb_386_bht[1] : _GEN_1929; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1935 = btb_387_tag == io_i_addr[12:3] ? btb_387_valid : _GEN_1930; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1936 = btb_387_tag == io_i_addr[12:3] ? btb_387_target_address : _GEN_1931; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1939 = btb_387_tag == io_i_addr[12:3] ? ~btb_387_bht[1] : _GEN_1934; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1940 = btb_388_tag == io_i_addr[12:3] ? btb_388_valid : _GEN_1935; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1941 = btb_388_tag == io_i_addr[12:3] ? btb_388_target_address : _GEN_1936; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1944 = btb_388_tag == io_i_addr[12:3] ? ~btb_388_bht[1] : _GEN_1939; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1945 = btb_389_tag == io_i_addr[12:3] ? btb_389_valid : _GEN_1940; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1946 = btb_389_tag == io_i_addr[12:3] ? btb_389_target_address : _GEN_1941; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1949 = btb_389_tag == io_i_addr[12:3] ? ~btb_389_bht[1] : _GEN_1944; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1950 = btb_390_tag == io_i_addr[12:3] ? btb_390_valid : _GEN_1945; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1951 = btb_390_tag == io_i_addr[12:3] ? btb_390_target_address : _GEN_1946; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1954 = btb_390_tag == io_i_addr[12:3] ? ~btb_390_bht[1] : _GEN_1949; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1955 = btb_391_tag == io_i_addr[12:3] ? btb_391_valid : _GEN_1950; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1956 = btb_391_tag == io_i_addr[12:3] ? btb_391_target_address : _GEN_1951; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1959 = btb_391_tag == io_i_addr[12:3] ? ~btb_391_bht[1] : _GEN_1954; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1960 = btb_392_tag == io_i_addr[12:3] ? btb_392_valid : _GEN_1955; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1961 = btb_392_tag == io_i_addr[12:3] ? btb_392_target_address : _GEN_1956; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1964 = btb_392_tag == io_i_addr[12:3] ? ~btb_392_bht[1] : _GEN_1959; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1965 = btb_393_tag == io_i_addr[12:3] ? btb_393_valid : _GEN_1960; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1966 = btb_393_tag == io_i_addr[12:3] ? btb_393_target_address : _GEN_1961; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1969 = btb_393_tag == io_i_addr[12:3] ? ~btb_393_bht[1] : _GEN_1964; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1970 = btb_394_tag == io_i_addr[12:3] ? btb_394_valid : _GEN_1965; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1971 = btb_394_tag == io_i_addr[12:3] ? btb_394_target_address : _GEN_1966; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1974 = btb_394_tag == io_i_addr[12:3] ? ~btb_394_bht[1] : _GEN_1969; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1975 = btb_395_tag == io_i_addr[12:3] ? btb_395_valid : _GEN_1970; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1976 = btb_395_tag == io_i_addr[12:3] ? btb_395_target_address : _GEN_1971; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1979 = btb_395_tag == io_i_addr[12:3] ? ~btb_395_bht[1] : _GEN_1974; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1980 = btb_396_tag == io_i_addr[12:3] ? btb_396_valid : _GEN_1975; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1981 = btb_396_tag == io_i_addr[12:3] ? btb_396_target_address : _GEN_1976; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1984 = btb_396_tag == io_i_addr[12:3] ? ~btb_396_bht[1] : _GEN_1979; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1985 = btb_397_tag == io_i_addr[12:3] ? btb_397_valid : _GEN_1980; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1986 = btb_397_tag == io_i_addr[12:3] ? btb_397_target_address : _GEN_1981; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1989 = btb_397_tag == io_i_addr[12:3] ? ~btb_397_bht[1] : _GEN_1984; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1990 = btb_398_tag == io_i_addr[12:3] ? btb_398_valid : _GEN_1985; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1991 = btb_398_tag == io_i_addr[12:3] ? btb_398_target_address : _GEN_1986; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1994 = btb_398_tag == io_i_addr[12:3] ? ~btb_398_bht[1] : _GEN_1989; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_1995 = btb_399_tag == io_i_addr[12:3] ? btb_399_valid : _GEN_1990; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_1996 = btb_399_tag == io_i_addr[12:3] ? btb_399_target_address : _GEN_1991; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_1999 = btb_399_tag == io_i_addr[12:3] ? ~btb_399_bht[1] : _GEN_1994; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2000 = btb_400_tag == io_i_addr[12:3] ? btb_400_valid : _GEN_1995; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2001 = btb_400_tag == io_i_addr[12:3] ? btb_400_target_address : _GEN_1996; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2004 = btb_400_tag == io_i_addr[12:3] ? ~btb_400_bht[1] : _GEN_1999; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2005 = btb_401_tag == io_i_addr[12:3] ? btb_401_valid : _GEN_2000; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2006 = btb_401_tag == io_i_addr[12:3] ? btb_401_target_address : _GEN_2001; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2009 = btb_401_tag == io_i_addr[12:3] ? ~btb_401_bht[1] : _GEN_2004; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2010 = btb_402_tag == io_i_addr[12:3] ? btb_402_valid : _GEN_2005; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2011 = btb_402_tag == io_i_addr[12:3] ? btb_402_target_address : _GEN_2006; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2014 = btb_402_tag == io_i_addr[12:3] ? ~btb_402_bht[1] : _GEN_2009; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2015 = btb_403_tag == io_i_addr[12:3] ? btb_403_valid : _GEN_2010; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2016 = btb_403_tag == io_i_addr[12:3] ? btb_403_target_address : _GEN_2011; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2019 = btb_403_tag == io_i_addr[12:3] ? ~btb_403_bht[1] : _GEN_2014; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2020 = btb_404_tag == io_i_addr[12:3] ? btb_404_valid : _GEN_2015; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2021 = btb_404_tag == io_i_addr[12:3] ? btb_404_target_address : _GEN_2016; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2024 = btb_404_tag == io_i_addr[12:3] ? ~btb_404_bht[1] : _GEN_2019; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2025 = btb_405_tag == io_i_addr[12:3] ? btb_405_valid : _GEN_2020; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2026 = btb_405_tag == io_i_addr[12:3] ? btb_405_target_address : _GEN_2021; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2029 = btb_405_tag == io_i_addr[12:3] ? ~btb_405_bht[1] : _GEN_2024; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2030 = btb_406_tag == io_i_addr[12:3] ? btb_406_valid : _GEN_2025; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2031 = btb_406_tag == io_i_addr[12:3] ? btb_406_target_address : _GEN_2026; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2034 = btb_406_tag == io_i_addr[12:3] ? ~btb_406_bht[1] : _GEN_2029; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2035 = btb_407_tag == io_i_addr[12:3] ? btb_407_valid : _GEN_2030; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2036 = btb_407_tag == io_i_addr[12:3] ? btb_407_target_address : _GEN_2031; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2039 = btb_407_tag == io_i_addr[12:3] ? ~btb_407_bht[1] : _GEN_2034; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2040 = btb_408_tag == io_i_addr[12:3] ? btb_408_valid : _GEN_2035; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2041 = btb_408_tag == io_i_addr[12:3] ? btb_408_target_address : _GEN_2036; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2044 = btb_408_tag == io_i_addr[12:3] ? ~btb_408_bht[1] : _GEN_2039; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2045 = btb_409_tag == io_i_addr[12:3] ? btb_409_valid : _GEN_2040; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2046 = btb_409_tag == io_i_addr[12:3] ? btb_409_target_address : _GEN_2041; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2049 = btb_409_tag == io_i_addr[12:3] ? ~btb_409_bht[1] : _GEN_2044; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2050 = btb_410_tag == io_i_addr[12:3] ? btb_410_valid : _GEN_2045; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2051 = btb_410_tag == io_i_addr[12:3] ? btb_410_target_address : _GEN_2046; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2054 = btb_410_tag == io_i_addr[12:3] ? ~btb_410_bht[1] : _GEN_2049; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2055 = btb_411_tag == io_i_addr[12:3] ? btb_411_valid : _GEN_2050; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2056 = btb_411_tag == io_i_addr[12:3] ? btb_411_target_address : _GEN_2051; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2059 = btb_411_tag == io_i_addr[12:3] ? ~btb_411_bht[1] : _GEN_2054; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2060 = btb_412_tag == io_i_addr[12:3] ? btb_412_valid : _GEN_2055; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2061 = btb_412_tag == io_i_addr[12:3] ? btb_412_target_address : _GEN_2056; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2064 = btb_412_tag == io_i_addr[12:3] ? ~btb_412_bht[1] : _GEN_2059; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2065 = btb_413_tag == io_i_addr[12:3] ? btb_413_valid : _GEN_2060; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2066 = btb_413_tag == io_i_addr[12:3] ? btb_413_target_address : _GEN_2061; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2069 = btb_413_tag == io_i_addr[12:3] ? ~btb_413_bht[1] : _GEN_2064; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2070 = btb_414_tag == io_i_addr[12:3] ? btb_414_valid : _GEN_2065; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2071 = btb_414_tag == io_i_addr[12:3] ? btb_414_target_address : _GEN_2066; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2074 = btb_414_tag == io_i_addr[12:3] ? ~btb_414_bht[1] : _GEN_2069; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2075 = btb_415_tag == io_i_addr[12:3] ? btb_415_valid : _GEN_2070; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2076 = btb_415_tag == io_i_addr[12:3] ? btb_415_target_address : _GEN_2071; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2079 = btb_415_tag == io_i_addr[12:3] ? ~btb_415_bht[1] : _GEN_2074; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2080 = btb_416_tag == io_i_addr[12:3] ? btb_416_valid : _GEN_2075; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2081 = btb_416_tag == io_i_addr[12:3] ? btb_416_target_address : _GEN_2076; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2084 = btb_416_tag == io_i_addr[12:3] ? ~btb_416_bht[1] : _GEN_2079; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2085 = btb_417_tag == io_i_addr[12:3] ? btb_417_valid : _GEN_2080; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2086 = btb_417_tag == io_i_addr[12:3] ? btb_417_target_address : _GEN_2081; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2089 = btb_417_tag == io_i_addr[12:3] ? ~btb_417_bht[1] : _GEN_2084; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2090 = btb_418_tag == io_i_addr[12:3] ? btb_418_valid : _GEN_2085; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2091 = btb_418_tag == io_i_addr[12:3] ? btb_418_target_address : _GEN_2086; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2094 = btb_418_tag == io_i_addr[12:3] ? ~btb_418_bht[1] : _GEN_2089; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2095 = btb_419_tag == io_i_addr[12:3] ? btb_419_valid : _GEN_2090; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2096 = btb_419_tag == io_i_addr[12:3] ? btb_419_target_address : _GEN_2091; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2099 = btb_419_tag == io_i_addr[12:3] ? ~btb_419_bht[1] : _GEN_2094; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2100 = btb_420_tag == io_i_addr[12:3] ? btb_420_valid : _GEN_2095; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2101 = btb_420_tag == io_i_addr[12:3] ? btb_420_target_address : _GEN_2096; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2104 = btb_420_tag == io_i_addr[12:3] ? ~btb_420_bht[1] : _GEN_2099; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2105 = btb_421_tag == io_i_addr[12:3] ? btb_421_valid : _GEN_2100; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2106 = btb_421_tag == io_i_addr[12:3] ? btb_421_target_address : _GEN_2101; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2109 = btb_421_tag == io_i_addr[12:3] ? ~btb_421_bht[1] : _GEN_2104; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2110 = btb_422_tag == io_i_addr[12:3] ? btb_422_valid : _GEN_2105; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2111 = btb_422_tag == io_i_addr[12:3] ? btb_422_target_address : _GEN_2106; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2114 = btb_422_tag == io_i_addr[12:3] ? ~btb_422_bht[1] : _GEN_2109; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2115 = btb_423_tag == io_i_addr[12:3] ? btb_423_valid : _GEN_2110; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2116 = btb_423_tag == io_i_addr[12:3] ? btb_423_target_address : _GEN_2111; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2119 = btb_423_tag == io_i_addr[12:3] ? ~btb_423_bht[1] : _GEN_2114; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2120 = btb_424_tag == io_i_addr[12:3] ? btb_424_valid : _GEN_2115; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2121 = btb_424_tag == io_i_addr[12:3] ? btb_424_target_address : _GEN_2116; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2124 = btb_424_tag == io_i_addr[12:3] ? ~btb_424_bht[1] : _GEN_2119; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2125 = btb_425_tag == io_i_addr[12:3] ? btb_425_valid : _GEN_2120; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2126 = btb_425_tag == io_i_addr[12:3] ? btb_425_target_address : _GEN_2121; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2129 = btb_425_tag == io_i_addr[12:3] ? ~btb_425_bht[1] : _GEN_2124; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2130 = btb_426_tag == io_i_addr[12:3] ? btb_426_valid : _GEN_2125; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2131 = btb_426_tag == io_i_addr[12:3] ? btb_426_target_address : _GEN_2126; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2134 = btb_426_tag == io_i_addr[12:3] ? ~btb_426_bht[1] : _GEN_2129; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2135 = btb_427_tag == io_i_addr[12:3] ? btb_427_valid : _GEN_2130; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2136 = btb_427_tag == io_i_addr[12:3] ? btb_427_target_address : _GEN_2131; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2139 = btb_427_tag == io_i_addr[12:3] ? ~btb_427_bht[1] : _GEN_2134; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2140 = btb_428_tag == io_i_addr[12:3] ? btb_428_valid : _GEN_2135; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2141 = btb_428_tag == io_i_addr[12:3] ? btb_428_target_address : _GEN_2136; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2144 = btb_428_tag == io_i_addr[12:3] ? ~btb_428_bht[1] : _GEN_2139; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2145 = btb_429_tag == io_i_addr[12:3] ? btb_429_valid : _GEN_2140; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2146 = btb_429_tag == io_i_addr[12:3] ? btb_429_target_address : _GEN_2141; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2149 = btb_429_tag == io_i_addr[12:3] ? ~btb_429_bht[1] : _GEN_2144; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2150 = btb_430_tag == io_i_addr[12:3] ? btb_430_valid : _GEN_2145; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2151 = btb_430_tag == io_i_addr[12:3] ? btb_430_target_address : _GEN_2146; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2154 = btb_430_tag == io_i_addr[12:3] ? ~btb_430_bht[1] : _GEN_2149; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2155 = btb_431_tag == io_i_addr[12:3] ? btb_431_valid : _GEN_2150; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2156 = btb_431_tag == io_i_addr[12:3] ? btb_431_target_address : _GEN_2151; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2159 = btb_431_tag == io_i_addr[12:3] ? ~btb_431_bht[1] : _GEN_2154; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2160 = btb_432_tag == io_i_addr[12:3] ? btb_432_valid : _GEN_2155; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2161 = btb_432_tag == io_i_addr[12:3] ? btb_432_target_address : _GEN_2156; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2164 = btb_432_tag == io_i_addr[12:3] ? ~btb_432_bht[1] : _GEN_2159; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2165 = btb_433_tag == io_i_addr[12:3] ? btb_433_valid : _GEN_2160; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2166 = btb_433_tag == io_i_addr[12:3] ? btb_433_target_address : _GEN_2161; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2169 = btb_433_tag == io_i_addr[12:3] ? ~btb_433_bht[1] : _GEN_2164; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2170 = btb_434_tag == io_i_addr[12:3] ? btb_434_valid : _GEN_2165; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2171 = btb_434_tag == io_i_addr[12:3] ? btb_434_target_address : _GEN_2166; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2174 = btb_434_tag == io_i_addr[12:3] ? ~btb_434_bht[1] : _GEN_2169; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2175 = btb_435_tag == io_i_addr[12:3] ? btb_435_valid : _GEN_2170; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2176 = btb_435_tag == io_i_addr[12:3] ? btb_435_target_address : _GEN_2171; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2179 = btb_435_tag == io_i_addr[12:3] ? ~btb_435_bht[1] : _GEN_2174; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2180 = btb_436_tag == io_i_addr[12:3] ? btb_436_valid : _GEN_2175; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2181 = btb_436_tag == io_i_addr[12:3] ? btb_436_target_address : _GEN_2176; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2184 = btb_436_tag == io_i_addr[12:3] ? ~btb_436_bht[1] : _GEN_2179; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2185 = btb_437_tag == io_i_addr[12:3] ? btb_437_valid : _GEN_2180; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2186 = btb_437_tag == io_i_addr[12:3] ? btb_437_target_address : _GEN_2181; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2189 = btb_437_tag == io_i_addr[12:3] ? ~btb_437_bht[1] : _GEN_2184; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2190 = btb_438_tag == io_i_addr[12:3] ? btb_438_valid : _GEN_2185; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2191 = btb_438_tag == io_i_addr[12:3] ? btb_438_target_address : _GEN_2186; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2194 = btb_438_tag == io_i_addr[12:3] ? ~btb_438_bht[1] : _GEN_2189; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2195 = btb_439_tag == io_i_addr[12:3] ? btb_439_valid : _GEN_2190; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2196 = btb_439_tag == io_i_addr[12:3] ? btb_439_target_address : _GEN_2191; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2199 = btb_439_tag == io_i_addr[12:3] ? ~btb_439_bht[1] : _GEN_2194; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2200 = btb_440_tag == io_i_addr[12:3] ? btb_440_valid : _GEN_2195; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2201 = btb_440_tag == io_i_addr[12:3] ? btb_440_target_address : _GEN_2196; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2204 = btb_440_tag == io_i_addr[12:3] ? ~btb_440_bht[1] : _GEN_2199; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2205 = btb_441_tag == io_i_addr[12:3] ? btb_441_valid : _GEN_2200; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2206 = btb_441_tag == io_i_addr[12:3] ? btb_441_target_address : _GEN_2201; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2209 = btb_441_tag == io_i_addr[12:3] ? ~btb_441_bht[1] : _GEN_2204; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2210 = btb_442_tag == io_i_addr[12:3] ? btb_442_valid : _GEN_2205; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2211 = btb_442_tag == io_i_addr[12:3] ? btb_442_target_address : _GEN_2206; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2214 = btb_442_tag == io_i_addr[12:3] ? ~btb_442_bht[1] : _GEN_2209; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2215 = btb_443_tag == io_i_addr[12:3] ? btb_443_valid : _GEN_2210; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2216 = btb_443_tag == io_i_addr[12:3] ? btb_443_target_address : _GEN_2211; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2219 = btb_443_tag == io_i_addr[12:3] ? ~btb_443_bht[1] : _GEN_2214; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2220 = btb_444_tag == io_i_addr[12:3] ? btb_444_valid : _GEN_2215; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2221 = btb_444_tag == io_i_addr[12:3] ? btb_444_target_address : _GEN_2216; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2224 = btb_444_tag == io_i_addr[12:3] ? ~btb_444_bht[1] : _GEN_2219; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2225 = btb_445_tag == io_i_addr[12:3] ? btb_445_valid : _GEN_2220; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2226 = btb_445_tag == io_i_addr[12:3] ? btb_445_target_address : _GEN_2221; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2229 = btb_445_tag == io_i_addr[12:3] ? ~btb_445_bht[1] : _GEN_2224; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2230 = btb_446_tag == io_i_addr[12:3] ? btb_446_valid : _GEN_2225; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2231 = btb_446_tag == io_i_addr[12:3] ? btb_446_target_address : _GEN_2226; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2234 = btb_446_tag == io_i_addr[12:3] ? ~btb_446_bht[1] : _GEN_2229; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2235 = btb_447_tag == io_i_addr[12:3] ? btb_447_valid : _GEN_2230; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2236 = btb_447_tag == io_i_addr[12:3] ? btb_447_target_address : _GEN_2231; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2239 = btb_447_tag == io_i_addr[12:3] ? ~btb_447_bht[1] : _GEN_2234; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2240 = btb_448_tag == io_i_addr[12:3] ? btb_448_valid : _GEN_2235; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2241 = btb_448_tag == io_i_addr[12:3] ? btb_448_target_address : _GEN_2236; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2244 = btb_448_tag == io_i_addr[12:3] ? ~btb_448_bht[1] : _GEN_2239; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2245 = btb_449_tag == io_i_addr[12:3] ? btb_449_valid : _GEN_2240; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2246 = btb_449_tag == io_i_addr[12:3] ? btb_449_target_address : _GEN_2241; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2249 = btb_449_tag == io_i_addr[12:3] ? ~btb_449_bht[1] : _GEN_2244; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2250 = btb_450_tag == io_i_addr[12:3] ? btb_450_valid : _GEN_2245; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2251 = btb_450_tag == io_i_addr[12:3] ? btb_450_target_address : _GEN_2246; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2254 = btb_450_tag == io_i_addr[12:3] ? ~btb_450_bht[1] : _GEN_2249; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2255 = btb_451_tag == io_i_addr[12:3] ? btb_451_valid : _GEN_2250; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2256 = btb_451_tag == io_i_addr[12:3] ? btb_451_target_address : _GEN_2251; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2259 = btb_451_tag == io_i_addr[12:3] ? ~btb_451_bht[1] : _GEN_2254; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2260 = btb_452_tag == io_i_addr[12:3] ? btb_452_valid : _GEN_2255; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2261 = btb_452_tag == io_i_addr[12:3] ? btb_452_target_address : _GEN_2256; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2264 = btb_452_tag == io_i_addr[12:3] ? ~btb_452_bht[1] : _GEN_2259; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2265 = btb_453_tag == io_i_addr[12:3] ? btb_453_valid : _GEN_2260; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2266 = btb_453_tag == io_i_addr[12:3] ? btb_453_target_address : _GEN_2261; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2269 = btb_453_tag == io_i_addr[12:3] ? ~btb_453_bht[1] : _GEN_2264; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2270 = btb_454_tag == io_i_addr[12:3] ? btb_454_valid : _GEN_2265; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2271 = btb_454_tag == io_i_addr[12:3] ? btb_454_target_address : _GEN_2266; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2274 = btb_454_tag == io_i_addr[12:3] ? ~btb_454_bht[1] : _GEN_2269; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2275 = btb_455_tag == io_i_addr[12:3] ? btb_455_valid : _GEN_2270; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2276 = btb_455_tag == io_i_addr[12:3] ? btb_455_target_address : _GEN_2271; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2279 = btb_455_tag == io_i_addr[12:3] ? ~btb_455_bht[1] : _GEN_2274; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2280 = btb_456_tag == io_i_addr[12:3] ? btb_456_valid : _GEN_2275; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2281 = btb_456_tag == io_i_addr[12:3] ? btb_456_target_address : _GEN_2276; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2284 = btb_456_tag == io_i_addr[12:3] ? ~btb_456_bht[1] : _GEN_2279; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2285 = btb_457_tag == io_i_addr[12:3] ? btb_457_valid : _GEN_2280; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2286 = btb_457_tag == io_i_addr[12:3] ? btb_457_target_address : _GEN_2281; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2289 = btb_457_tag == io_i_addr[12:3] ? ~btb_457_bht[1] : _GEN_2284; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2290 = btb_458_tag == io_i_addr[12:3] ? btb_458_valid : _GEN_2285; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2291 = btb_458_tag == io_i_addr[12:3] ? btb_458_target_address : _GEN_2286; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2294 = btb_458_tag == io_i_addr[12:3] ? ~btb_458_bht[1] : _GEN_2289; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2295 = btb_459_tag == io_i_addr[12:3] ? btb_459_valid : _GEN_2290; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2296 = btb_459_tag == io_i_addr[12:3] ? btb_459_target_address : _GEN_2291; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2299 = btb_459_tag == io_i_addr[12:3] ? ~btb_459_bht[1] : _GEN_2294; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2300 = btb_460_tag == io_i_addr[12:3] ? btb_460_valid : _GEN_2295; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2301 = btb_460_tag == io_i_addr[12:3] ? btb_460_target_address : _GEN_2296; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2304 = btb_460_tag == io_i_addr[12:3] ? ~btb_460_bht[1] : _GEN_2299; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2305 = btb_461_tag == io_i_addr[12:3] ? btb_461_valid : _GEN_2300; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2306 = btb_461_tag == io_i_addr[12:3] ? btb_461_target_address : _GEN_2301; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2309 = btb_461_tag == io_i_addr[12:3] ? ~btb_461_bht[1] : _GEN_2304; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2310 = btb_462_tag == io_i_addr[12:3] ? btb_462_valid : _GEN_2305; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2311 = btb_462_tag == io_i_addr[12:3] ? btb_462_target_address : _GEN_2306; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2314 = btb_462_tag == io_i_addr[12:3] ? ~btb_462_bht[1] : _GEN_2309; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2315 = btb_463_tag == io_i_addr[12:3] ? btb_463_valid : _GEN_2310; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2316 = btb_463_tag == io_i_addr[12:3] ? btb_463_target_address : _GEN_2311; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2319 = btb_463_tag == io_i_addr[12:3] ? ~btb_463_bht[1] : _GEN_2314; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2320 = btb_464_tag == io_i_addr[12:3] ? btb_464_valid : _GEN_2315; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2321 = btb_464_tag == io_i_addr[12:3] ? btb_464_target_address : _GEN_2316; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2324 = btb_464_tag == io_i_addr[12:3] ? ~btb_464_bht[1] : _GEN_2319; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2325 = btb_465_tag == io_i_addr[12:3] ? btb_465_valid : _GEN_2320; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2326 = btb_465_tag == io_i_addr[12:3] ? btb_465_target_address : _GEN_2321; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2329 = btb_465_tag == io_i_addr[12:3] ? ~btb_465_bht[1] : _GEN_2324; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2330 = btb_466_tag == io_i_addr[12:3] ? btb_466_valid : _GEN_2325; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2331 = btb_466_tag == io_i_addr[12:3] ? btb_466_target_address : _GEN_2326; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2334 = btb_466_tag == io_i_addr[12:3] ? ~btb_466_bht[1] : _GEN_2329; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2335 = btb_467_tag == io_i_addr[12:3] ? btb_467_valid : _GEN_2330; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2336 = btb_467_tag == io_i_addr[12:3] ? btb_467_target_address : _GEN_2331; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2339 = btb_467_tag == io_i_addr[12:3] ? ~btb_467_bht[1] : _GEN_2334; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2340 = btb_468_tag == io_i_addr[12:3] ? btb_468_valid : _GEN_2335; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2341 = btb_468_tag == io_i_addr[12:3] ? btb_468_target_address : _GEN_2336; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2344 = btb_468_tag == io_i_addr[12:3] ? ~btb_468_bht[1] : _GEN_2339; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2345 = btb_469_tag == io_i_addr[12:3] ? btb_469_valid : _GEN_2340; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2346 = btb_469_tag == io_i_addr[12:3] ? btb_469_target_address : _GEN_2341; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2349 = btb_469_tag == io_i_addr[12:3] ? ~btb_469_bht[1] : _GEN_2344; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2350 = btb_470_tag == io_i_addr[12:3] ? btb_470_valid : _GEN_2345; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2351 = btb_470_tag == io_i_addr[12:3] ? btb_470_target_address : _GEN_2346; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2354 = btb_470_tag == io_i_addr[12:3] ? ~btb_470_bht[1] : _GEN_2349; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2355 = btb_471_tag == io_i_addr[12:3] ? btb_471_valid : _GEN_2350; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2356 = btb_471_tag == io_i_addr[12:3] ? btb_471_target_address : _GEN_2351; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2359 = btb_471_tag == io_i_addr[12:3] ? ~btb_471_bht[1] : _GEN_2354; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2360 = btb_472_tag == io_i_addr[12:3] ? btb_472_valid : _GEN_2355; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2361 = btb_472_tag == io_i_addr[12:3] ? btb_472_target_address : _GEN_2356; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2364 = btb_472_tag == io_i_addr[12:3] ? ~btb_472_bht[1] : _GEN_2359; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2365 = btb_473_tag == io_i_addr[12:3] ? btb_473_valid : _GEN_2360; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2366 = btb_473_tag == io_i_addr[12:3] ? btb_473_target_address : _GEN_2361; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2369 = btb_473_tag == io_i_addr[12:3] ? ~btb_473_bht[1] : _GEN_2364; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2370 = btb_474_tag == io_i_addr[12:3] ? btb_474_valid : _GEN_2365; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2371 = btb_474_tag == io_i_addr[12:3] ? btb_474_target_address : _GEN_2366; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2374 = btb_474_tag == io_i_addr[12:3] ? ~btb_474_bht[1] : _GEN_2369; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2375 = btb_475_tag == io_i_addr[12:3] ? btb_475_valid : _GEN_2370; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2376 = btb_475_tag == io_i_addr[12:3] ? btb_475_target_address : _GEN_2371; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2379 = btb_475_tag == io_i_addr[12:3] ? ~btb_475_bht[1] : _GEN_2374; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2380 = btb_476_tag == io_i_addr[12:3] ? btb_476_valid : _GEN_2375; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2381 = btb_476_tag == io_i_addr[12:3] ? btb_476_target_address : _GEN_2376; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2384 = btb_476_tag == io_i_addr[12:3] ? ~btb_476_bht[1] : _GEN_2379; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2385 = btb_477_tag == io_i_addr[12:3] ? btb_477_valid : _GEN_2380; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2386 = btb_477_tag == io_i_addr[12:3] ? btb_477_target_address : _GEN_2381; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2389 = btb_477_tag == io_i_addr[12:3] ? ~btb_477_bht[1] : _GEN_2384; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2390 = btb_478_tag == io_i_addr[12:3] ? btb_478_valid : _GEN_2385; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2391 = btb_478_tag == io_i_addr[12:3] ? btb_478_target_address : _GEN_2386; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2394 = btb_478_tag == io_i_addr[12:3] ? ~btb_478_bht[1] : _GEN_2389; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2395 = btb_479_tag == io_i_addr[12:3] ? btb_479_valid : _GEN_2390; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2396 = btb_479_tag == io_i_addr[12:3] ? btb_479_target_address : _GEN_2391; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2399 = btb_479_tag == io_i_addr[12:3] ? ~btb_479_bht[1] : _GEN_2394; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2400 = btb_480_tag == io_i_addr[12:3] ? btb_480_valid : _GEN_2395; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2401 = btb_480_tag == io_i_addr[12:3] ? btb_480_target_address : _GEN_2396; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2404 = btb_480_tag == io_i_addr[12:3] ? ~btb_480_bht[1] : _GEN_2399; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2405 = btb_481_tag == io_i_addr[12:3] ? btb_481_valid : _GEN_2400; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2406 = btb_481_tag == io_i_addr[12:3] ? btb_481_target_address : _GEN_2401; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2409 = btb_481_tag == io_i_addr[12:3] ? ~btb_481_bht[1] : _GEN_2404; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2410 = btb_482_tag == io_i_addr[12:3] ? btb_482_valid : _GEN_2405; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2411 = btb_482_tag == io_i_addr[12:3] ? btb_482_target_address : _GEN_2406; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2414 = btb_482_tag == io_i_addr[12:3] ? ~btb_482_bht[1] : _GEN_2409; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2415 = btb_483_tag == io_i_addr[12:3] ? btb_483_valid : _GEN_2410; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2416 = btb_483_tag == io_i_addr[12:3] ? btb_483_target_address : _GEN_2411; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2419 = btb_483_tag == io_i_addr[12:3] ? ~btb_483_bht[1] : _GEN_2414; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2420 = btb_484_tag == io_i_addr[12:3] ? btb_484_valid : _GEN_2415; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2421 = btb_484_tag == io_i_addr[12:3] ? btb_484_target_address : _GEN_2416; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2424 = btb_484_tag == io_i_addr[12:3] ? ~btb_484_bht[1] : _GEN_2419; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2425 = btb_485_tag == io_i_addr[12:3] ? btb_485_valid : _GEN_2420; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2426 = btb_485_tag == io_i_addr[12:3] ? btb_485_target_address : _GEN_2421; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2429 = btb_485_tag == io_i_addr[12:3] ? ~btb_485_bht[1] : _GEN_2424; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2430 = btb_486_tag == io_i_addr[12:3] ? btb_486_valid : _GEN_2425; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2431 = btb_486_tag == io_i_addr[12:3] ? btb_486_target_address : _GEN_2426; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2434 = btb_486_tag == io_i_addr[12:3] ? ~btb_486_bht[1] : _GEN_2429; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2435 = btb_487_tag == io_i_addr[12:3] ? btb_487_valid : _GEN_2430; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2436 = btb_487_tag == io_i_addr[12:3] ? btb_487_target_address : _GEN_2431; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2439 = btb_487_tag == io_i_addr[12:3] ? ~btb_487_bht[1] : _GEN_2434; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2440 = btb_488_tag == io_i_addr[12:3] ? btb_488_valid : _GEN_2435; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2441 = btb_488_tag == io_i_addr[12:3] ? btb_488_target_address : _GEN_2436; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2444 = btb_488_tag == io_i_addr[12:3] ? ~btb_488_bht[1] : _GEN_2439; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2445 = btb_489_tag == io_i_addr[12:3] ? btb_489_valid : _GEN_2440; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2446 = btb_489_tag == io_i_addr[12:3] ? btb_489_target_address : _GEN_2441; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2449 = btb_489_tag == io_i_addr[12:3] ? ~btb_489_bht[1] : _GEN_2444; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2450 = btb_490_tag == io_i_addr[12:3] ? btb_490_valid : _GEN_2445; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2451 = btb_490_tag == io_i_addr[12:3] ? btb_490_target_address : _GEN_2446; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2454 = btb_490_tag == io_i_addr[12:3] ? ~btb_490_bht[1] : _GEN_2449; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2455 = btb_491_tag == io_i_addr[12:3] ? btb_491_valid : _GEN_2450; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2456 = btb_491_tag == io_i_addr[12:3] ? btb_491_target_address : _GEN_2451; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2459 = btb_491_tag == io_i_addr[12:3] ? ~btb_491_bht[1] : _GEN_2454; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2460 = btb_492_tag == io_i_addr[12:3] ? btb_492_valid : _GEN_2455; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2461 = btb_492_tag == io_i_addr[12:3] ? btb_492_target_address : _GEN_2456; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2464 = btb_492_tag == io_i_addr[12:3] ? ~btb_492_bht[1] : _GEN_2459; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2465 = btb_493_tag == io_i_addr[12:3] ? btb_493_valid : _GEN_2460; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2466 = btb_493_tag == io_i_addr[12:3] ? btb_493_target_address : _GEN_2461; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2469 = btb_493_tag == io_i_addr[12:3] ? ~btb_493_bht[1] : _GEN_2464; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2470 = btb_494_tag == io_i_addr[12:3] ? btb_494_valid : _GEN_2465; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2471 = btb_494_tag == io_i_addr[12:3] ? btb_494_target_address : _GEN_2466; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2474 = btb_494_tag == io_i_addr[12:3] ? ~btb_494_bht[1] : _GEN_2469; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2475 = btb_495_tag == io_i_addr[12:3] ? btb_495_valid : _GEN_2470; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2476 = btb_495_tag == io_i_addr[12:3] ? btb_495_target_address : _GEN_2471; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2479 = btb_495_tag == io_i_addr[12:3] ? ~btb_495_bht[1] : _GEN_2474; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2480 = btb_496_tag == io_i_addr[12:3] ? btb_496_valid : _GEN_2475; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2481 = btb_496_tag == io_i_addr[12:3] ? btb_496_target_address : _GEN_2476; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2484 = btb_496_tag == io_i_addr[12:3] ? ~btb_496_bht[1] : _GEN_2479; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2485 = btb_497_tag == io_i_addr[12:3] ? btb_497_valid : _GEN_2480; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2486 = btb_497_tag == io_i_addr[12:3] ? btb_497_target_address : _GEN_2481; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2489 = btb_497_tag == io_i_addr[12:3] ? ~btb_497_bht[1] : _GEN_2484; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2490 = btb_498_tag == io_i_addr[12:3] ? btb_498_valid : _GEN_2485; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2491 = btb_498_tag == io_i_addr[12:3] ? btb_498_target_address : _GEN_2486; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2494 = btb_498_tag == io_i_addr[12:3] ? ~btb_498_bht[1] : _GEN_2489; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2495 = btb_499_tag == io_i_addr[12:3] ? btb_499_valid : _GEN_2490; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2496 = btb_499_tag == io_i_addr[12:3] ? btb_499_target_address : _GEN_2491; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2499 = btb_499_tag == io_i_addr[12:3] ? ~btb_499_bht[1] : _GEN_2494; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2500 = btb_500_tag == io_i_addr[12:3] ? btb_500_valid : _GEN_2495; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2501 = btb_500_tag == io_i_addr[12:3] ? btb_500_target_address : _GEN_2496; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2504 = btb_500_tag == io_i_addr[12:3] ? ~btb_500_bht[1] : _GEN_2499; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2505 = btb_501_tag == io_i_addr[12:3] ? btb_501_valid : _GEN_2500; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2506 = btb_501_tag == io_i_addr[12:3] ? btb_501_target_address : _GEN_2501; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2509 = btb_501_tag == io_i_addr[12:3] ? ~btb_501_bht[1] : _GEN_2504; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2510 = btb_502_tag == io_i_addr[12:3] ? btb_502_valid : _GEN_2505; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2511 = btb_502_tag == io_i_addr[12:3] ? btb_502_target_address : _GEN_2506; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2514 = btb_502_tag == io_i_addr[12:3] ? ~btb_502_bht[1] : _GEN_2509; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2515 = btb_503_tag == io_i_addr[12:3] ? btb_503_valid : _GEN_2510; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2516 = btb_503_tag == io_i_addr[12:3] ? btb_503_target_address : _GEN_2511; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2519 = btb_503_tag == io_i_addr[12:3] ? ~btb_503_bht[1] : _GEN_2514; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2520 = btb_504_tag == io_i_addr[12:3] ? btb_504_valid : _GEN_2515; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2521 = btb_504_tag == io_i_addr[12:3] ? btb_504_target_address : _GEN_2516; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2524 = btb_504_tag == io_i_addr[12:3] ? ~btb_504_bht[1] : _GEN_2519; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2525 = btb_505_tag == io_i_addr[12:3] ? btb_505_valid : _GEN_2520; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2526 = btb_505_tag == io_i_addr[12:3] ? btb_505_target_address : _GEN_2521; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2529 = btb_505_tag == io_i_addr[12:3] ? ~btb_505_bht[1] : _GEN_2524; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2530 = btb_506_tag == io_i_addr[12:3] ? btb_506_valid : _GEN_2525; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2531 = btb_506_tag == io_i_addr[12:3] ? btb_506_target_address : _GEN_2526; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2534 = btb_506_tag == io_i_addr[12:3] ? ~btb_506_bht[1] : _GEN_2529; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2535 = btb_507_tag == io_i_addr[12:3] ? btb_507_valid : _GEN_2530; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2536 = btb_507_tag == io_i_addr[12:3] ? btb_507_target_address : _GEN_2531; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2539 = btb_507_tag == io_i_addr[12:3] ? ~btb_507_bht[1] : _GEN_2534; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2540 = btb_508_tag == io_i_addr[12:3] ? btb_508_valid : _GEN_2535; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2541 = btb_508_tag == io_i_addr[12:3] ? btb_508_target_address : _GEN_2536; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2544 = btb_508_tag == io_i_addr[12:3] ? ~btb_508_bht[1] : _GEN_2539; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2545 = btb_509_tag == io_i_addr[12:3] ? btb_509_valid : _GEN_2540; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2546 = btb_509_tag == io_i_addr[12:3] ? btb_509_target_address : _GEN_2541; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2549 = btb_509_tag == io_i_addr[12:3] ? ~btb_509_bht[1] : _GEN_2544; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_2550 = btb_510_tag == io_i_addr[12:3] ? btb_510_valid : _GEN_2545; // @[branch_predictor.scala 40:45 41:44]
  wire [63:0] _GEN_2551 = btb_510_tag == io_i_addr[12:3] ? btb_510_target_address : _GEN_2546; // @[branch_predictor.scala 40:45 42:45]
  wire  _GEN_2554 = btb_510_tag == io_i_addr[12:3] ? ~btb_510_bht[1] : _GEN_2549; // @[branch_predictor.scala 40:45 45:44]
  wire  _GEN_19459 = 9'h0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2560 = 9'h0 == btb_victim_ptr | btb_0_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19460 = 9'h1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2561 = 9'h1 == btb_victim_ptr | btb_1_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19461 = 9'h2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2562 = 9'h2 == btb_victim_ptr | btb_2_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19462 = 9'h3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2563 = 9'h3 == btb_victim_ptr | btb_3_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19463 = 9'h4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2564 = 9'h4 == btb_victim_ptr | btb_4_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19464 = 9'h5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2565 = 9'h5 == btb_victim_ptr | btb_5_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19465 = 9'h6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2566 = 9'h6 == btb_victim_ptr | btb_6_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19466 = 9'h7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2567 = 9'h7 == btb_victim_ptr | btb_7_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19467 = 9'h8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2568 = 9'h8 == btb_victim_ptr | btb_8_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19468 = 9'h9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2569 = 9'h9 == btb_victim_ptr | btb_9_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19469 = 9'ha == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2570 = 9'ha == btb_victim_ptr | btb_10_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19470 = 9'hb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2571 = 9'hb == btb_victim_ptr | btb_11_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19471 = 9'hc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2572 = 9'hc == btb_victim_ptr | btb_12_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19472 = 9'hd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2573 = 9'hd == btb_victim_ptr | btb_13_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19473 = 9'he == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2574 = 9'he == btb_victim_ptr | btb_14_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19474 = 9'hf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2575 = 9'hf == btb_victim_ptr | btb_15_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19475 = 9'h10 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2576 = 9'h10 == btb_victim_ptr | btb_16_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19476 = 9'h11 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2577 = 9'h11 == btb_victim_ptr | btb_17_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19477 = 9'h12 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2578 = 9'h12 == btb_victim_ptr | btb_18_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19478 = 9'h13 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2579 = 9'h13 == btb_victim_ptr | btb_19_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19479 = 9'h14 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2580 = 9'h14 == btb_victim_ptr | btb_20_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19480 = 9'h15 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2581 = 9'h15 == btb_victim_ptr | btb_21_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19481 = 9'h16 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2582 = 9'h16 == btb_victim_ptr | btb_22_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19482 = 9'h17 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2583 = 9'h17 == btb_victim_ptr | btb_23_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19483 = 9'h18 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2584 = 9'h18 == btb_victim_ptr | btb_24_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19484 = 9'h19 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2585 = 9'h19 == btb_victim_ptr | btb_25_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19485 = 9'h1a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2586 = 9'h1a == btb_victim_ptr | btb_26_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19486 = 9'h1b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2587 = 9'h1b == btb_victim_ptr | btb_27_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19487 = 9'h1c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2588 = 9'h1c == btb_victim_ptr | btb_28_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19488 = 9'h1d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2589 = 9'h1d == btb_victim_ptr | btb_29_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19489 = 9'h1e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2590 = 9'h1e == btb_victim_ptr | btb_30_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19490 = 9'h1f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2591 = 9'h1f == btb_victim_ptr | btb_31_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19491 = 9'h20 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2592 = 9'h20 == btb_victim_ptr | btb_32_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19492 = 9'h21 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2593 = 9'h21 == btb_victim_ptr | btb_33_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19493 = 9'h22 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2594 = 9'h22 == btb_victim_ptr | btb_34_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19494 = 9'h23 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2595 = 9'h23 == btb_victim_ptr | btb_35_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19495 = 9'h24 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2596 = 9'h24 == btb_victim_ptr | btb_36_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19496 = 9'h25 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2597 = 9'h25 == btb_victim_ptr | btb_37_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19497 = 9'h26 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2598 = 9'h26 == btb_victim_ptr | btb_38_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19498 = 9'h27 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2599 = 9'h27 == btb_victim_ptr | btb_39_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19499 = 9'h28 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2600 = 9'h28 == btb_victim_ptr | btb_40_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19500 = 9'h29 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2601 = 9'h29 == btb_victim_ptr | btb_41_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19501 = 9'h2a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2602 = 9'h2a == btb_victim_ptr | btb_42_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19502 = 9'h2b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2603 = 9'h2b == btb_victim_ptr | btb_43_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19503 = 9'h2c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2604 = 9'h2c == btb_victim_ptr | btb_44_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19504 = 9'h2d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2605 = 9'h2d == btb_victim_ptr | btb_45_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19505 = 9'h2e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2606 = 9'h2e == btb_victim_ptr | btb_46_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19506 = 9'h2f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2607 = 9'h2f == btb_victim_ptr | btb_47_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19507 = 9'h30 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2608 = 9'h30 == btb_victim_ptr | btb_48_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19508 = 9'h31 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2609 = 9'h31 == btb_victim_ptr | btb_49_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19509 = 9'h32 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2610 = 9'h32 == btb_victim_ptr | btb_50_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19510 = 9'h33 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2611 = 9'h33 == btb_victim_ptr | btb_51_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19511 = 9'h34 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2612 = 9'h34 == btb_victim_ptr | btb_52_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19512 = 9'h35 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2613 = 9'h35 == btb_victim_ptr | btb_53_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19513 = 9'h36 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2614 = 9'h36 == btb_victim_ptr | btb_54_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19514 = 9'h37 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2615 = 9'h37 == btb_victim_ptr | btb_55_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19515 = 9'h38 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2616 = 9'h38 == btb_victim_ptr | btb_56_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19516 = 9'h39 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2617 = 9'h39 == btb_victim_ptr | btb_57_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19517 = 9'h3a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2618 = 9'h3a == btb_victim_ptr | btb_58_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19518 = 9'h3b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2619 = 9'h3b == btb_victim_ptr | btb_59_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19519 = 9'h3c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2620 = 9'h3c == btb_victim_ptr | btb_60_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19520 = 9'h3d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2621 = 9'h3d == btb_victim_ptr | btb_61_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19521 = 9'h3e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2622 = 9'h3e == btb_victim_ptr | btb_62_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19522 = 9'h3f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2623 = 9'h3f == btb_victim_ptr | btb_63_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19523 = 9'h40 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2624 = 9'h40 == btb_victim_ptr | btb_64_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19524 = 9'h41 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2625 = 9'h41 == btb_victim_ptr | btb_65_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19525 = 9'h42 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2626 = 9'h42 == btb_victim_ptr | btb_66_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19526 = 9'h43 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2627 = 9'h43 == btb_victim_ptr | btb_67_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19527 = 9'h44 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2628 = 9'h44 == btb_victim_ptr | btb_68_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19528 = 9'h45 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2629 = 9'h45 == btb_victim_ptr | btb_69_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19529 = 9'h46 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2630 = 9'h46 == btb_victim_ptr | btb_70_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19530 = 9'h47 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2631 = 9'h47 == btb_victim_ptr | btb_71_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19531 = 9'h48 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2632 = 9'h48 == btb_victim_ptr | btb_72_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19532 = 9'h49 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2633 = 9'h49 == btb_victim_ptr | btb_73_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19533 = 9'h4a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2634 = 9'h4a == btb_victim_ptr | btb_74_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19534 = 9'h4b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2635 = 9'h4b == btb_victim_ptr | btb_75_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19535 = 9'h4c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2636 = 9'h4c == btb_victim_ptr | btb_76_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19536 = 9'h4d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2637 = 9'h4d == btb_victim_ptr | btb_77_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19537 = 9'h4e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2638 = 9'h4e == btb_victim_ptr | btb_78_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19538 = 9'h4f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2639 = 9'h4f == btb_victim_ptr | btb_79_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19539 = 9'h50 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2640 = 9'h50 == btb_victim_ptr | btb_80_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19540 = 9'h51 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2641 = 9'h51 == btb_victim_ptr | btb_81_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19541 = 9'h52 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2642 = 9'h52 == btb_victim_ptr | btb_82_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19542 = 9'h53 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2643 = 9'h53 == btb_victim_ptr | btb_83_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19543 = 9'h54 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2644 = 9'h54 == btb_victim_ptr | btb_84_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19544 = 9'h55 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2645 = 9'h55 == btb_victim_ptr | btb_85_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19545 = 9'h56 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2646 = 9'h56 == btb_victim_ptr | btb_86_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19546 = 9'h57 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2647 = 9'h57 == btb_victim_ptr | btb_87_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19547 = 9'h58 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2648 = 9'h58 == btb_victim_ptr | btb_88_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19548 = 9'h59 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2649 = 9'h59 == btb_victim_ptr | btb_89_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19549 = 9'h5a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2650 = 9'h5a == btb_victim_ptr | btb_90_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19550 = 9'h5b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2651 = 9'h5b == btb_victim_ptr | btb_91_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19551 = 9'h5c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2652 = 9'h5c == btb_victim_ptr | btb_92_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19552 = 9'h5d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2653 = 9'h5d == btb_victim_ptr | btb_93_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19553 = 9'h5e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2654 = 9'h5e == btb_victim_ptr | btb_94_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19554 = 9'h5f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2655 = 9'h5f == btb_victim_ptr | btb_95_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19555 = 9'h60 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2656 = 9'h60 == btb_victim_ptr | btb_96_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19556 = 9'h61 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2657 = 9'h61 == btb_victim_ptr | btb_97_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19557 = 9'h62 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2658 = 9'h62 == btb_victim_ptr | btb_98_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19558 = 9'h63 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2659 = 9'h63 == btb_victim_ptr | btb_99_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19559 = 9'h64 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2660 = 9'h64 == btb_victim_ptr | btb_100_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19560 = 9'h65 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2661 = 9'h65 == btb_victim_ptr | btb_101_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19561 = 9'h66 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2662 = 9'h66 == btb_victim_ptr | btb_102_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19562 = 9'h67 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2663 = 9'h67 == btb_victim_ptr | btb_103_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19563 = 9'h68 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2664 = 9'h68 == btb_victim_ptr | btb_104_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19564 = 9'h69 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2665 = 9'h69 == btb_victim_ptr | btb_105_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19565 = 9'h6a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2666 = 9'h6a == btb_victim_ptr | btb_106_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19566 = 9'h6b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2667 = 9'h6b == btb_victim_ptr | btb_107_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19567 = 9'h6c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2668 = 9'h6c == btb_victim_ptr | btb_108_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19568 = 9'h6d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2669 = 9'h6d == btb_victim_ptr | btb_109_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19569 = 9'h6e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2670 = 9'h6e == btb_victim_ptr | btb_110_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19570 = 9'h6f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2671 = 9'h6f == btb_victim_ptr | btb_111_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19571 = 9'h70 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2672 = 9'h70 == btb_victim_ptr | btb_112_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19572 = 9'h71 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2673 = 9'h71 == btb_victim_ptr | btb_113_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19573 = 9'h72 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2674 = 9'h72 == btb_victim_ptr | btb_114_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19574 = 9'h73 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2675 = 9'h73 == btb_victim_ptr | btb_115_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19575 = 9'h74 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2676 = 9'h74 == btb_victim_ptr | btb_116_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19576 = 9'h75 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2677 = 9'h75 == btb_victim_ptr | btb_117_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19577 = 9'h76 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2678 = 9'h76 == btb_victim_ptr | btb_118_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19578 = 9'h77 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2679 = 9'h77 == btb_victim_ptr | btb_119_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19579 = 9'h78 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2680 = 9'h78 == btb_victim_ptr | btb_120_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19580 = 9'h79 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2681 = 9'h79 == btb_victim_ptr | btb_121_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19581 = 9'h7a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2682 = 9'h7a == btb_victim_ptr | btb_122_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19582 = 9'h7b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2683 = 9'h7b == btb_victim_ptr | btb_123_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19583 = 9'h7c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2684 = 9'h7c == btb_victim_ptr | btb_124_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19584 = 9'h7d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2685 = 9'h7d == btb_victim_ptr | btb_125_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19585 = 9'h7e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2686 = 9'h7e == btb_victim_ptr | btb_126_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19586 = 9'h7f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2687 = 9'h7f == btb_victim_ptr | btb_127_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19587 = 9'h80 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2688 = 9'h80 == btb_victim_ptr | btb_128_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19588 = 9'h81 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2689 = 9'h81 == btb_victim_ptr | btb_129_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19589 = 9'h82 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2690 = 9'h82 == btb_victim_ptr | btb_130_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19590 = 9'h83 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2691 = 9'h83 == btb_victim_ptr | btb_131_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19591 = 9'h84 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2692 = 9'h84 == btb_victim_ptr | btb_132_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19592 = 9'h85 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2693 = 9'h85 == btb_victim_ptr | btb_133_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19593 = 9'h86 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2694 = 9'h86 == btb_victim_ptr | btb_134_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19594 = 9'h87 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2695 = 9'h87 == btb_victim_ptr | btb_135_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19595 = 9'h88 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2696 = 9'h88 == btb_victim_ptr | btb_136_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19596 = 9'h89 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2697 = 9'h89 == btb_victim_ptr | btb_137_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19597 = 9'h8a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2698 = 9'h8a == btb_victim_ptr | btb_138_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19598 = 9'h8b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2699 = 9'h8b == btb_victim_ptr | btb_139_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19599 = 9'h8c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2700 = 9'h8c == btb_victim_ptr | btb_140_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19600 = 9'h8d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2701 = 9'h8d == btb_victim_ptr | btb_141_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19601 = 9'h8e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2702 = 9'h8e == btb_victim_ptr | btb_142_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19602 = 9'h8f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2703 = 9'h8f == btb_victim_ptr | btb_143_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19603 = 9'h90 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2704 = 9'h90 == btb_victim_ptr | btb_144_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19604 = 9'h91 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2705 = 9'h91 == btb_victim_ptr | btb_145_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19605 = 9'h92 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2706 = 9'h92 == btb_victim_ptr | btb_146_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19606 = 9'h93 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2707 = 9'h93 == btb_victim_ptr | btb_147_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19607 = 9'h94 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2708 = 9'h94 == btb_victim_ptr | btb_148_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19608 = 9'h95 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2709 = 9'h95 == btb_victim_ptr | btb_149_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19609 = 9'h96 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2710 = 9'h96 == btb_victim_ptr | btb_150_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19610 = 9'h97 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2711 = 9'h97 == btb_victim_ptr | btb_151_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19611 = 9'h98 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2712 = 9'h98 == btb_victim_ptr | btb_152_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19612 = 9'h99 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2713 = 9'h99 == btb_victim_ptr | btb_153_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19613 = 9'h9a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2714 = 9'h9a == btb_victim_ptr | btb_154_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19614 = 9'h9b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2715 = 9'h9b == btb_victim_ptr | btb_155_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19615 = 9'h9c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2716 = 9'h9c == btb_victim_ptr | btb_156_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19616 = 9'h9d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2717 = 9'h9d == btb_victim_ptr | btb_157_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19617 = 9'h9e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2718 = 9'h9e == btb_victim_ptr | btb_158_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19618 = 9'h9f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2719 = 9'h9f == btb_victim_ptr | btb_159_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19619 = 9'ha0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2720 = 9'ha0 == btb_victim_ptr | btb_160_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19620 = 9'ha1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2721 = 9'ha1 == btb_victim_ptr | btb_161_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19621 = 9'ha2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2722 = 9'ha2 == btb_victim_ptr | btb_162_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19622 = 9'ha3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2723 = 9'ha3 == btb_victim_ptr | btb_163_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19623 = 9'ha4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2724 = 9'ha4 == btb_victim_ptr | btb_164_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19624 = 9'ha5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2725 = 9'ha5 == btb_victim_ptr | btb_165_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19625 = 9'ha6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2726 = 9'ha6 == btb_victim_ptr | btb_166_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19626 = 9'ha7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2727 = 9'ha7 == btb_victim_ptr | btb_167_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19627 = 9'ha8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2728 = 9'ha8 == btb_victim_ptr | btb_168_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19628 = 9'ha9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2729 = 9'ha9 == btb_victim_ptr | btb_169_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19629 = 9'haa == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2730 = 9'haa == btb_victim_ptr | btb_170_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19630 = 9'hab == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2731 = 9'hab == btb_victim_ptr | btb_171_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19631 = 9'hac == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2732 = 9'hac == btb_victim_ptr | btb_172_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19632 = 9'had == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2733 = 9'had == btb_victim_ptr | btb_173_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19633 = 9'hae == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2734 = 9'hae == btb_victim_ptr | btb_174_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19634 = 9'haf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2735 = 9'haf == btb_victim_ptr | btb_175_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19635 = 9'hb0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2736 = 9'hb0 == btb_victim_ptr | btb_176_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19636 = 9'hb1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2737 = 9'hb1 == btb_victim_ptr | btb_177_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19637 = 9'hb2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2738 = 9'hb2 == btb_victim_ptr | btb_178_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19638 = 9'hb3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2739 = 9'hb3 == btb_victim_ptr | btb_179_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19639 = 9'hb4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2740 = 9'hb4 == btb_victim_ptr | btb_180_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19640 = 9'hb5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2741 = 9'hb5 == btb_victim_ptr | btb_181_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19641 = 9'hb6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2742 = 9'hb6 == btb_victim_ptr | btb_182_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19642 = 9'hb7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2743 = 9'hb7 == btb_victim_ptr | btb_183_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19643 = 9'hb8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2744 = 9'hb8 == btb_victim_ptr | btb_184_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19644 = 9'hb9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2745 = 9'hb9 == btb_victim_ptr | btb_185_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19645 = 9'hba == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2746 = 9'hba == btb_victim_ptr | btb_186_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19646 = 9'hbb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2747 = 9'hbb == btb_victim_ptr | btb_187_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19647 = 9'hbc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2748 = 9'hbc == btb_victim_ptr | btb_188_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19648 = 9'hbd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2749 = 9'hbd == btb_victim_ptr | btb_189_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19649 = 9'hbe == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2750 = 9'hbe == btb_victim_ptr | btb_190_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19650 = 9'hbf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2751 = 9'hbf == btb_victim_ptr | btb_191_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19651 = 9'hc0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2752 = 9'hc0 == btb_victim_ptr | btb_192_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19652 = 9'hc1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2753 = 9'hc1 == btb_victim_ptr | btb_193_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19653 = 9'hc2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2754 = 9'hc2 == btb_victim_ptr | btb_194_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19654 = 9'hc3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2755 = 9'hc3 == btb_victim_ptr | btb_195_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19655 = 9'hc4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2756 = 9'hc4 == btb_victim_ptr | btb_196_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19656 = 9'hc5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2757 = 9'hc5 == btb_victim_ptr | btb_197_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19657 = 9'hc6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2758 = 9'hc6 == btb_victim_ptr | btb_198_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19658 = 9'hc7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2759 = 9'hc7 == btb_victim_ptr | btb_199_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19659 = 9'hc8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2760 = 9'hc8 == btb_victim_ptr | btb_200_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19660 = 9'hc9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2761 = 9'hc9 == btb_victim_ptr | btb_201_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19661 = 9'hca == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2762 = 9'hca == btb_victim_ptr | btb_202_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19662 = 9'hcb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2763 = 9'hcb == btb_victim_ptr | btb_203_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19663 = 9'hcc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2764 = 9'hcc == btb_victim_ptr | btb_204_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19664 = 9'hcd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2765 = 9'hcd == btb_victim_ptr | btb_205_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19665 = 9'hce == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2766 = 9'hce == btb_victim_ptr | btb_206_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19666 = 9'hcf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2767 = 9'hcf == btb_victim_ptr | btb_207_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19667 = 9'hd0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2768 = 9'hd0 == btb_victim_ptr | btb_208_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19668 = 9'hd1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2769 = 9'hd1 == btb_victim_ptr | btb_209_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19669 = 9'hd2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2770 = 9'hd2 == btb_victim_ptr | btb_210_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19670 = 9'hd3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2771 = 9'hd3 == btb_victim_ptr | btb_211_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19671 = 9'hd4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2772 = 9'hd4 == btb_victim_ptr | btb_212_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19672 = 9'hd5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2773 = 9'hd5 == btb_victim_ptr | btb_213_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19673 = 9'hd6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2774 = 9'hd6 == btb_victim_ptr | btb_214_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19674 = 9'hd7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2775 = 9'hd7 == btb_victim_ptr | btb_215_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19675 = 9'hd8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2776 = 9'hd8 == btb_victim_ptr | btb_216_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19676 = 9'hd9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2777 = 9'hd9 == btb_victim_ptr | btb_217_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19677 = 9'hda == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2778 = 9'hda == btb_victim_ptr | btb_218_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19678 = 9'hdb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2779 = 9'hdb == btb_victim_ptr | btb_219_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19679 = 9'hdc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2780 = 9'hdc == btb_victim_ptr | btb_220_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19680 = 9'hdd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2781 = 9'hdd == btb_victim_ptr | btb_221_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19681 = 9'hde == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2782 = 9'hde == btb_victim_ptr | btb_222_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19682 = 9'hdf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2783 = 9'hdf == btb_victim_ptr | btb_223_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19683 = 9'he0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2784 = 9'he0 == btb_victim_ptr | btb_224_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19684 = 9'he1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2785 = 9'he1 == btb_victim_ptr | btb_225_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19685 = 9'he2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2786 = 9'he2 == btb_victim_ptr | btb_226_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19686 = 9'he3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2787 = 9'he3 == btb_victim_ptr | btb_227_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19687 = 9'he4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2788 = 9'he4 == btb_victim_ptr | btb_228_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19688 = 9'he5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2789 = 9'he5 == btb_victim_ptr | btb_229_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19689 = 9'he6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2790 = 9'he6 == btb_victim_ptr | btb_230_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19690 = 9'he7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2791 = 9'he7 == btb_victim_ptr | btb_231_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19691 = 9'he8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2792 = 9'he8 == btb_victim_ptr | btb_232_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19692 = 9'he9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2793 = 9'he9 == btb_victim_ptr | btb_233_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19693 = 9'hea == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2794 = 9'hea == btb_victim_ptr | btb_234_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19694 = 9'heb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2795 = 9'heb == btb_victim_ptr | btb_235_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19695 = 9'hec == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2796 = 9'hec == btb_victim_ptr | btb_236_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19696 = 9'hed == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2797 = 9'hed == btb_victim_ptr | btb_237_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19697 = 9'hee == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2798 = 9'hee == btb_victim_ptr | btb_238_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19698 = 9'hef == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2799 = 9'hef == btb_victim_ptr | btb_239_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19699 = 9'hf0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2800 = 9'hf0 == btb_victim_ptr | btb_240_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19700 = 9'hf1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2801 = 9'hf1 == btb_victim_ptr | btb_241_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19701 = 9'hf2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2802 = 9'hf2 == btb_victim_ptr | btb_242_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19702 = 9'hf3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2803 = 9'hf3 == btb_victim_ptr | btb_243_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19703 = 9'hf4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2804 = 9'hf4 == btb_victim_ptr | btb_244_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19704 = 9'hf5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2805 = 9'hf5 == btb_victim_ptr | btb_245_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19705 = 9'hf6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2806 = 9'hf6 == btb_victim_ptr | btb_246_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19706 = 9'hf7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2807 = 9'hf7 == btb_victim_ptr | btb_247_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19707 = 9'hf8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2808 = 9'hf8 == btb_victim_ptr | btb_248_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19708 = 9'hf9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2809 = 9'hf9 == btb_victim_ptr | btb_249_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19709 = 9'hfa == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2810 = 9'hfa == btb_victim_ptr | btb_250_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19710 = 9'hfb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2811 = 9'hfb == btb_victim_ptr | btb_251_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19711 = 9'hfc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2812 = 9'hfc == btb_victim_ptr | btb_252_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19712 = 9'hfd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2813 = 9'hfd == btb_victim_ptr | btb_253_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19713 = 9'hfe == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2814 = 9'hfe == btb_victim_ptr | btb_254_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19714 = 9'hff == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2815 = 9'hff == btb_victim_ptr | btb_255_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19715 = 9'h100 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2816 = 9'h100 == btb_victim_ptr | btb_256_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19716 = 9'h101 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2817 = 9'h101 == btb_victim_ptr | btb_257_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19717 = 9'h102 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2818 = 9'h102 == btb_victim_ptr | btb_258_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19718 = 9'h103 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2819 = 9'h103 == btb_victim_ptr | btb_259_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19719 = 9'h104 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2820 = 9'h104 == btb_victim_ptr | btb_260_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19720 = 9'h105 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2821 = 9'h105 == btb_victim_ptr | btb_261_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19721 = 9'h106 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2822 = 9'h106 == btb_victim_ptr | btb_262_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19722 = 9'h107 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2823 = 9'h107 == btb_victim_ptr | btb_263_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19723 = 9'h108 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2824 = 9'h108 == btb_victim_ptr | btb_264_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19724 = 9'h109 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2825 = 9'h109 == btb_victim_ptr | btb_265_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19725 = 9'h10a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2826 = 9'h10a == btb_victim_ptr | btb_266_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19726 = 9'h10b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2827 = 9'h10b == btb_victim_ptr | btb_267_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19727 = 9'h10c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2828 = 9'h10c == btb_victim_ptr | btb_268_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19728 = 9'h10d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2829 = 9'h10d == btb_victim_ptr | btb_269_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19729 = 9'h10e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2830 = 9'h10e == btb_victim_ptr | btb_270_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19730 = 9'h10f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2831 = 9'h10f == btb_victim_ptr | btb_271_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19731 = 9'h110 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2832 = 9'h110 == btb_victim_ptr | btb_272_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19732 = 9'h111 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2833 = 9'h111 == btb_victim_ptr | btb_273_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19733 = 9'h112 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2834 = 9'h112 == btb_victim_ptr | btb_274_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19734 = 9'h113 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2835 = 9'h113 == btb_victim_ptr | btb_275_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19735 = 9'h114 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2836 = 9'h114 == btb_victim_ptr | btb_276_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19736 = 9'h115 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2837 = 9'h115 == btb_victim_ptr | btb_277_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19737 = 9'h116 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2838 = 9'h116 == btb_victim_ptr | btb_278_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19738 = 9'h117 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2839 = 9'h117 == btb_victim_ptr | btb_279_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19739 = 9'h118 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2840 = 9'h118 == btb_victim_ptr | btb_280_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19740 = 9'h119 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2841 = 9'h119 == btb_victim_ptr | btb_281_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19741 = 9'h11a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2842 = 9'h11a == btb_victim_ptr | btb_282_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19742 = 9'h11b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2843 = 9'h11b == btb_victim_ptr | btb_283_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19743 = 9'h11c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2844 = 9'h11c == btb_victim_ptr | btb_284_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19744 = 9'h11d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2845 = 9'h11d == btb_victim_ptr | btb_285_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19745 = 9'h11e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2846 = 9'h11e == btb_victim_ptr | btb_286_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19746 = 9'h11f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2847 = 9'h11f == btb_victim_ptr | btb_287_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19747 = 9'h120 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2848 = 9'h120 == btb_victim_ptr | btb_288_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19748 = 9'h121 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2849 = 9'h121 == btb_victim_ptr | btb_289_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19749 = 9'h122 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2850 = 9'h122 == btb_victim_ptr | btb_290_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19750 = 9'h123 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2851 = 9'h123 == btb_victim_ptr | btb_291_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19751 = 9'h124 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2852 = 9'h124 == btb_victim_ptr | btb_292_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19752 = 9'h125 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2853 = 9'h125 == btb_victim_ptr | btb_293_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19753 = 9'h126 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2854 = 9'h126 == btb_victim_ptr | btb_294_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19754 = 9'h127 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2855 = 9'h127 == btb_victim_ptr | btb_295_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19755 = 9'h128 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2856 = 9'h128 == btb_victim_ptr | btb_296_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19756 = 9'h129 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2857 = 9'h129 == btb_victim_ptr | btb_297_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19757 = 9'h12a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2858 = 9'h12a == btb_victim_ptr | btb_298_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19758 = 9'h12b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2859 = 9'h12b == btb_victim_ptr | btb_299_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19759 = 9'h12c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2860 = 9'h12c == btb_victim_ptr | btb_300_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19760 = 9'h12d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2861 = 9'h12d == btb_victim_ptr | btb_301_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19761 = 9'h12e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2862 = 9'h12e == btb_victim_ptr | btb_302_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19762 = 9'h12f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2863 = 9'h12f == btb_victim_ptr | btb_303_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19763 = 9'h130 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2864 = 9'h130 == btb_victim_ptr | btb_304_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19764 = 9'h131 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2865 = 9'h131 == btb_victim_ptr | btb_305_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19765 = 9'h132 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2866 = 9'h132 == btb_victim_ptr | btb_306_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19766 = 9'h133 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2867 = 9'h133 == btb_victim_ptr | btb_307_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19767 = 9'h134 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2868 = 9'h134 == btb_victim_ptr | btb_308_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19768 = 9'h135 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2869 = 9'h135 == btb_victim_ptr | btb_309_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19769 = 9'h136 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2870 = 9'h136 == btb_victim_ptr | btb_310_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19770 = 9'h137 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2871 = 9'h137 == btb_victim_ptr | btb_311_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19771 = 9'h138 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2872 = 9'h138 == btb_victim_ptr | btb_312_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19772 = 9'h139 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2873 = 9'h139 == btb_victim_ptr | btb_313_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19773 = 9'h13a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2874 = 9'h13a == btb_victim_ptr | btb_314_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19774 = 9'h13b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2875 = 9'h13b == btb_victim_ptr | btb_315_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19775 = 9'h13c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2876 = 9'h13c == btb_victim_ptr | btb_316_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19776 = 9'h13d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2877 = 9'h13d == btb_victim_ptr | btb_317_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19777 = 9'h13e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2878 = 9'h13e == btb_victim_ptr | btb_318_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19778 = 9'h13f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2879 = 9'h13f == btb_victim_ptr | btb_319_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19779 = 9'h140 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2880 = 9'h140 == btb_victim_ptr | btb_320_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19780 = 9'h141 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2881 = 9'h141 == btb_victim_ptr | btb_321_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19781 = 9'h142 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2882 = 9'h142 == btb_victim_ptr | btb_322_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19782 = 9'h143 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2883 = 9'h143 == btb_victim_ptr | btb_323_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19783 = 9'h144 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2884 = 9'h144 == btb_victim_ptr | btb_324_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19784 = 9'h145 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2885 = 9'h145 == btb_victim_ptr | btb_325_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19785 = 9'h146 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2886 = 9'h146 == btb_victim_ptr | btb_326_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19786 = 9'h147 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2887 = 9'h147 == btb_victim_ptr | btb_327_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19787 = 9'h148 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2888 = 9'h148 == btb_victim_ptr | btb_328_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19788 = 9'h149 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2889 = 9'h149 == btb_victim_ptr | btb_329_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19789 = 9'h14a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2890 = 9'h14a == btb_victim_ptr | btb_330_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19790 = 9'h14b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2891 = 9'h14b == btb_victim_ptr | btb_331_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19791 = 9'h14c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2892 = 9'h14c == btb_victim_ptr | btb_332_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19792 = 9'h14d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2893 = 9'h14d == btb_victim_ptr | btb_333_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19793 = 9'h14e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2894 = 9'h14e == btb_victim_ptr | btb_334_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19794 = 9'h14f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2895 = 9'h14f == btb_victim_ptr | btb_335_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19795 = 9'h150 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2896 = 9'h150 == btb_victim_ptr | btb_336_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19796 = 9'h151 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2897 = 9'h151 == btb_victim_ptr | btb_337_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19797 = 9'h152 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2898 = 9'h152 == btb_victim_ptr | btb_338_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19798 = 9'h153 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2899 = 9'h153 == btb_victim_ptr | btb_339_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19799 = 9'h154 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2900 = 9'h154 == btb_victim_ptr | btb_340_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19800 = 9'h155 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2901 = 9'h155 == btb_victim_ptr | btb_341_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19801 = 9'h156 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2902 = 9'h156 == btb_victim_ptr | btb_342_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19802 = 9'h157 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2903 = 9'h157 == btb_victim_ptr | btb_343_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19803 = 9'h158 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2904 = 9'h158 == btb_victim_ptr | btb_344_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19804 = 9'h159 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2905 = 9'h159 == btb_victim_ptr | btb_345_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19805 = 9'h15a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2906 = 9'h15a == btb_victim_ptr | btb_346_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19806 = 9'h15b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2907 = 9'h15b == btb_victim_ptr | btb_347_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19807 = 9'h15c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2908 = 9'h15c == btb_victim_ptr | btb_348_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19808 = 9'h15d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2909 = 9'h15d == btb_victim_ptr | btb_349_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19809 = 9'h15e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2910 = 9'h15e == btb_victim_ptr | btb_350_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19810 = 9'h15f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2911 = 9'h15f == btb_victim_ptr | btb_351_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19811 = 9'h160 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2912 = 9'h160 == btb_victim_ptr | btb_352_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19812 = 9'h161 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2913 = 9'h161 == btb_victim_ptr | btb_353_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19813 = 9'h162 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2914 = 9'h162 == btb_victim_ptr | btb_354_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19814 = 9'h163 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2915 = 9'h163 == btb_victim_ptr | btb_355_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19815 = 9'h164 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2916 = 9'h164 == btb_victim_ptr | btb_356_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19816 = 9'h165 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2917 = 9'h165 == btb_victim_ptr | btb_357_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19817 = 9'h166 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2918 = 9'h166 == btb_victim_ptr | btb_358_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19818 = 9'h167 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2919 = 9'h167 == btb_victim_ptr | btb_359_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19819 = 9'h168 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2920 = 9'h168 == btb_victim_ptr | btb_360_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19820 = 9'h169 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2921 = 9'h169 == btb_victim_ptr | btb_361_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19821 = 9'h16a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2922 = 9'h16a == btb_victim_ptr | btb_362_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19822 = 9'h16b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2923 = 9'h16b == btb_victim_ptr | btb_363_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19823 = 9'h16c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2924 = 9'h16c == btb_victim_ptr | btb_364_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19824 = 9'h16d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2925 = 9'h16d == btb_victim_ptr | btb_365_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19825 = 9'h16e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2926 = 9'h16e == btb_victim_ptr | btb_366_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19826 = 9'h16f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2927 = 9'h16f == btb_victim_ptr | btb_367_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19827 = 9'h170 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2928 = 9'h170 == btb_victim_ptr | btb_368_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19828 = 9'h171 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2929 = 9'h171 == btb_victim_ptr | btb_369_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19829 = 9'h172 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2930 = 9'h172 == btb_victim_ptr | btb_370_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19830 = 9'h173 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2931 = 9'h173 == btb_victim_ptr | btb_371_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19831 = 9'h174 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2932 = 9'h174 == btb_victim_ptr | btb_372_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19832 = 9'h175 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2933 = 9'h175 == btb_victim_ptr | btb_373_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19833 = 9'h176 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2934 = 9'h176 == btb_victim_ptr | btb_374_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19834 = 9'h177 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2935 = 9'h177 == btb_victim_ptr | btb_375_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19835 = 9'h178 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2936 = 9'h178 == btb_victim_ptr | btb_376_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19836 = 9'h179 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2937 = 9'h179 == btb_victim_ptr | btb_377_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19837 = 9'h17a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2938 = 9'h17a == btb_victim_ptr | btb_378_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19838 = 9'h17b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2939 = 9'h17b == btb_victim_ptr | btb_379_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19839 = 9'h17c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2940 = 9'h17c == btb_victim_ptr | btb_380_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19840 = 9'h17d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2941 = 9'h17d == btb_victim_ptr | btb_381_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19841 = 9'h17e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2942 = 9'h17e == btb_victim_ptr | btb_382_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19842 = 9'h17f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2943 = 9'h17f == btb_victim_ptr | btb_383_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19843 = 9'h180 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2944 = 9'h180 == btb_victim_ptr | btb_384_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19844 = 9'h181 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2945 = 9'h181 == btb_victim_ptr | btb_385_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19845 = 9'h182 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2946 = 9'h182 == btb_victim_ptr | btb_386_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19846 = 9'h183 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2947 = 9'h183 == btb_victim_ptr | btb_387_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19847 = 9'h184 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2948 = 9'h184 == btb_victim_ptr | btb_388_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19848 = 9'h185 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2949 = 9'h185 == btb_victim_ptr | btb_389_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19849 = 9'h186 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2950 = 9'h186 == btb_victim_ptr | btb_390_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19850 = 9'h187 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2951 = 9'h187 == btb_victim_ptr | btb_391_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19851 = 9'h188 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2952 = 9'h188 == btb_victim_ptr | btb_392_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19852 = 9'h189 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2953 = 9'h189 == btb_victim_ptr | btb_393_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19853 = 9'h18a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2954 = 9'h18a == btb_victim_ptr | btb_394_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19854 = 9'h18b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2955 = 9'h18b == btb_victim_ptr | btb_395_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19855 = 9'h18c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2956 = 9'h18c == btb_victim_ptr | btb_396_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19856 = 9'h18d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2957 = 9'h18d == btb_victim_ptr | btb_397_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19857 = 9'h18e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2958 = 9'h18e == btb_victim_ptr | btb_398_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19858 = 9'h18f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2959 = 9'h18f == btb_victim_ptr | btb_399_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19859 = 9'h190 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2960 = 9'h190 == btb_victim_ptr | btb_400_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19860 = 9'h191 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2961 = 9'h191 == btb_victim_ptr | btb_401_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19861 = 9'h192 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2962 = 9'h192 == btb_victim_ptr | btb_402_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19862 = 9'h193 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2963 = 9'h193 == btb_victim_ptr | btb_403_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19863 = 9'h194 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2964 = 9'h194 == btb_victim_ptr | btb_404_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19864 = 9'h195 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2965 = 9'h195 == btb_victim_ptr | btb_405_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19865 = 9'h196 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2966 = 9'h196 == btb_victim_ptr | btb_406_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19866 = 9'h197 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2967 = 9'h197 == btb_victim_ptr | btb_407_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19867 = 9'h198 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2968 = 9'h198 == btb_victim_ptr | btb_408_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19868 = 9'h199 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2969 = 9'h199 == btb_victim_ptr | btb_409_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19869 = 9'h19a == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2970 = 9'h19a == btb_victim_ptr | btb_410_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19870 = 9'h19b == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2971 = 9'h19b == btb_victim_ptr | btb_411_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19871 = 9'h19c == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2972 = 9'h19c == btb_victim_ptr | btb_412_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19872 = 9'h19d == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2973 = 9'h19d == btb_victim_ptr | btb_413_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19873 = 9'h19e == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2974 = 9'h19e == btb_victim_ptr | btb_414_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19874 = 9'h19f == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2975 = 9'h19f == btb_victim_ptr | btb_415_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19875 = 9'h1a0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2976 = 9'h1a0 == btb_victim_ptr | btb_416_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19876 = 9'h1a1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2977 = 9'h1a1 == btb_victim_ptr | btb_417_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19877 = 9'h1a2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2978 = 9'h1a2 == btb_victim_ptr | btb_418_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19878 = 9'h1a3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2979 = 9'h1a3 == btb_victim_ptr | btb_419_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19879 = 9'h1a4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2980 = 9'h1a4 == btb_victim_ptr | btb_420_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19880 = 9'h1a5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2981 = 9'h1a5 == btb_victim_ptr | btb_421_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19881 = 9'h1a6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2982 = 9'h1a6 == btb_victim_ptr | btb_422_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19882 = 9'h1a7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2983 = 9'h1a7 == btb_victim_ptr | btb_423_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19883 = 9'h1a8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2984 = 9'h1a8 == btb_victim_ptr | btb_424_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19884 = 9'h1a9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2985 = 9'h1a9 == btb_victim_ptr | btb_425_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19885 = 9'h1aa == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2986 = 9'h1aa == btb_victim_ptr | btb_426_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19886 = 9'h1ab == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2987 = 9'h1ab == btb_victim_ptr | btb_427_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19887 = 9'h1ac == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2988 = 9'h1ac == btb_victim_ptr | btb_428_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19888 = 9'h1ad == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2989 = 9'h1ad == btb_victim_ptr | btb_429_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19889 = 9'h1ae == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2990 = 9'h1ae == btb_victim_ptr | btb_430_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19890 = 9'h1af == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2991 = 9'h1af == btb_victim_ptr | btb_431_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19891 = 9'h1b0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2992 = 9'h1b0 == btb_victim_ptr | btb_432_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19892 = 9'h1b1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2993 = 9'h1b1 == btb_victim_ptr | btb_433_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19893 = 9'h1b2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2994 = 9'h1b2 == btb_victim_ptr | btb_434_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19894 = 9'h1b3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2995 = 9'h1b3 == btb_victim_ptr | btb_435_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19895 = 9'h1b4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2996 = 9'h1b4 == btb_victim_ptr | btb_436_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19896 = 9'h1b5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2997 = 9'h1b5 == btb_victim_ptr | btb_437_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19897 = 9'h1b6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2998 = 9'h1b6 == btb_victim_ptr | btb_438_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19898 = 9'h1b7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_2999 = 9'h1b7 == btb_victim_ptr | btb_439_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19899 = 9'h1b8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3000 = 9'h1b8 == btb_victim_ptr | btb_440_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19900 = 9'h1b9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3001 = 9'h1b9 == btb_victim_ptr | btb_441_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19901 = 9'h1ba == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3002 = 9'h1ba == btb_victim_ptr | btb_442_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19902 = 9'h1bb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3003 = 9'h1bb == btb_victim_ptr | btb_443_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19903 = 9'h1bc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3004 = 9'h1bc == btb_victim_ptr | btb_444_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19904 = 9'h1bd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3005 = 9'h1bd == btb_victim_ptr | btb_445_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19905 = 9'h1be == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3006 = 9'h1be == btb_victim_ptr | btb_446_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19906 = 9'h1bf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3007 = 9'h1bf == btb_victim_ptr | btb_447_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19907 = 9'h1c0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3008 = 9'h1c0 == btb_victim_ptr | btb_448_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19908 = 9'h1c1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3009 = 9'h1c1 == btb_victim_ptr | btb_449_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19909 = 9'h1c2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3010 = 9'h1c2 == btb_victim_ptr | btb_450_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19910 = 9'h1c3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3011 = 9'h1c3 == btb_victim_ptr | btb_451_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19911 = 9'h1c4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3012 = 9'h1c4 == btb_victim_ptr | btb_452_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19912 = 9'h1c5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3013 = 9'h1c5 == btb_victim_ptr | btb_453_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19913 = 9'h1c6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3014 = 9'h1c6 == btb_victim_ptr | btb_454_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19914 = 9'h1c7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3015 = 9'h1c7 == btb_victim_ptr | btb_455_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19915 = 9'h1c8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3016 = 9'h1c8 == btb_victim_ptr | btb_456_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19916 = 9'h1c9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3017 = 9'h1c9 == btb_victim_ptr | btb_457_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19917 = 9'h1ca == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3018 = 9'h1ca == btb_victim_ptr | btb_458_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19918 = 9'h1cb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3019 = 9'h1cb == btb_victim_ptr | btb_459_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19919 = 9'h1cc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3020 = 9'h1cc == btb_victim_ptr | btb_460_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19920 = 9'h1cd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3021 = 9'h1cd == btb_victim_ptr | btb_461_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19921 = 9'h1ce == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3022 = 9'h1ce == btb_victim_ptr | btb_462_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19922 = 9'h1cf == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3023 = 9'h1cf == btb_victim_ptr | btb_463_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19923 = 9'h1d0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3024 = 9'h1d0 == btb_victim_ptr | btb_464_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19924 = 9'h1d1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3025 = 9'h1d1 == btb_victim_ptr | btb_465_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19925 = 9'h1d2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3026 = 9'h1d2 == btb_victim_ptr | btb_466_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19926 = 9'h1d3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3027 = 9'h1d3 == btb_victim_ptr | btb_467_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19927 = 9'h1d4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3028 = 9'h1d4 == btb_victim_ptr | btb_468_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19928 = 9'h1d5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3029 = 9'h1d5 == btb_victim_ptr | btb_469_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19929 = 9'h1d6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3030 = 9'h1d6 == btb_victim_ptr | btb_470_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19930 = 9'h1d7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3031 = 9'h1d7 == btb_victim_ptr | btb_471_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19931 = 9'h1d8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3032 = 9'h1d8 == btb_victim_ptr | btb_472_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19932 = 9'h1d9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3033 = 9'h1d9 == btb_victim_ptr | btb_473_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19933 = 9'h1da == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3034 = 9'h1da == btb_victim_ptr | btb_474_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19934 = 9'h1db == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3035 = 9'h1db == btb_victim_ptr | btb_475_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19935 = 9'h1dc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3036 = 9'h1dc == btb_victim_ptr | btb_476_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19936 = 9'h1dd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3037 = 9'h1dd == btb_victim_ptr | btb_477_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19937 = 9'h1de == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3038 = 9'h1de == btb_victim_ptr | btb_478_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19938 = 9'h1df == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3039 = 9'h1df == btb_victim_ptr | btb_479_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19939 = 9'h1e0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3040 = 9'h1e0 == btb_victim_ptr | btb_480_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19940 = 9'h1e1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3041 = 9'h1e1 == btb_victim_ptr | btb_481_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19941 = 9'h1e2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3042 = 9'h1e2 == btb_victim_ptr | btb_482_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19942 = 9'h1e3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3043 = 9'h1e3 == btb_victim_ptr | btb_483_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19943 = 9'h1e4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3044 = 9'h1e4 == btb_victim_ptr | btb_484_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19944 = 9'h1e5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3045 = 9'h1e5 == btb_victim_ptr | btb_485_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19945 = 9'h1e6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3046 = 9'h1e6 == btb_victim_ptr | btb_486_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19946 = 9'h1e7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3047 = 9'h1e7 == btb_victim_ptr | btb_487_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19947 = 9'h1e8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3048 = 9'h1e8 == btb_victim_ptr | btb_488_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19948 = 9'h1e9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3049 = 9'h1e9 == btb_victim_ptr | btb_489_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19949 = 9'h1ea == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3050 = 9'h1ea == btb_victim_ptr | btb_490_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19950 = 9'h1eb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3051 = 9'h1eb == btb_victim_ptr | btb_491_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19951 = 9'h1ec == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3052 = 9'h1ec == btb_victim_ptr | btb_492_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19952 = 9'h1ed == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3053 = 9'h1ed == btb_victim_ptr | btb_493_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19953 = 9'h1ee == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3054 = 9'h1ee == btb_victim_ptr | btb_494_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19954 = 9'h1ef == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3055 = 9'h1ef == btb_victim_ptr | btb_495_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19955 = 9'h1f0 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3056 = 9'h1f0 == btb_victim_ptr | btb_496_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19956 = 9'h1f1 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3057 = 9'h1f1 == btb_victim_ptr | btb_497_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19957 = 9'h1f2 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3058 = 9'h1f2 == btb_victim_ptr | btb_498_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19958 = 9'h1f3 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3059 = 9'h1f3 == btb_victim_ptr | btb_499_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19959 = 9'h1f4 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3060 = 9'h1f4 == btb_victim_ptr | btb_500_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19960 = 9'h1f5 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3061 = 9'h1f5 == btb_victim_ptr | btb_501_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19961 = 9'h1f6 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3062 = 9'h1f6 == btb_victim_ptr | btb_502_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19962 = 9'h1f7 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3063 = 9'h1f7 == btb_victim_ptr | btb_503_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19963 = 9'h1f8 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3064 = 9'h1f8 == btb_victim_ptr | btb_504_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19964 = 9'h1f9 == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3065 = 9'h1f9 == btb_victim_ptr | btb_505_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19965 = 9'h1fa == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3066 = 9'h1fa == btb_victim_ptr | btb_506_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19966 = 9'h1fb == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3067 = 9'h1fb == btb_victim_ptr | btb_507_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19967 = 9'h1fc == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3068 = 9'h1fc == btb_victim_ptr | btb_508_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19968 = 9'h1fd == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3069 = 9'h1fd == btb_victim_ptr | btb_509_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19969 = 9'h1fe == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3070 = 9'h1fe == btb_victim_ptr | btb_510_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_19970 = 9'h1ff == btb_victim_ptr; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire  _GEN_3071 = 9'h1ff == btb_victim_ptr | btb_511_valid; // @[branch_predictor.scala 30:22 63:{35,35}]
  wire [9:0] _GEN_3072 = 9'h0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_0_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3073 = 9'h1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_1_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3074 = 9'h2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_2_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3075 = 9'h3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_3_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3076 = 9'h4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_4_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3077 = 9'h5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_5_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3078 = 9'h6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_6_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3079 = 9'h7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_7_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3080 = 9'h8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_8_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3081 = 9'h9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_9_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3082 = 9'ha == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_10_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3083 = 9'hb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_11_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3084 = 9'hc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_12_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3085 = 9'hd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_13_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3086 = 9'he == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_14_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3087 = 9'hf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_15_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3088 = 9'h10 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_16_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3089 = 9'h11 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_17_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3090 = 9'h12 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_18_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3091 = 9'h13 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_19_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3092 = 9'h14 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_20_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3093 = 9'h15 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_21_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3094 = 9'h16 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_22_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3095 = 9'h17 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_23_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3096 = 9'h18 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_24_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3097 = 9'h19 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_25_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3098 = 9'h1a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_26_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3099 = 9'h1b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_27_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3100 = 9'h1c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_28_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3101 = 9'h1d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_29_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3102 = 9'h1e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_30_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3103 = 9'h1f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_31_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3104 = 9'h20 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_32_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3105 = 9'h21 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_33_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3106 = 9'h22 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_34_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3107 = 9'h23 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_35_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3108 = 9'h24 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_36_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3109 = 9'h25 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_37_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3110 = 9'h26 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_38_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3111 = 9'h27 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_39_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3112 = 9'h28 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_40_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3113 = 9'h29 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_41_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3114 = 9'h2a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_42_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3115 = 9'h2b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_43_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3116 = 9'h2c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_44_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3117 = 9'h2d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_45_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3118 = 9'h2e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_46_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3119 = 9'h2f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_47_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3120 = 9'h30 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_48_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3121 = 9'h31 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_49_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3122 = 9'h32 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_50_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3123 = 9'h33 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_51_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3124 = 9'h34 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_52_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3125 = 9'h35 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_53_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3126 = 9'h36 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_54_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3127 = 9'h37 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_55_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3128 = 9'h38 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_56_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3129 = 9'h39 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_57_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3130 = 9'h3a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_58_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3131 = 9'h3b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_59_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3132 = 9'h3c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_60_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3133 = 9'h3d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_61_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3134 = 9'h3e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_62_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3135 = 9'h3f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_63_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3136 = 9'h40 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_64_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3137 = 9'h41 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_65_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3138 = 9'h42 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_66_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3139 = 9'h43 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_67_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3140 = 9'h44 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_68_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3141 = 9'h45 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_69_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3142 = 9'h46 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_70_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3143 = 9'h47 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_71_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3144 = 9'h48 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_72_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3145 = 9'h49 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_73_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3146 = 9'h4a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_74_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3147 = 9'h4b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_75_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3148 = 9'h4c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_76_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3149 = 9'h4d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_77_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3150 = 9'h4e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_78_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3151 = 9'h4f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_79_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3152 = 9'h50 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_80_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3153 = 9'h51 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_81_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3154 = 9'h52 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_82_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3155 = 9'h53 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_83_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3156 = 9'h54 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_84_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3157 = 9'h55 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_85_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3158 = 9'h56 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_86_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3159 = 9'h57 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_87_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3160 = 9'h58 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_88_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3161 = 9'h59 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_89_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3162 = 9'h5a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_90_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3163 = 9'h5b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_91_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3164 = 9'h5c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_92_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3165 = 9'h5d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_93_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3166 = 9'h5e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_94_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3167 = 9'h5f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_95_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3168 = 9'h60 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_96_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3169 = 9'h61 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_97_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3170 = 9'h62 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_98_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3171 = 9'h63 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_99_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3172 = 9'h64 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_100_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3173 = 9'h65 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_101_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3174 = 9'h66 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_102_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3175 = 9'h67 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_103_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3176 = 9'h68 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_104_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3177 = 9'h69 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_105_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3178 = 9'h6a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_106_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3179 = 9'h6b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_107_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3180 = 9'h6c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_108_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3181 = 9'h6d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_109_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3182 = 9'h6e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_110_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3183 = 9'h6f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_111_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3184 = 9'h70 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_112_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3185 = 9'h71 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_113_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3186 = 9'h72 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_114_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3187 = 9'h73 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_115_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3188 = 9'h74 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_116_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3189 = 9'h75 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_117_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3190 = 9'h76 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_118_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3191 = 9'h77 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_119_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3192 = 9'h78 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_120_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3193 = 9'h79 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_121_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3194 = 9'h7a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_122_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3195 = 9'h7b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_123_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3196 = 9'h7c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_124_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3197 = 9'h7d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_125_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3198 = 9'h7e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_126_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3199 = 9'h7f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_127_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3200 = 9'h80 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_128_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3201 = 9'h81 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_129_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3202 = 9'h82 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_130_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3203 = 9'h83 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_131_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3204 = 9'h84 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_132_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3205 = 9'h85 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_133_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3206 = 9'h86 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_134_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3207 = 9'h87 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_135_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3208 = 9'h88 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_136_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3209 = 9'h89 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_137_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3210 = 9'h8a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_138_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3211 = 9'h8b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_139_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3212 = 9'h8c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_140_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3213 = 9'h8d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_141_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3214 = 9'h8e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_142_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3215 = 9'h8f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_143_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3216 = 9'h90 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_144_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3217 = 9'h91 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_145_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3218 = 9'h92 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_146_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3219 = 9'h93 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_147_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3220 = 9'h94 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_148_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3221 = 9'h95 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_149_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3222 = 9'h96 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_150_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3223 = 9'h97 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_151_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3224 = 9'h98 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_152_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3225 = 9'h99 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_153_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3226 = 9'h9a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_154_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3227 = 9'h9b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_155_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3228 = 9'h9c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_156_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3229 = 9'h9d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_157_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3230 = 9'h9e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_158_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3231 = 9'h9f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_159_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3232 = 9'ha0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_160_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3233 = 9'ha1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_161_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3234 = 9'ha2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_162_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3235 = 9'ha3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_163_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3236 = 9'ha4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_164_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3237 = 9'ha5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_165_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3238 = 9'ha6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_166_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3239 = 9'ha7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_167_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3240 = 9'ha8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_168_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3241 = 9'ha9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_169_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3242 = 9'haa == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_170_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3243 = 9'hab == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_171_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3244 = 9'hac == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_172_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3245 = 9'had == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_173_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3246 = 9'hae == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_174_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3247 = 9'haf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_175_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3248 = 9'hb0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_176_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3249 = 9'hb1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_177_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3250 = 9'hb2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_178_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3251 = 9'hb3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_179_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3252 = 9'hb4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_180_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3253 = 9'hb5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_181_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3254 = 9'hb6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_182_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3255 = 9'hb7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_183_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3256 = 9'hb8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_184_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3257 = 9'hb9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_185_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3258 = 9'hba == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_186_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3259 = 9'hbb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_187_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3260 = 9'hbc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_188_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3261 = 9'hbd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_189_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3262 = 9'hbe == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_190_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3263 = 9'hbf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_191_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3264 = 9'hc0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_192_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3265 = 9'hc1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_193_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3266 = 9'hc2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_194_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3267 = 9'hc3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_195_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3268 = 9'hc4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_196_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3269 = 9'hc5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_197_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3270 = 9'hc6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_198_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3271 = 9'hc7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_199_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3272 = 9'hc8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_200_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3273 = 9'hc9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_201_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3274 = 9'hca == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_202_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3275 = 9'hcb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_203_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3276 = 9'hcc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_204_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3277 = 9'hcd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_205_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3278 = 9'hce == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_206_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3279 = 9'hcf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_207_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3280 = 9'hd0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_208_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3281 = 9'hd1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_209_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3282 = 9'hd2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_210_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3283 = 9'hd3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_211_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3284 = 9'hd4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_212_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3285 = 9'hd5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_213_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3286 = 9'hd6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_214_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3287 = 9'hd7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_215_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3288 = 9'hd8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_216_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3289 = 9'hd9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_217_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3290 = 9'hda == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_218_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3291 = 9'hdb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_219_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3292 = 9'hdc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_220_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3293 = 9'hdd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_221_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3294 = 9'hde == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_222_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3295 = 9'hdf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_223_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3296 = 9'he0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_224_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3297 = 9'he1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_225_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3298 = 9'he2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_226_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3299 = 9'he3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_227_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3300 = 9'he4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_228_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3301 = 9'he5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_229_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3302 = 9'he6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_230_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3303 = 9'he7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_231_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3304 = 9'he8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_232_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3305 = 9'he9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_233_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3306 = 9'hea == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_234_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3307 = 9'heb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_235_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3308 = 9'hec == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_236_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3309 = 9'hed == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_237_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3310 = 9'hee == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_238_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3311 = 9'hef == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_239_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3312 = 9'hf0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_240_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3313 = 9'hf1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_241_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3314 = 9'hf2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_242_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3315 = 9'hf3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_243_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3316 = 9'hf4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_244_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3317 = 9'hf5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_245_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3318 = 9'hf6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_246_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3319 = 9'hf7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_247_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3320 = 9'hf8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_248_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3321 = 9'hf9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_249_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3322 = 9'hfa == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_250_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3323 = 9'hfb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_251_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3324 = 9'hfc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_252_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3325 = 9'hfd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_253_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3326 = 9'hfe == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_254_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3327 = 9'hff == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_255_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3328 = 9'h100 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_256_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3329 = 9'h101 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_257_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3330 = 9'h102 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_258_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3331 = 9'h103 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_259_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3332 = 9'h104 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_260_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3333 = 9'h105 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_261_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3334 = 9'h106 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_262_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3335 = 9'h107 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_263_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3336 = 9'h108 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_264_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3337 = 9'h109 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_265_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3338 = 9'h10a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_266_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3339 = 9'h10b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_267_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3340 = 9'h10c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_268_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3341 = 9'h10d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_269_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3342 = 9'h10e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_270_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3343 = 9'h10f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_271_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3344 = 9'h110 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_272_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3345 = 9'h111 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_273_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3346 = 9'h112 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_274_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3347 = 9'h113 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_275_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3348 = 9'h114 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_276_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3349 = 9'h115 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_277_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3350 = 9'h116 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_278_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3351 = 9'h117 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_279_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3352 = 9'h118 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_280_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3353 = 9'h119 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_281_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3354 = 9'h11a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_282_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3355 = 9'h11b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_283_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3356 = 9'h11c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_284_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3357 = 9'h11d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_285_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3358 = 9'h11e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_286_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3359 = 9'h11f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_287_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3360 = 9'h120 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_288_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3361 = 9'h121 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_289_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3362 = 9'h122 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_290_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3363 = 9'h123 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_291_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3364 = 9'h124 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_292_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3365 = 9'h125 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_293_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3366 = 9'h126 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_294_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3367 = 9'h127 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_295_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3368 = 9'h128 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_296_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3369 = 9'h129 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_297_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3370 = 9'h12a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_298_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3371 = 9'h12b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_299_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3372 = 9'h12c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_300_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3373 = 9'h12d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_301_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3374 = 9'h12e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_302_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3375 = 9'h12f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_303_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3376 = 9'h130 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_304_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3377 = 9'h131 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_305_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3378 = 9'h132 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_306_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3379 = 9'h133 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_307_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3380 = 9'h134 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_308_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3381 = 9'h135 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_309_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3382 = 9'h136 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_310_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3383 = 9'h137 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_311_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3384 = 9'h138 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_312_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3385 = 9'h139 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_313_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3386 = 9'h13a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_314_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3387 = 9'h13b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_315_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3388 = 9'h13c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_316_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3389 = 9'h13d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_317_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3390 = 9'h13e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_318_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3391 = 9'h13f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_319_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3392 = 9'h140 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_320_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3393 = 9'h141 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_321_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3394 = 9'h142 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_322_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3395 = 9'h143 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_323_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3396 = 9'h144 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_324_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3397 = 9'h145 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_325_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3398 = 9'h146 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_326_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3399 = 9'h147 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_327_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3400 = 9'h148 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_328_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3401 = 9'h149 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_329_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3402 = 9'h14a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_330_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3403 = 9'h14b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_331_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3404 = 9'h14c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_332_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3405 = 9'h14d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_333_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3406 = 9'h14e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_334_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3407 = 9'h14f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_335_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3408 = 9'h150 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_336_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3409 = 9'h151 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_337_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3410 = 9'h152 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_338_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3411 = 9'h153 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_339_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3412 = 9'h154 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_340_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3413 = 9'h155 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_341_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3414 = 9'h156 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_342_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3415 = 9'h157 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_343_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3416 = 9'h158 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_344_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3417 = 9'h159 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_345_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3418 = 9'h15a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_346_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3419 = 9'h15b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_347_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3420 = 9'h15c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_348_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3421 = 9'h15d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_349_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3422 = 9'h15e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_350_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3423 = 9'h15f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_351_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3424 = 9'h160 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_352_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3425 = 9'h161 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_353_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3426 = 9'h162 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_354_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3427 = 9'h163 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_355_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3428 = 9'h164 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_356_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3429 = 9'h165 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_357_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3430 = 9'h166 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_358_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3431 = 9'h167 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_359_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3432 = 9'h168 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_360_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3433 = 9'h169 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_361_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3434 = 9'h16a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_362_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3435 = 9'h16b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_363_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3436 = 9'h16c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_364_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3437 = 9'h16d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_365_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3438 = 9'h16e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_366_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3439 = 9'h16f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_367_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3440 = 9'h170 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_368_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3441 = 9'h171 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_369_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3442 = 9'h172 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_370_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3443 = 9'h173 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_371_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3444 = 9'h174 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_372_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3445 = 9'h175 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_373_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3446 = 9'h176 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_374_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3447 = 9'h177 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_375_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3448 = 9'h178 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_376_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3449 = 9'h179 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_377_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3450 = 9'h17a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_378_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3451 = 9'h17b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_379_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3452 = 9'h17c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_380_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3453 = 9'h17d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_381_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3454 = 9'h17e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_382_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3455 = 9'h17f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_383_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3456 = 9'h180 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_384_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3457 = 9'h181 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_385_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3458 = 9'h182 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_386_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3459 = 9'h183 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_387_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3460 = 9'h184 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_388_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3461 = 9'h185 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_389_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3462 = 9'h186 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_390_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3463 = 9'h187 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_391_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3464 = 9'h188 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_392_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3465 = 9'h189 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_393_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3466 = 9'h18a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_394_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3467 = 9'h18b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_395_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3468 = 9'h18c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_396_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3469 = 9'h18d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_397_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3470 = 9'h18e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_398_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3471 = 9'h18f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_399_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3472 = 9'h190 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_400_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3473 = 9'h191 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_401_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3474 = 9'h192 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_402_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3475 = 9'h193 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_403_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3476 = 9'h194 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_404_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3477 = 9'h195 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_405_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3478 = 9'h196 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_406_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3479 = 9'h197 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_407_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3480 = 9'h198 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_408_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3481 = 9'h199 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_409_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3482 = 9'h19a == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_410_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3483 = 9'h19b == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_411_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3484 = 9'h19c == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_412_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3485 = 9'h19d == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_413_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3486 = 9'h19e == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_414_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3487 = 9'h19f == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_415_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3488 = 9'h1a0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_416_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3489 = 9'h1a1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_417_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3490 = 9'h1a2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_418_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3491 = 9'h1a3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_419_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3492 = 9'h1a4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_420_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3493 = 9'h1a5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_421_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3494 = 9'h1a6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_422_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3495 = 9'h1a7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_423_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3496 = 9'h1a8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_424_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3497 = 9'h1a9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_425_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3498 = 9'h1aa == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_426_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3499 = 9'h1ab == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_427_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3500 = 9'h1ac == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_428_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3501 = 9'h1ad == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_429_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3502 = 9'h1ae == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_430_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3503 = 9'h1af == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_431_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3504 = 9'h1b0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_432_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3505 = 9'h1b1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_433_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3506 = 9'h1b2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_434_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3507 = 9'h1b3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_435_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3508 = 9'h1b4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_436_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3509 = 9'h1b5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_437_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3510 = 9'h1b6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_438_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3511 = 9'h1b7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_439_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3512 = 9'h1b8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_440_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3513 = 9'h1b9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_441_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3514 = 9'h1ba == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_442_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3515 = 9'h1bb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_443_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3516 = 9'h1bc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_444_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3517 = 9'h1bd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_445_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3518 = 9'h1be == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_446_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3519 = 9'h1bf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_447_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3520 = 9'h1c0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_448_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3521 = 9'h1c1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_449_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3522 = 9'h1c2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_450_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3523 = 9'h1c3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_451_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3524 = 9'h1c4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_452_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3525 = 9'h1c5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_453_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3526 = 9'h1c6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_454_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3527 = 9'h1c7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_455_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3528 = 9'h1c8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_456_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3529 = 9'h1c9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_457_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3530 = 9'h1ca == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_458_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3531 = 9'h1cb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_459_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3532 = 9'h1cc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_460_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3533 = 9'h1cd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_461_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3534 = 9'h1ce == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_462_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3535 = 9'h1cf == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_463_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3536 = 9'h1d0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_464_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3537 = 9'h1d1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_465_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3538 = 9'h1d2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_466_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3539 = 9'h1d3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_467_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3540 = 9'h1d4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_468_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3541 = 9'h1d5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_469_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3542 = 9'h1d6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_470_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3543 = 9'h1d7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_471_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3544 = 9'h1d8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_472_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3545 = 9'h1d9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_473_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3546 = 9'h1da == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_474_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3547 = 9'h1db == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_475_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3548 = 9'h1dc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_476_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3549 = 9'h1dd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_477_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3550 = 9'h1de == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_478_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3551 = 9'h1df == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_479_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3552 = 9'h1e0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_480_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3553 = 9'h1e1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_481_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3554 = 9'h1e2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_482_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3555 = 9'h1e3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_483_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3556 = 9'h1e4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_484_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3557 = 9'h1e5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_485_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3558 = 9'h1e6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_486_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3559 = 9'h1e7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_487_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3560 = 9'h1e8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_488_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3561 = 9'h1e9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_489_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3562 = 9'h1ea == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_490_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3563 = 9'h1eb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_491_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3564 = 9'h1ec == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_492_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3565 = 9'h1ed == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_493_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3566 = 9'h1ee == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_494_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3567 = 9'h1ef == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_495_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3568 = 9'h1f0 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_496_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3569 = 9'h1f1 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_497_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3570 = 9'h1f2 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_498_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3571 = 9'h1f3 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_499_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3572 = 9'h1f4 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_500_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3573 = 9'h1f5 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_501_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3574 = 9'h1f6 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_502_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3575 = 9'h1f7 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_503_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3576 = 9'h1f8 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_504_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3577 = 9'h1f9 == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_505_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3578 = 9'h1fa == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_506_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3579 = 9'h1fb == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_507_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3580 = 9'h1fc == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_508_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3581 = 9'h1fd == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_509_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3582 = 9'h1fe == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_510_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [9:0] _GEN_3583 = 9'h1ff == btb_victim_ptr ? io_i_branch_resolve_pack_pc[12:3] : btb_511_tag; // @[branch_predictor.scala 30:22 64:{33,33}]
  wire [63:0] _GEN_3584 = 9'h0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_0_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3585 = 9'h1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_1_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3586 = 9'h2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_2_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3587 = 9'h3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_3_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3588 = 9'h4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_4_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3589 = 9'h5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_5_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3590 = 9'h6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_6_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3591 = 9'h7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_7_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3592 = 9'h8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_8_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3593 = 9'h9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_9_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3594 = 9'ha == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_10_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3595 = 9'hb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_11_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3596 = 9'hc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_12_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3597 = 9'hd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_13_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3598 = 9'he == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_14_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3599 = 9'hf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_15_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3600 = 9'h10 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_16_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3601 = 9'h11 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_17_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3602 = 9'h12 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_18_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3603 = 9'h13 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_19_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3604 = 9'h14 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_20_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3605 = 9'h15 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_21_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3606 = 9'h16 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_22_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3607 = 9'h17 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_23_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3608 = 9'h18 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_24_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3609 = 9'h19 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_25_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3610 = 9'h1a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_26_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3611 = 9'h1b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_27_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3612 = 9'h1c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_28_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3613 = 9'h1d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_29_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3614 = 9'h1e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_30_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3615 = 9'h1f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_31_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3616 = 9'h20 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_32_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3617 = 9'h21 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_33_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3618 = 9'h22 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_34_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3619 = 9'h23 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_35_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3620 = 9'h24 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_36_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3621 = 9'h25 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_37_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3622 = 9'h26 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_38_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3623 = 9'h27 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_39_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3624 = 9'h28 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_40_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3625 = 9'h29 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_41_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3626 = 9'h2a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_42_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3627 = 9'h2b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_43_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3628 = 9'h2c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_44_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3629 = 9'h2d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_45_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3630 = 9'h2e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_46_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3631 = 9'h2f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_47_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3632 = 9'h30 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_48_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3633 = 9'h31 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_49_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3634 = 9'h32 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_50_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3635 = 9'h33 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_51_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3636 = 9'h34 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_52_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3637 = 9'h35 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_53_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3638 = 9'h36 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_54_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3639 = 9'h37 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_55_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3640 = 9'h38 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_56_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3641 = 9'h39 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_57_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3642 = 9'h3a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_58_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3643 = 9'h3b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_59_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3644 = 9'h3c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_60_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3645 = 9'h3d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_61_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3646 = 9'h3e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_62_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3647 = 9'h3f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_63_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3648 = 9'h40 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_64_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3649 = 9'h41 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_65_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3650 = 9'h42 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_66_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3651 = 9'h43 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_67_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3652 = 9'h44 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_68_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3653 = 9'h45 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_69_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3654 = 9'h46 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_70_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3655 = 9'h47 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_71_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3656 = 9'h48 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_72_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3657 = 9'h49 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_73_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3658 = 9'h4a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_74_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3659 = 9'h4b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_75_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3660 = 9'h4c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_76_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3661 = 9'h4d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_77_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3662 = 9'h4e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_78_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3663 = 9'h4f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_79_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3664 = 9'h50 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_80_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3665 = 9'h51 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_81_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3666 = 9'h52 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_82_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3667 = 9'h53 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_83_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3668 = 9'h54 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_84_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3669 = 9'h55 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_85_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3670 = 9'h56 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_86_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3671 = 9'h57 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_87_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3672 = 9'h58 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_88_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3673 = 9'h59 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_89_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3674 = 9'h5a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_90_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3675 = 9'h5b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_91_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3676 = 9'h5c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_92_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3677 = 9'h5d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_93_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3678 = 9'h5e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_94_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3679 = 9'h5f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_95_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3680 = 9'h60 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_96_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3681 = 9'h61 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_97_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3682 = 9'h62 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_98_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3683 = 9'h63 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_99_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3684 = 9'h64 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_100_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3685 = 9'h65 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_101_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3686 = 9'h66 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_102_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3687 = 9'h67 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_103_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3688 = 9'h68 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_104_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3689 = 9'h69 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_105_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3690 = 9'h6a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_106_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3691 = 9'h6b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_107_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3692 = 9'h6c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_108_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3693 = 9'h6d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_109_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3694 = 9'h6e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_110_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3695 = 9'h6f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_111_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3696 = 9'h70 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_112_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3697 = 9'h71 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_113_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3698 = 9'h72 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_114_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3699 = 9'h73 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_115_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3700 = 9'h74 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_116_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3701 = 9'h75 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_117_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3702 = 9'h76 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_118_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3703 = 9'h77 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_119_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3704 = 9'h78 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_120_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3705 = 9'h79 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_121_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3706 = 9'h7a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_122_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3707 = 9'h7b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_123_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3708 = 9'h7c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_124_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3709 = 9'h7d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_125_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3710 = 9'h7e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_126_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3711 = 9'h7f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_127_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3712 = 9'h80 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_128_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3713 = 9'h81 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_129_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3714 = 9'h82 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_130_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3715 = 9'h83 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_131_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3716 = 9'h84 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_132_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3717 = 9'h85 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_133_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3718 = 9'h86 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_134_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3719 = 9'h87 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_135_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3720 = 9'h88 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_136_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3721 = 9'h89 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_137_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3722 = 9'h8a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_138_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3723 = 9'h8b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_139_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3724 = 9'h8c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_140_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3725 = 9'h8d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_141_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3726 = 9'h8e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_142_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3727 = 9'h8f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_143_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3728 = 9'h90 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_144_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3729 = 9'h91 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_145_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3730 = 9'h92 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_146_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3731 = 9'h93 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_147_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3732 = 9'h94 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_148_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3733 = 9'h95 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_149_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3734 = 9'h96 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_150_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3735 = 9'h97 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_151_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3736 = 9'h98 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_152_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3737 = 9'h99 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_153_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3738 = 9'h9a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_154_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3739 = 9'h9b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_155_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3740 = 9'h9c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_156_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3741 = 9'h9d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_157_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3742 = 9'h9e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_158_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3743 = 9'h9f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_159_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3744 = 9'ha0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_160_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3745 = 9'ha1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_161_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3746 = 9'ha2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_162_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3747 = 9'ha3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_163_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3748 = 9'ha4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_164_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3749 = 9'ha5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_165_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3750 = 9'ha6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_166_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3751 = 9'ha7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_167_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3752 = 9'ha8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_168_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3753 = 9'ha9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_169_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3754 = 9'haa == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_170_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3755 = 9'hab == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_171_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3756 = 9'hac == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_172_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3757 = 9'had == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_173_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3758 = 9'hae == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_174_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3759 = 9'haf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_175_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3760 = 9'hb0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_176_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3761 = 9'hb1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_177_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3762 = 9'hb2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_178_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3763 = 9'hb3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_179_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3764 = 9'hb4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_180_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3765 = 9'hb5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_181_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3766 = 9'hb6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_182_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3767 = 9'hb7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_183_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3768 = 9'hb8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_184_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3769 = 9'hb9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_185_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3770 = 9'hba == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_186_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3771 = 9'hbb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_187_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3772 = 9'hbc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_188_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3773 = 9'hbd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_189_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3774 = 9'hbe == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_190_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3775 = 9'hbf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_191_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3776 = 9'hc0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_192_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3777 = 9'hc1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_193_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3778 = 9'hc2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_194_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3779 = 9'hc3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_195_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3780 = 9'hc4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_196_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3781 = 9'hc5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_197_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3782 = 9'hc6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_198_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3783 = 9'hc7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_199_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3784 = 9'hc8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_200_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3785 = 9'hc9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_201_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3786 = 9'hca == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_202_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3787 = 9'hcb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_203_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3788 = 9'hcc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_204_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3789 = 9'hcd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_205_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3790 = 9'hce == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_206_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3791 = 9'hcf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_207_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3792 = 9'hd0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_208_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3793 = 9'hd1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_209_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3794 = 9'hd2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_210_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3795 = 9'hd3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_211_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3796 = 9'hd4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_212_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3797 = 9'hd5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_213_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3798 = 9'hd6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_214_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3799 = 9'hd7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_215_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3800 = 9'hd8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_216_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3801 = 9'hd9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_217_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3802 = 9'hda == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_218_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3803 = 9'hdb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_219_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3804 = 9'hdc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_220_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3805 = 9'hdd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_221_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3806 = 9'hde == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_222_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3807 = 9'hdf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_223_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3808 = 9'he0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_224_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3809 = 9'he1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_225_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3810 = 9'he2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_226_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3811 = 9'he3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_227_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3812 = 9'he4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_228_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3813 = 9'he5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_229_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3814 = 9'he6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_230_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3815 = 9'he7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_231_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3816 = 9'he8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_232_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3817 = 9'he9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_233_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3818 = 9'hea == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_234_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3819 = 9'heb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_235_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3820 = 9'hec == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_236_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3821 = 9'hed == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_237_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3822 = 9'hee == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_238_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3823 = 9'hef == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_239_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3824 = 9'hf0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_240_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3825 = 9'hf1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_241_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3826 = 9'hf2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_242_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3827 = 9'hf3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_243_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3828 = 9'hf4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_244_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3829 = 9'hf5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_245_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3830 = 9'hf6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_246_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3831 = 9'hf7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_247_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3832 = 9'hf8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_248_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3833 = 9'hf9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_249_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3834 = 9'hfa == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_250_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3835 = 9'hfb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_251_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3836 = 9'hfc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_252_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3837 = 9'hfd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_253_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3838 = 9'hfe == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_254_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3839 = 9'hff == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_255_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3840 = 9'h100 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_256_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3841 = 9'h101 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_257_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3842 = 9'h102 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_258_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3843 = 9'h103 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_259_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3844 = 9'h104 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_260_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3845 = 9'h105 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_261_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3846 = 9'h106 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_262_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3847 = 9'h107 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_263_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3848 = 9'h108 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_264_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3849 = 9'h109 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_265_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3850 = 9'h10a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_266_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3851 = 9'h10b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_267_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3852 = 9'h10c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_268_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3853 = 9'h10d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_269_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3854 = 9'h10e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_270_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3855 = 9'h10f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_271_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3856 = 9'h110 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_272_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3857 = 9'h111 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_273_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3858 = 9'h112 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_274_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3859 = 9'h113 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_275_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3860 = 9'h114 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_276_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3861 = 9'h115 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_277_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3862 = 9'h116 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_278_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3863 = 9'h117 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_279_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3864 = 9'h118 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_280_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3865 = 9'h119 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_281_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3866 = 9'h11a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_282_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3867 = 9'h11b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_283_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3868 = 9'h11c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_284_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3869 = 9'h11d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_285_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3870 = 9'h11e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_286_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3871 = 9'h11f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_287_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3872 = 9'h120 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_288_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3873 = 9'h121 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_289_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3874 = 9'h122 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_290_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3875 = 9'h123 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_291_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3876 = 9'h124 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_292_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3877 = 9'h125 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_293_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3878 = 9'h126 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_294_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3879 = 9'h127 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_295_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3880 = 9'h128 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_296_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3881 = 9'h129 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_297_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3882 = 9'h12a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_298_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3883 = 9'h12b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_299_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3884 = 9'h12c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_300_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3885 = 9'h12d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_301_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3886 = 9'h12e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_302_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3887 = 9'h12f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_303_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3888 = 9'h130 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_304_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3889 = 9'h131 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_305_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3890 = 9'h132 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_306_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3891 = 9'h133 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_307_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3892 = 9'h134 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_308_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3893 = 9'h135 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_309_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3894 = 9'h136 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_310_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3895 = 9'h137 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_311_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3896 = 9'h138 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_312_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3897 = 9'h139 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_313_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3898 = 9'h13a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_314_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3899 = 9'h13b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_315_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3900 = 9'h13c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_316_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3901 = 9'h13d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_317_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3902 = 9'h13e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_318_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3903 = 9'h13f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_319_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3904 = 9'h140 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_320_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3905 = 9'h141 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_321_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3906 = 9'h142 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_322_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3907 = 9'h143 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_323_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3908 = 9'h144 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_324_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3909 = 9'h145 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_325_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3910 = 9'h146 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_326_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3911 = 9'h147 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_327_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3912 = 9'h148 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_328_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3913 = 9'h149 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_329_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3914 = 9'h14a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_330_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3915 = 9'h14b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_331_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3916 = 9'h14c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_332_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3917 = 9'h14d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_333_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3918 = 9'h14e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_334_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3919 = 9'h14f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_335_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3920 = 9'h150 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_336_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3921 = 9'h151 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_337_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3922 = 9'h152 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_338_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3923 = 9'h153 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_339_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3924 = 9'h154 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_340_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3925 = 9'h155 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_341_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3926 = 9'h156 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_342_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3927 = 9'h157 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_343_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3928 = 9'h158 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_344_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3929 = 9'h159 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_345_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3930 = 9'h15a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_346_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3931 = 9'h15b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_347_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3932 = 9'h15c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_348_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3933 = 9'h15d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_349_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3934 = 9'h15e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_350_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3935 = 9'h15f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_351_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3936 = 9'h160 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_352_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3937 = 9'h161 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_353_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3938 = 9'h162 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_354_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3939 = 9'h163 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_355_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3940 = 9'h164 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_356_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3941 = 9'h165 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_357_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3942 = 9'h166 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_358_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3943 = 9'h167 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_359_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3944 = 9'h168 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_360_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3945 = 9'h169 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_361_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3946 = 9'h16a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_362_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3947 = 9'h16b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_363_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3948 = 9'h16c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_364_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3949 = 9'h16d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_365_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3950 = 9'h16e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_366_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3951 = 9'h16f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_367_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3952 = 9'h170 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_368_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3953 = 9'h171 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_369_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3954 = 9'h172 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_370_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3955 = 9'h173 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_371_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3956 = 9'h174 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_372_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3957 = 9'h175 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_373_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3958 = 9'h176 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_374_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3959 = 9'h177 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_375_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3960 = 9'h178 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_376_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3961 = 9'h179 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_377_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3962 = 9'h17a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_378_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3963 = 9'h17b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_379_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3964 = 9'h17c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_380_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3965 = 9'h17d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_381_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3966 = 9'h17e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_382_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3967 = 9'h17f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_383_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3968 = 9'h180 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_384_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3969 = 9'h181 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_385_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3970 = 9'h182 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_386_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3971 = 9'h183 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_387_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3972 = 9'h184 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_388_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3973 = 9'h185 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_389_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3974 = 9'h186 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_390_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3975 = 9'h187 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_391_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3976 = 9'h188 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_392_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3977 = 9'h189 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_393_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3978 = 9'h18a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_394_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3979 = 9'h18b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_395_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3980 = 9'h18c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_396_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3981 = 9'h18d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_397_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3982 = 9'h18e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_398_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3983 = 9'h18f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_399_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3984 = 9'h190 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_400_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3985 = 9'h191 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_401_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3986 = 9'h192 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_402_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3987 = 9'h193 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_403_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3988 = 9'h194 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_404_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3989 = 9'h195 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_405_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3990 = 9'h196 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_406_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3991 = 9'h197 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_407_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3992 = 9'h198 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_408_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3993 = 9'h199 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_409_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3994 = 9'h19a == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_410_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3995 = 9'h19b == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_411_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3996 = 9'h19c == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_412_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3997 = 9'h19d == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_413_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3998 = 9'h19e == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_414_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_3999 = 9'h19f == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_415_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4000 = 9'h1a0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_416_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4001 = 9'h1a1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_417_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4002 = 9'h1a2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_418_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4003 = 9'h1a3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_419_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4004 = 9'h1a4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_420_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4005 = 9'h1a5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_421_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4006 = 9'h1a6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_422_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4007 = 9'h1a7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_423_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4008 = 9'h1a8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_424_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4009 = 9'h1a9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_425_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4010 = 9'h1aa == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_426_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4011 = 9'h1ab == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_427_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4012 = 9'h1ac == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_428_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4013 = 9'h1ad == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_429_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4014 = 9'h1ae == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_430_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4015 = 9'h1af == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_431_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4016 = 9'h1b0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_432_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4017 = 9'h1b1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_433_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4018 = 9'h1b2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_434_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4019 = 9'h1b3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_435_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4020 = 9'h1b4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_436_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4021 = 9'h1b5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_437_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4022 = 9'h1b6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_438_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4023 = 9'h1b7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_439_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4024 = 9'h1b8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_440_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4025 = 9'h1b9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_441_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4026 = 9'h1ba == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_442_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4027 = 9'h1bb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_443_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4028 = 9'h1bc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_444_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4029 = 9'h1bd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_445_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4030 = 9'h1be == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_446_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4031 = 9'h1bf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_447_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4032 = 9'h1c0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_448_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4033 = 9'h1c1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_449_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4034 = 9'h1c2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_450_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4035 = 9'h1c3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_451_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4036 = 9'h1c4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_452_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4037 = 9'h1c5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_453_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4038 = 9'h1c6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_454_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4039 = 9'h1c7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_455_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4040 = 9'h1c8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_456_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4041 = 9'h1c9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_457_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4042 = 9'h1ca == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_458_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4043 = 9'h1cb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_459_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4044 = 9'h1cc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_460_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4045 = 9'h1cd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_461_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4046 = 9'h1ce == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_462_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4047 = 9'h1cf == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_463_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4048 = 9'h1d0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_464_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4049 = 9'h1d1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_465_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4050 = 9'h1d2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_466_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4051 = 9'h1d3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_467_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4052 = 9'h1d4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_468_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4053 = 9'h1d5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_469_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4054 = 9'h1d6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_470_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4055 = 9'h1d7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_471_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4056 = 9'h1d8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_472_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4057 = 9'h1d9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_473_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4058 = 9'h1da == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_474_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4059 = 9'h1db == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_475_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4060 = 9'h1dc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_476_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4061 = 9'h1dd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_477_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4062 = 9'h1de == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_478_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4063 = 9'h1df == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_479_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4064 = 9'h1e0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_480_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4065 = 9'h1e1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_481_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4066 = 9'h1e2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_482_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4067 = 9'h1e3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_483_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4068 = 9'h1e4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_484_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4069 = 9'h1e5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_485_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4070 = 9'h1e6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_486_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4071 = 9'h1e7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_487_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4072 = 9'h1e8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_488_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4073 = 9'h1e9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_489_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4074 = 9'h1ea == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_490_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4075 = 9'h1eb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_491_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4076 = 9'h1ec == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_492_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4077 = 9'h1ed == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_493_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4078 = 9'h1ee == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_494_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4079 = 9'h1ef == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_495_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4080 = 9'h1f0 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_496_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4081 = 9'h1f1 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_497_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4082 = 9'h1f2 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_498_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4083 = 9'h1f3 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_499_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4084 = 9'h1f4 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_500_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4085 = 9'h1f5 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_501_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4086 = 9'h1f6 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_502_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4087 = 9'h1f7 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_503_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4088 = 9'h1f8 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_504_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4089 = 9'h1f9 == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_505_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4090 = 9'h1fa == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_506_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4091 = 9'h1fb == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_507_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4092 = 9'h1fc == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_508_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4093 = 9'h1fd == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_509_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4094 = 9'h1fe == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_510_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [63:0] _GEN_4095 = 9'h1ff == btb_victim_ptr ? io_i_branch_resolve_pack_target : btb_511_target_address; // @[branch_predictor.scala 30:22 65:{44,44}]
  wire [1:0] _btb_bht_T = io_i_branch_resolve_pack_taken ? 2'h1 : 2'h0; // @[branch_predictor.scala 68:39]
  wire [1:0] _GEN_5120 = 9'h0 == btb_victim_ptr ? _btb_bht_T : btb_0_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5121 = 9'h1 == btb_victim_ptr ? _btb_bht_T : btb_1_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5122 = 9'h2 == btb_victim_ptr ? _btb_bht_T : btb_2_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5123 = 9'h3 == btb_victim_ptr ? _btb_bht_T : btb_3_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5124 = 9'h4 == btb_victim_ptr ? _btb_bht_T : btb_4_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5125 = 9'h5 == btb_victim_ptr ? _btb_bht_T : btb_5_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5126 = 9'h6 == btb_victim_ptr ? _btb_bht_T : btb_6_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5127 = 9'h7 == btb_victim_ptr ? _btb_bht_T : btb_7_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5128 = 9'h8 == btb_victim_ptr ? _btb_bht_T : btb_8_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5129 = 9'h9 == btb_victim_ptr ? _btb_bht_T : btb_9_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5130 = 9'ha == btb_victim_ptr ? _btb_bht_T : btb_10_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5131 = 9'hb == btb_victim_ptr ? _btb_bht_T : btb_11_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5132 = 9'hc == btb_victim_ptr ? _btb_bht_T : btb_12_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5133 = 9'hd == btb_victim_ptr ? _btb_bht_T : btb_13_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5134 = 9'he == btb_victim_ptr ? _btb_bht_T : btb_14_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5135 = 9'hf == btb_victim_ptr ? _btb_bht_T : btb_15_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5136 = 9'h10 == btb_victim_ptr ? _btb_bht_T : btb_16_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5137 = 9'h11 == btb_victim_ptr ? _btb_bht_T : btb_17_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5138 = 9'h12 == btb_victim_ptr ? _btb_bht_T : btb_18_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5139 = 9'h13 == btb_victim_ptr ? _btb_bht_T : btb_19_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5140 = 9'h14 == btb_victim_ptr ? _btb_bht_T : btb_20_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5141 = 9'h15 == btb_victim_ptr ? _btb_bht_T : btb_21_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5142 = 9'h16 == btb_victim_ptr ? _btb_bht_T : btb_22_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5143 = 9'h17 == btb_victim_ptr ? _btb_bht_T : btb_23_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5144 = 9'h18 == btb_victim_ptr ? _btb_bht_T : btb_24_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5145 = 9'h19 == btb_victim_ptr ? _btb_bht_T : btb_25_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5146 = 9'h1a == btb_victim_ptr ? _btb_bht_T : btb_26_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5147 = 9'h1b == btb_victim_ptr ? _btb_bht_T : btb_27_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5148 = 9'h1c == btb_victim_ptr ? _btb_bht_T : btb_28_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5149 = 9'h1d == btb_victim_ptr ? _btb_bht_T : btb_29_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5150 = 9'h1e == btb_victim_ptr ? _btb_bht_T : btb_30_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5151 = 9'h1f == btb_victim_ptr ? _btb_bht_T : btb_31_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5152 = 9'h20 == btb_victim_ptr ? _btb_bht_T : btb_32_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5153 = 9'h21 == btb_victim_ptr ? _btb_bht_T : btb_33_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5154 = 9'h22 == btb_victim_ptr ? _btb_bht_T : btb_34_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5155 = 9'h23 == btb_victim_ptr ? _btb_bht_T : btb_35_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5156 = 9'h24 == btb_victim_ptr ? _btb_bht_T : btb_36_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5157 = 9'h25 == btb_victim_ptr ? _btb_bht_T : btb_37_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5158 = 9'h26 == btb_victim_ptr ? _btb_bht_T : btb_38_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5159 = 9'h27 == btb_victim_ptr ? _btb_bht_T : btb_39_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5160 = 9'h28 == btb_victim_ptr ? _btb_bht_T : btb_40_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5161 = 9'h29 == btb_victim_ptr ? _btb_bht_T : btb_41_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5162 = 9'h2a == btb_victim_ptr ? _btb_bht_T : btb_42_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5163 = 9'h2b == btb_victim_ptr ? _btb_bht_T : btb_43_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5164 = 9'h2c == btb_victim_ptr ? _btb_bht_T : btb_44_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5165 = 9'h2d == btb_victim_ptr ? _btb_bht_T : btb_45_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5166 = 9'h2e == btb_victim_ptr ? _btb_bht_T : btb_46_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5167 = 9'h2f == btb_victim_ptr ? _btb_bht_T : btb_47_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5168 = 9'h30 == btb_victim_ptr ? _btb_bht_T : btb_48_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5169 = 9'h31 == btb_victim_ptr ? _btb_bht_T : btb_49_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5170 = 9'h32 == btb_victim_ptr ? _btb_bht_T : btb_50_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5171 = 9'h33 == btb_victim_ptr ? _btb_bht_T : btb_51_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5172 = 9'h34 == btb_victim_ptr ? _btb_bht_T : btb_52_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5173 = 9'h35 == btb_victim_ptr ? _btb_bht_T : btb_53_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5174 = 9'h36 == btb_victim_ptr ? _btb_bht_T : btb_54_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5175 = 9'h37 == btb_victim_ptr ? _btb_bht_T : btb_55_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5176 = 9'h38 == btb_victim_ptr ? _btb_bht_T : btb_56_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5177 = 9'h39 == btb_victim_ptr ? _btb_bht_T : btb_57_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5178 = 9'h3a == btb_victim_ptr ? _btb_bht_T : btb_58_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5179 = 9'h3b == btb_victim_ptr ? _btb_bht_T : btb_59_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5180 = 9'h3c == btb_victim_ptr ? _btb_bht_T : btb_60_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5181 = 9'h3d == btb_victim_ptr ? _btb_bht_T : btb_61_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5182 = 9'h3e == btb_victim_ptr ? _btb_bht_T : btb_62_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5183 = 9'h3f == btb_victim_ptr ? _btb_bht_T : btb_63_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5184 = 9'h40 == btb_victim_ptr ? _btb_bht_T : btb_64_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5185 = 9'h41 == btb_victim_ptr ? _btb_bht_T : btb_65_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5186 = 9'h42 == btb_victim_ptr ? _btb_bht_T : btb_66_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5187 = 9'h43 == btb_victim_ptr ? _btb_bht_T : btb_67_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5188 = 9'h44 == btb_victim_ptr ? _btb_bht_T : btb_68_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5189 = 9'h45 == btb_victim_ptr ? _btb_bht_T : btb_69_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5190 = 9'h46 == btb_victim_ptr ? _btb_bht_T : btb_70_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5191 = 9'h47 == btb_victim_ptr ? _btb_bht_T : btb_71_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5192 = 9'h48 == btb_victim_ptr ? _btb_bht_T : btb_72_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5193 = 9'h49 == btb_victim_ptr ? _btb_bht_T : btb_73_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5194 = 9'h4a == btb_victim_ptr ? _btb_bht_T : btb_74_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5195 = 9'h4b == btb_victim_ptr ? _btb_bht_T : btb_75_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5196 = 9'h4c == btb_victim_ptr ? _btb_bht_T : btb_76_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5197 = 9'h4d == btb_victim_ptr ? _btb_bht_T : btb_77_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5198 = 9'h4e == btb_victim_ptr ? _btb_bht_T : btb_78_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5199 = 9'h4f == btb_victim_ptr ? _btb_bht_T : btb_79_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5200 = 9'h50 == btb_victim_ptr ? _btb_bht_T : btb_80_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5201 = 9'h51 == btb_victim_ptr ? _btb_bht_T : btb_81_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5202 = 9'h52 == btb_victim_ptr ? _btb_bht_T : btb_82_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5203 = 9'h53 == btb_victim_ptr ? _btb_bht_T : btb_83_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5204 = 9'h54 == btb_victim_ptr ? _btb_bht_T : btb_84_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5205 = 9'h55 == btb_victim_ptr ? _btb_bht_T : btb_85_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5206 = 9'h56 == btb_victim_ptr ? _btb_bht_T : btb_86_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5207 = 9'h57 == btb_victim_ptr ? _btb_bht_T : btb_87_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5208 = 9'h58 == btb_victim_ptr ? _btb_bht_T : btb_88_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5209 = 9'h59 == btb_victim_ptr ? _btb_bht_T : btb_89_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5210 = 9'h5a == btb_victim_ptr ? _btb_bht_T : btb_90_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5211 = 9'h5b == btb_victim_ptr ? _btb_bht_T : btb_91_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5212 = 9'h5c == btb_victim_ptr ? _btb_bht_T : btb_92_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5213 = 9'h5d == btb_victim_ptr ? _btb_bht_T : btb_93_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5214 = 9'h5e == btb_victim_ptr ? _btb_bht_T : btb_94_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5215 = 9'h5f == btb_victim_ptr ? _btb_bht_T : btb_95_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5216 = 9'h60 == btb_victim_ptr ? _btb_bht_T : btb_96_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5217 = 9'h61 == btb_victim_ptr ? _btb_bht_T : btb_97_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5218 = 9'h62 == btb_victim_ptr ? _btb_bht_T : btb_98_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5219 = 9'h63 == btb_victim_ptr ? _btb_bht_T : btb_99_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5220 = 9'h64 == btb_victim_ptr ? _btb_bht_T : btb_100_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5221 = 9'h65 == btb_victim_ptr ? _btb_bht_T : btb_101_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5222 = 9'h66 == btb_victim_ptr ? _btb_bht_T : btb_102_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5223 = 9'h67 == btb_victim_ptr ? _btb_bht_T : btb_103_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5224 = 9'h68 == btb_victim_ptr ? _btb_bht_T : btb_104_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5225 = 9'h69 == btb_victim_ptr ? _btb_bht_T : btb_105_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5226 = 9'h6a == btb_victim_ptr ? _btb_bht_T : btb_106_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5227 = 9'h6b == btb_victim_ptr ? _btb_bht_T : btb_107_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5228 = 9'h6c == btb_victim_ptr ? _btb_bht_T : btb_108_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5229 = 9'h6d == btb_victim_ptr ? _btb_bht_T : btb_109_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5230 = 9'h6e == btb_victim_ptr ? _btb_bht_T : btb_110_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5231 = 9'h6f == btb_victim_ptr ? _btb_bht_T : btb_111_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5232 = 9'h70 == btb_victim_ptr ? _btb_bht_T : btb_112_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5233 = 9'h71 == btb_victim_ptr ? _btb_bht_T : btb_113_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5234 = 9'h72 == btb_victim_ptr ? _btb_bht_T : btb_114_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5235 = 9'h73 == btb_victim_ptr ? _btb_bht_T : btb_115_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5236 = 9'h74 == btb_victim_ptr ? _btb_bht_T : btb_116_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5237 = 9'h75 == btb_victim_ptr ? _btb_bht_T : btb_117_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5238 = 9'h76 == btb_victim_ptr ? _btb_bht_T : btb_118_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5239 = 9'h77 == btb_victim_ptr ? _btb_bht_T : btb_119_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5240 = 9'h78 == btb_victim_ptr ? _btb_bht_T : btb_120_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5241 = 9'h79 == btb_victim_ptr ? _btb_bht_T : btb_121_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5242 = 9'h7a == btb_victim_ptr ? _btb_bht_T : btb_122_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5243 = 9'h7b == btb_victim_ptr ? _btb_bht_T : btb_123_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5244 = 9'h7c == btb_victim_ptr ? _btb_bht_T : btb_124_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5245 = 9'h7d == btb_victim_ptr ? _btb_bht_T : btb_125_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5246 = 9'h7e == btb_victim_ptr ? _btb_bht_T : btb_126_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5247 = 9'h7f == btb_victim_ptr ? _btb_bht_T : btb_127_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5248 = 9'h80 == btb_victim_ptr ? _btb_bht_T : btb_128_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5249 = 9'h81 == btb_victim_ptr ? _btb_bht_T : btb_129_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5250 = 9'h82 == btb_victim_ptr ? _btb_bht_T : btb_130_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5251 = 9'h83 == btb_victim_ptr ? _btb_bht_T : btb_131_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5252 = 9'h84 == btb_victim_ptr ? _btb_bht_T : btb_132_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5253 = 9'h85 == btb_victim_ptr ? _btb_bht_T : btb_133_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5254 = 9'h86 == btb_victim_ptr ? _btb_bht_T : btb_134_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5255 = 9'h87 == btb_victim_ptr ? _btb_bht_T : btb_135_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5256 = 9'h88 == btb_victim_ptr ? _btb_bht_T : btb_136_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5257 = 9'h89 == btb_victim_ptr ? _btb_bht_T : btb_137_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5258 = 9'h8a == btb_victim_ptr ? _btb_bht_T : btb_138_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5259 = 9'h8b == btb_victim_ptr ? _btb_bht_T : btb_139_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5260 = 9'h8c == btb_victim_ptr ? _btb_bht_T : btb_140_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5261 = 9'h8d == btb_victim_ptr ? _btb_bht_T : btb_141_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5262 = 9'h8e == btb_victim_ptr ? _btb_bht_T : btb_142_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5263 = 9'h8f == btb_victim_ptr ? _btb_bht_T : btb_143_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5264 = 9'h90 == btb_victim_ptr ? _btb_bht_T : btb_144_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5265 = 9'h91 == btb_victim_ptr ? _btb_bht_T : btb_145_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5266 = 9'h92 == btb_victim_ptr ? _btb_bht_T : btb_146_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5267 = 9'h93 == btb_victim_ptr ? _btb_bht_T : btb_147_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5268 = 9'h94 == btb_victim_ptr ? _btb_bht_T : btb_148_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5269 = 9'h95 == btb_victim_ptr ? _btb_bht_T : btb_149_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5270 = 9'h96 == btb_victim_ptr ? _btb_bht_T : btb_150_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5271 = 9'h97 == btb_victim_ptr ? _btb_bht_T : btb_151_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5272 = 9'h98 == btb_victim_ptr ? _btb_bht_T : btb_152_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5273 = 9'h99 == btb_victim_ptr ? _btb_bht_T : btb_153_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5274 = 9'h9a == btb_victim_ptr ? _btb_bht_T : btb_154_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5275 = 9'h9b == btb_victim_ptr ? _btb_bht_T : btb_155_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5276 = 9'h9c == btb_victim_ptr ? _btb_bht_T : btb_156_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5277 = 9'h9d == btb_victim_ptr ? _btb_bht_T : btb_157_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5278 = 9'h9e == btb_victim_ptr ? _btb_bht_T : btb_158_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5279 = 9'h9f == btb_victim_ptr ? _btb_bht_T : btb_159_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5280 = 9'ha0 == btb_victim_ptr ? _btb_bht_T : btb_160_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5281 = 9'ha1 == btb_victim_ptr ? _btb_bht_T : btb_161_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5282 = 9'ha2 == btb_victim_ptr ? _btb_bht_T : btb_162_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5283 = 9'ha3 == btb_victim_ptr ? _btb_bht_T : btb_163_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5284 = 9'ha4 == btb_victim_ptr ? _btb_bht_T : btb_164_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5285 = 9'ha5 == btb_victim_ptr ? _btb_bht_T : btb_165_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5286 = 9'ha6 == btb_victim_ptr ? _btb_bht_T : btb_166_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5287 = 9'ha7 == btb_victim_ptr ? _btb_bht_T : btb_167_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5288 = 9'ha8 == btb_victim_ptr ? _btb_bht_T : btb_168_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5289 = 9'ha9 == btb_victim_ptr ? _btb_bht_T : btb_169_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5290 = 9'haa == btb_victim_ptr ? _btb_bht_T : btb_170_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5291 = 9'hab == btb_victim_ptr ? _btb_bht_T : btb_171_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5292 = 9'hac == btb_victim_ptr ? _btb_bht_T : btb_172_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5293 = 9'had == btb_victim_ptr ? _btb_bht_T : btb_173_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5294 = 9'hae == btb_victim_ptr ? _btb_bht_T : btb_174_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5295 = 9'haf == btb_victim_ptr ? _btb_bht_T : btb_175_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5296 = 9'hb0 == btb_victim_ptr ? _btb_bht_T : btb_176_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5297 = 9'hb1 == btb_victim_ptr ? _btb_bht_T : btb_177_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5298 = 9'hb2 == btb_victim_ptr ? _btb_bht_T : btb_178_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5299 = 9'hb3 == btb_victim_ptr ? _btb_bht_T : btb_179_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5300 = 9'hb4 == btb_victim_ptr ? _btb_bht_T : btb_180_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5301 = 9'hb5 == btb_victim_ptr ? _btb_bht_T : btb_181_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5302 = 9'hb6 == btb_victim_ptr ? _btb_bht_T : btb_182_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5303 = 9'hb7 == btb_victim_ptr ? _btb_bht_T : btb_183_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5304 = 9'hb8 == btb_victim_ptr ? _btb_bht_T : btb_184_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5305 = 9'hb9 == btb_victim_ptr ? _btb_bht_T : btb_185_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5306 = 9'hba == btb_victim_ptr ? _btb_bht_T : btb_186_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5307 = 9'hbb == btb_victim_ptr ? _btb_bht_T : btb_187_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5308 = 9'hbc == btb_victim_ptr ? _btb_bht_T : btb_188_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5309 = 9'hbd == btb_victim_ptr ? _btb_bht_T : btb_189_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5310 = 9'hbe == btb_victim_ptr ? _btb_bht_T : btb_190_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5311 = 9'hbf == btb_victim_ptr ? _btb_bht_T : btb_191_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5312 = 9'hc0 == btb_victim_ptr ? _btb_bht_T : btb_192_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5313 = 9'hc1 == btb_victim_ptr ? _btb_bht_T : btb_193_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5314 = 9'hc2 == btb_victim_ptr ? _btb_bht_T : btb_194_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5315 = 9'hc3 == btb_victim_ptr ? _btb_bht_T : btb_195_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5316 = 9'hc4 == btb_victim_ptr ? _btb_bht_T : btb_196_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5317 = 9'hc5 == btb_victim_ptr ? _btb_bht_T : btb_197_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5318 = 9'hc6 == btb_victim_ptr ? _btb_bht_T : btb_198_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5319 = 9'hc7 == btb_victim_ptr ? _btb_bht_T : btb_199_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5320 = 9'hc8 == btb_victim_ptr ? _btb_bht_T : btb_200_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5321 = 9'hc9 == btb_victim_ptr ? _btb_bht_T : btb_201_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5322 = 9'hca == btb_victim_ptr ? _btb_bht_T : btb_202_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5323 = 9'hcb == btb_victim_ptr ? _btb_bht_T : btb_203_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5324 = 9'hcc == btb_victim_ptr ? _btb_bht_T : btb_204_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5325 = 9'hcd == btb_victim_ptr ? _btb_bht_T : btb_205_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5326 = 9'hce == btb_victim_ptr ? _btb_bht_T : btb_206_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5327 = 9'hcf == btb_victim_ptr ? _btb_bht_T : btb_207_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5328 = 9'hd0 == btb_victim_ptr ? _btb_bht_T : btb_208_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5329 = 9'hd1 == btb_victim_ptr ? _btb_bht_T : btb_209_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5330 = 9'hd2 == btb_victim_ptr ? _btb_bht_T : btb_210_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5331 = 9'hd3 == btb_victim_ptr ? _btb_bht_T : btb_211_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5332 = 9'hd4 == btb_victim_ptr ? _btb_bht_T : btb_212_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5333 = 9'hd5 == btb_victim_ptr ? _btb_bht_T : btb_213_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5334 = 9'hd6 == btb_victim_ptr ? _btb_bht_T : btb_214_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5335 = 9'hd7 == btb_victim_ptr ? _btb_bht_T : btb_215_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5336 = 9'hd8 == btb_victim_ptr ? _btb_bht_T : btb_216_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5337 = 9'hd9 == btb_victim_ptr ? _btb_bht_T : btb_217_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5338 = 9'hda == btb_victim_ptr ? _btb_bht_T : btb_218_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5339 = 9'hdb == btb_victim_ptr ? _btb_bht_T : btb_219_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5340 = 9'hdc == btb_victim_ptr ? _btb_bht_T : btb_220_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5341 = 9'hdd == btb_victim_ptr ? _btb_bht_T : btb_221_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5342 = 9'hde == btb_victim_ptr ? _btb_bht_T : btb_222_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5343 = 9'hdf == btb_victim_ptr ? _btb_bht_T : btb_223_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5344 = 9'he0 == btb_victim_ptr ? _btb_bht_T : btb_224_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5345 = 9'he1 == btb_victim_ptr ? _btb_bht_T : btb_225_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5346 = 9'he2 == btb_victim_ptr ? _btb_bht_T : btb_226_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5347 = 9'he3 == btb_victim_ptr ? _btb_bht_T : btb_227_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5348 = 9'he4 == btb_victim_ptr ? _btb_bht_T : btb_228_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5349 = 9'he5 == btb_victim_ptr ? _btb_bht_T : btb_229_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5350 = 9'he6 == btb_victim_ptr ? _btb_bht_T : btb_230_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5351 = 9'he7 == btb_victim_ptr ? _btb_bht_T : btb_231_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5352 = 9'he8 == btb_victim_ptr ? _btb_bht_T : btb_232_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5353 = 9'he9 == btb_victim_ptr ? _btb_bht_T : btb_233_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5354 = 9'hea == btb_victim_ptr ? _btb_bht_T : btb_234_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5355 = 9'heb == btb_victim_ptr ? _btb_bht_T : btb_235_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5356 = 9'hec == btb_victim_ptr ? _btb_bht_T : btb_236_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5357 = 9'hed == btb_victim_ptr ? _btb_bht_T : btb_237_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5358 = 9'hee == btb_victim_ptr ? _btb_bht_T : btb_238_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5359 = 9'hef == btb_victim_ptr ? _btb_bht_T : btb_239_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5360 = 9'hf0 == btb_victim_ptr ? _btb_bht_T : btb_240_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5361 = 9'hf1 == btb_victim_ptr ? _btb_bht_T : btb_241_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5362 = 9'hf2 == btb_victim_ptr ? _btb_bht_T : btb_242_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5363 = 9'hf3 == btb_victim_ptr ? _btb_bht_T : btb_243_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5364 = 9'hf4 == btb_victim_ptr ? _btb_bht_T : btb_244_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5365 = 9'hf5 == btb_victim_ptr ? _btb_bht_T : btb_245_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5366 = 9'hf6 == btb_victim_ptr ? _btb_bht_T : btb_246_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5367 = 9'hf7 == btb_victim_ptr ? _btb_bht_T : btb_247_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5368 = 9'hf8 == btb_victim_ptr ? _btb_bht_T : btb_248_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5369 = 9'hf9 == btb_victim_ptr ? _btb_bht_T : btb_249_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5370 = 9'hfa == btb_victim_ptr ? _btb_bht_T : btb_250_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5371 = 9'hfb == btb_victim_ptr ? _btb_bht_T : btb_251_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5372 = 9'hfc == btb_victim_ptr ? _btb_bht_T : btb_252_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5373 = 9'hfd == btb_victim_ptr ? _btb_bht_T : btb_253_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5374 = 9'hfe == btb_victim_ptr ? _btb_bht_T : btb_254_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5375 = 9'hff == btb_victim_ptr ? _btb_bht_T : btb_255_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5376 = 9'h100 == btb_victim_ptr ? _btb_bht_T : btb_256_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5377 = 9'h101 == btb_victim_ptr ? _btb_bht_T : btb_257_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5378 = 9'h102 == btb_victim_ptr ? _btb_bht_T : btb_258_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5379 = 9'h103 == btb_victim_ptr ? _btb_bht_T : btb_259_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5380 = 9'h104 == btb_victim_ptr ? _btb_bht_T : btb_260_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5381 = 9'h105 == btb_victim_ptr ? _btb_bht_T : btb_261_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5382 = 9'h106 == btb_victim_ptr ? _btb_bht_T : btb_262_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5383 = 9'h107 == btb_victim_ptr ? _btb_bht_T : btb_263_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5384 = 9'h108 == btb_victim_ptr ? _btb_bht_T : btb_264_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5385 = 9'h109 == btb_victim_ptr ? _btb_bht_T : btb_265_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5386 = 9'h10a == btb_victim_ptr ? _btb_bht_T : btb_266_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5387 = 9'h10b == btb_victim_ptr ? _btb_bht_T : btb_267_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5388 = 9'h10c == btb_victim_ptr ? _btb_bht_T : btb_268_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5389 = 9'h10d == btb_victim_ptr ? _btb_bht_T : btb_269_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5390 = 9'h10e == btb_victim_ptr ? _btb_bht_T : btb_270_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5391 = 9'h10f == btb_victim_ptr ? _btb_bht_T : btb_271_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5392 = 9'h110 == btb_victim_ptr ? _btb_bht_T : btb_272_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5393 = 9'h111 == btb_victim_ptr ? _btb_bht_T : btb_273_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5394 = 9'h112 == btb_victim_ptr ? _btb_bht_T : btb_274_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5395 = 9'h113 == btb_victim_ptr ? _btb_bht_T : btb_275_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5396 = 9'h114 == btb_victim_ptr ? _btb_bht_T : btb_276_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5397 = 9'h115 == btb_victim_ptr ? _btb_bht_T : btb_277_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5398 = 9'h116 == btb_victim_ptr ? _btb_bht_T : btb_278_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5399 = 9'h117 == btb_victim_ptr ? _btb_bht_T : btb_279_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5400 = 9'h118 == btb_victim_ptr ? _btb_bht_T : btb_280_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5401 = 9'h119 == btb_victim_ptr ? _btb_bht_T : btb_281_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5402 = 9'h11a == btb_victim_ptr ? _btb_bht_T : btb_282_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5403 = 9'h11b == btb_victim_ptr ? _btb_bht_T : btb_283_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5404 = 9'h11c == btb_victim_ptr ? _btb_bht_T : btb_284_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5405 = 9'h11d == btb_victim_ptr ? _btb_bht_T : btb_285_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5406 = 9'h11e == btb_victim_ptr ? _btb_bht_T : btb_286_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5407 = 9'h11f == btb_victim_ptr ? _btb_bht_T : btb_287_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5408 = 9'h120 == btb_victim_ptr ? _btb_bht_T : btb_288_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5409 = 9'h121 == btb_victim_ptr ? _btb_bht_T : btb_289_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5410 = 9'h122 == btb_victim_ptr ? _btb_bht_T : btb_290_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5411 = 9'h123 == btb_victim_ptr ? _btb_bht_T : btb_291_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5412 = 9'h124 == btb_victim_ptr ? _btb_bht_T : btb_292_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5413 = 9'h125 == btb_victim_ptr ? _btb_bht_T : btb_293_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5414 = 9'h126 == btb_victim_ptr ? _btb_bht_T : btb_294_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5415 = 9'h127 == btb_victim_ptr ? _btb_bht_T : btb_295_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5416 = 9'h128 == btb_victim_ptr ? _btb_bht_T : btb_296_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5417 = 9'h129 == btb_victim_ptr ? _btb_bht_T : btb_297_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5418 = 9'h12a == btb_victim_ptr ? _btb_bht_T : btb_298_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5419 = 9'h12b == btb_victim_ptr ? _btb_bht_T : btb_299_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5420 = 9'h12c == btb_victim_ptr ? _btb_bht_T : btb_300_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5421 = 9'h12d == btb_victim_ptr ? _btb_bht_T : btb_301_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5422 = 9'h12e == btb_victim_ptr ? _btb_bht_T : btb_302_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5423 = 9'h12f == btb_victim_ptr ? _btb_bht_T : btb_303_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5424 = 9'h130 == btb_victim_ptr ? _btb_bht_T : btb_304_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5425 = 9'h131 == btb_victim_ptr ? _btb_bht_T : btb_305_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5426 = 9'h132 == btb_victim_ptr ? _btb_bht_T : btb_306_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5427 = 9'h133 == btb_victim_ptr ? _btb_bht_T : btb_307_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5428 = 9'h134 == btb_victim_ptr ? _btb_bht_T : btb_308_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5429 = 9'h135 == btb_victim_ptr ? _btb_bht_T : btb_309_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5430 = 9'h136 == btb_victim_ptr ? _btb_bht_T : btb_310_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5431 = 9'h137 == btb_victim_ptr ? _btb_bht_T : btb_311_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5432 = 9'h138 == btb_victim_ptr ? _btb_bht_T : btb_312_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5433 = 9'h139 == btb_victim_ptr ? _btb_bht_T : btb_313_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5434 = 9'h13a == btb_victim_ptr ? _btb_bht_T : btb_314_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5435 = 9'h13b == btb_victim_ptr ? _btb_bht_T : btb_315_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5436 = 9'h13c == btb_victim_ptr ? _btb_bht_T : btb_316_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5437 = 9'h13d == btb_victim_ptr ? _btb_bht_T : btb_317_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5438 = 9'h13e == btb_victim_ptr ? _btb_bht_T : btb_318_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5439 = 9'h13f == btb_victim_ptr ? _btb_bht_T : btb_319_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5440 = 9'h140 == btb_victim_ptr ? _btb_bht_T : btb_320_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5441 = 9'h141 == btb_victim_ptr ? _btb_bht_T : btb_321_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5442 = 9'h142 == btb_victim_ptr ? _btb_bht_T : btb_322_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5443 = 9'h143 == btb_victim_ptr ? _btb_bht_T : btb_323_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5444 = 9'h144 == btb_victim_ptr ? _btb_bht_T : btb_324_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5445 = 9'h145 == btb_victim_ptr ? _btb_bht_T : btb_325_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5446 = 9'h146 == btb_victim_ptr ? _btb_bht_T : btb_326_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5447 = 9'h147 == btb_victim_ptr ? _btb_bht_T : btb_327_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5448 = 9'h148 == btb_victim_ptr ? _btb_bht_T : btb_328_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5449 = 9'h149 == btb_victim_ptr ? _btb_bht_T : btb_329_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5450 = 9'h14a == btb_victim_ptr ? _btb_bht_T : btb_330_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5451 = 9'h14b == btb_victim_ptr ? _btb_bht_T : btb_331_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5452 = 9'h14c == btb_victim_ptr ? _btb_bht_T : btb_332_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5453 = 9'h14d == btb_victim_ptr ? _btb_bht_T : btb_333_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5454 = 9'h14e == btb_victim_ptr ? _btb_bht_T : btb_334_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5455 = 9'h14f == btb_victim_ptr ? _btb_bht_T : btb_335_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5456 = 9'h150 == btb_victim_ptr ? _btb_bht_T : btb_336_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5457 = 9'h151 == btb_victim_ptr ? _btb_bht_T : btb_337_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5458 = 9'h152 == btb_victim_ptr ? _btb_bht_T : btb_338_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5459 = 9'h153 == btb_victim_ptr ? _btb_bht_T : btb_339_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5460 = 9'h154 == btb_victim_ptr ? _btb_bht_T : btb_340_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5461 = 9'h155 == btb_victim_ptr ? _btb_bht_T : btb_341_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5462 = 9'h156 == btb_victim_ptr ? _btb_bht_T : btb_342_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5463 = 9'h157 == btb_victim_ptr ? _btb_bht_T : btb_343_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5464 = 9'h158 == btb_victim_ptr ? _btb_bht_T : btb_344_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5465 = 9'h159 == btb_victim_ptr ? _btb_bht_T : btb_345_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5466 = 9'h15a == btb_victim_ptr ? _btb_bht_T : btb_346_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5467 = 9'h15b == btb_victim_ptr ? _btb_bht_T : btb_347_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5468 = 9'h15c == btb_victim_ptr ? _btb_bht_T : btb_348_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5469 = 9'h15d == btb_victim_ptr ? _btb_bht_T : btb_349_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5470 = 9'h15e == btb_victim_ptr ? _btb_bht_T : btb_350_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5471 = 9'h15f == btb_victim_ptr ? _btb_bht_T : btb_351_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5472 = 9'h160 == btb_victim_ptr ? _btb_bht_T : btb_352_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5473 = 9'h161 == btb_victim_ptr ? _btb_bht_T : btb_353_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5474 = 9'h162 == btb_victim_ptr ? _btb_bht_T : btb_354_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5475 = 9'h163 == btb_victim_ptr ? _btb_bht_T : btb_355_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5476 = 9'h164 == btb_victim_ptr ? _btb_bht_T : btb_356_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5477 = 9'h165 == btb_victim_ptr ? _btb_bht_T : btb_357_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5478 = 9'h166 == btb_victim_ptr ? _btb_bht_T : btb_358_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5479 = 9'h167 == btb_victim_ptr ? _btb_bht_T : btb_359_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5480 = 9'h168 == btb_victim_ptr ? _btb_bht_T : btb_360_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5481 = 9'h169 == btb_victim_ptr ? _btb_bht_T : btb_361_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5482 = 9'h16a == btb_victim_ptr ? _btb_bht_T : btb_362_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5483 = 9'h16b == btb_victim_ptr ? _btb_bht_T : btb_363_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5484 = 9'h16c == btb_victim_ptr ? _btb_bht_T : btb_364_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5485 = 9'h16d == btb_victim_ptr ? _btb_bht_T : btb_365_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5486 = 9'h16e == btb_victim_ptr ? _btb_bht_T : btb_366_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5487 = 9'h16f == btb_victim_ptr ? _btb_bht_T : btb_367_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5488 = 9'h170 == btb_victim_ptr ? _btb_bht_T : btb_368_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5489 = 9'h171 == btb_victim_ptr ? _btb_bht_T : btb_369_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5490 = 9'h172 == btb_victim_ptr ? _btb_bht_T : btb_370_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5491 = 9'h173 == btb_victim_ptr ? _btb_bht_T : btb_371_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5492 = 9'h174 == btb_victim_ptr ? _btb_bht_T : btb_372_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5493 = 9'h175 == btb_victim_ptr ? _btb_bht_T : btb_373_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5494 = 9'h176 == btb_victim_ptr ? _btb_bht_T : btb_374_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5495 = 9'h177 == btb_victim_ptr ? _btb_bht_T : btb_375_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5496 = 9'h178 == btb_victim_ptr ? _btb_bht_T : btb_376_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5497 = 9'h179 == btb_victim_ptr ? _btb_bht_T : btb_377_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5498 = 9'h17a == btb_victim_ptr ? _btb_bht_T : btb_378_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5499 = 9'h17b == btb_victim_ptr ? _btb_bht_T : btb_379_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5500 = 9'h17c == btb_victim_ptr ? _btb_bht_T : btb_380_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5501 = 9'h17d == btb_victim_ptr ? _btb_bht_T : btb_381_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5502 = 9'h17e == btb_victim_ptr ? _btb_bht_T : btb_382_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5503 = 9'h17f == btb_victim_ptr ? _btb_bht_T : btb_383_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5504 = 9'h180 == btb_victim_ptr ? _btb_bht_T : btb_384_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5505 = 9'h181 == btb_victim_ptr ? _btb_bht_T : btb_385_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5506 = 9'h182 == btb_victim_ptr ? _btb_bht_T : btb_386_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5507 = 9'h183 == btb_victim_ptr ? _btb_bht_T : btb_387_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5508 = 9'h184 == btb_victim_ptr ? _btb_bht_T : btb_388_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5509 = 9'h185 == btb_victim_ptr ? _btb_bht_T : btb_389_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5510 = 9'h186 == btb_victim_ptr ? _btb_bht_T : btb_390_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5511 = 9'h187 == btb_victim_ptr ? _btb_bht_T : btb_391_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5512 = 9'h188 == btb_victim_ptr ? _btb_bht_T : btb_392_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5513 = 9'h189 == btb_victim_ptr ? _btb_bht_T : btb_393_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5514 = 9'h18a == btb_victim_ptr ? _btb_bht_T : btb_394_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5515 = 9'h18b == btb_victim_ptr ? _btb_bht_T : btb_395_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5516 = 9'h18c == btb_victim_ptr ? _btb_bht_T : btb_396_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5517 = 9'h18d == btb_victim_ptr ? _btb_bht_T : btb_397_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5518 = 9'h18e == btb_victim_ptr ? _btb_bht_T : btb_398_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5519 = 9'h18f == btb_victim_ptr ? _btb_bht_T : btb_399_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5520 = 9'h190 == btb_victim_ptr ? _btb_bht_T : btb_400_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5521 = 9'h191 == btb_victim_ptr ? _btb_bht_T : btb_401_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5522 = 9'h192 == btb_victim_ptr ? _btb_bht_T : btb_402_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5523 = 9'h193 == btb_victim_ptr ? _btb_bht_T : btb_403_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5524 = 9'h194 == btb_victim_ptr ? _btb_bht_T : btb_404_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5525 = 9'h195 == btb_victim_ptr ? _btb_bht_T : btb_405_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5526 = 9'h196 == btb_victim_ptr ? _btb_bht_T : btb_406_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5527 = 9'h197 == btb_victim_ptr ? _btb_bht_T : btb_407_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5528 = 9'h198 == btb_victim_ptr ? _btb_bht_T : btb_408_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5529 = 9'h199 == btb_victim_ptr ? _btb_bht_T : btb_409_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5530 = 9'h19a == btb_victim_ptr ? _btb_bht_T : btb_410_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5531 = 9'h19b == btb_victim_ptr ? _btb_bht_T : btb_411_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5532 = 9'h19c == btb_victim_ptr ? _btb_bht_T : btb_412_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5533 = 9'h19d == btb_victim_ptr ? _btb_bht_T : btb_413_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5534 = 9'h19e == btb_victim_ptr ? _btb_bht_T : btb_414_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5535 = 9'h19f == btb_victim_ptr ? _btb_bht_T : btb_415_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5536 = 9'h1a0 == btb_victim_ptr ? _btb_bht_T : btb_416_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5537 = 9'h1a1 == btb_victim_ptr ? _btb_bht_T : btb_417_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5538 = 9'h1a2 == btb_victim_ptr ? _btb_bht_T : btb_418_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5539 = 9'h1a3 == btb_victim_ptr ? _btb_bht_T : btb_419_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5540 = 9'h1a4 == btb_victim_ptr ? _btb_bht_T : btb_420_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5541 = 9'h1a5 == btb_victim_ptr ? _btb_bht_T : btb_421_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5542 = 9'h1a6 == btb_victim_ptr ? _btb_bht_T : btb_422_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5543 = 9'h1a7 == btb_victim_ptr ? _btb_bht_T : btb_423_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5544 = 9'h1a8 == btb_victim_ptr ? _btb_bht_T : btb_424_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5545 = 9'h1a9 == btb_victim_ptr ? _btb_bht_T : btb_425_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5546 = 9'h1aa == btb_victim_ptr ? _btb_bht_T : btb_426_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5547 = 9'h1ab == btb_victim_ptr ? _btb_bht_T : btb_427_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5548 = 9'h1ac == btb_victim_ptr ? _btb_bht_T : btb_428_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5549 = 9'h1ad == btb_victim_ptr ? _btb_bht_T : btb_429_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5550 = 9'h1ae == btb_victim_ptr ? _btb_bht_T : btb_430_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5551 = 9'h1af == btb_victim_ptr ? _btb_bht_T : btb_431_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5552 = 9'h1b0 == btb_victim_ptr ? _btb_bht_T : btb_432_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5553 = 9'h1b1 == btb_victim_ptr ? _btb_bht_T : btb_433_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5554 = 9'h1b2 == btb_victim_ptr ? _btb_bht_T : btb_434_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5555 = 9'h1b3 == btb_victim_ptr ? _btb_bht_T : btb_435_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5556 = 9'h1b4 == btb_victim_ptr ? _btb_bht_T : btb_436_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5557 = 9'h1b5 == btb_victim_ptr ? _btb_bht_T : btb_437_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5558 = 9'h1b6 == btb_victim_ptr ? _btb_bht_T : btb_438_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5559 = 9'h1b7 == btb_victim_ptr ? _btb_bht_T : btb_439_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5560 = 9'h1b8 == btb_victim_ptr ? _btb_bht_T : btb_440_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5561 = 9'h1b9 == btb_victim_ptr ? _btb_bht_T : btb_441_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5562 = 9'h1ba == btb_victim_ptr ? _btb_bht_T : btb_442_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5563 = 9'h1bb == btb_victim_ptr ? _btb_bht_T : btb_443_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5564 = 9'h1bc == btb_victim_ptr ? _btb_bht_T : btb_444_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5565 = 9'h1bd == btb_victim_ptr ? _btb_bht_T : btb_445_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5566 = 9'h1be == btb_victim_ptr ? _btb_bht_T : btb_446_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5567 = 9'h1bf == btb_victim_ptr ? _btb_bht_T : btb_447_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5568 = 9'h1c0 == btb_victim_ptr ? _btb_bht_T : btb_448_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5569 = 9'h1c1 == btb_victim_ptr ? _btb_bht_T : btb_449_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5570 = 9'h1c2 == btb_victim_ptr ? _btb_bht_T : btb_450_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5571 = 9'h1c3 == btb_victim_ptr ? _btb_bht_T : btb_451_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5572 = 9'h1c4 == btb_victim_ptr ? _btb_bht_T : btb_452_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5573 = 9'h1c5 == btb_victim_ptr ? _btb_bht_T : btb_453_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5574 = 9'h1c6 == btb_victim_ptr ? _btb_bht_T : btb_454_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5575 = 9'h1c7 == btb_victim_ptr ? _btb_bht_T : btb_455_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5576 = 9'h1c8 == btb_victim_ptr ? _btb_bht_T : btb_456_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5577 = 9'h1c9 == btb_victim_ptr ? _btb_bht_T : btb_457_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5578 = 9'h1ca == btb_victim_ptr ? _btb_bht_T : btb_458_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5579 = 9'h1cb == btb_victim_ptr ? _btb_bht_T : btb_459_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5580 = 9'h1cc == btb_victim_ptr ? _btb_bht_T : btb_460_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5581 = 9'h1cd == btb_victim_ptr ? _btb_bht_T : btb_461_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5582 = 9'h1ce == btb_victim_ptr ? _btb_bht_T : btb_462_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5583 = 9'h1cf == btb_victim_ptr ? _btb_bht_T : btb_463_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5584 = 9'h1d0 == btb_victim_ptr ? _btb_bht_T : btb_464_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5585 = 9'h1d1 == btb_victim_ptr ? _btb_bht_T : btb_465_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5586 = 9'h1d2 == btb_victim_ptr ? _btb_bht_T : btb_466_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5587 = 9'h1d3 == btb_victim_ptr ? _btb_bht_T : btb_467_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5588 = 9'h1d4 == btb_victim_ptr ? _btb_bht_T : btb_468_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5589 = 9'h1d5 == btb_victim_ptr ? _btb_bht_T : btb_469_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5590 = 9'h1d6 == btb_victim_ptr ? _btb_bht_T : btb_470_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5591 = 9'h1d7 == btb_victim_ptr ? _btb_bht_T : btb_471_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5592 = 9'h1d8 == btb_victim_ptr ? _btb_bht_T : btb_472_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5593 = 9'h1d9 == btb_victim_ptr ? _btb_bht_T : btb_473_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5594 = 9'h1da == btb_victim_ptr ? _btb_bht_T : btb_474_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5595 = 9'h1db == btb_victim_ptr ? _btb_bht_T : btb_475_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5596 = 9'h1dc == btb_victim_ptr ? _btb_bht_T : btb_476_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5597 = 9'h1dd == btb_victim_ptr ? _btb_bht_T : btb_477_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5598 = 9'h1de == btb_victim_ptr ? _btb_bht_T : btb_478_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5599 = 9'h1df == btb_victim_ptr ? _btb_bht_T : btb_479_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5600 = 9'h1e0 == btb_victim_ptr ? _btb_bht_T : btb_480_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5601 = 9'h1e1 == btb_victim_ptr ? _btb_bht_T : btb_481_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5602 = 9'h1e2 == btb_victim_ptr ? _btb_bht_T : btb_482_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5603 = 9'h1e3 == btb_victim_ptr ? _btb_bht_T : btb_483_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5604 = 9'h1e4 == btb_victim_ptr ? _btb_bht_T : btb_484_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5605 = 9'h1e5 == btb_victim_ptr ? _btb_bht_T : btb_485_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5606 = 9'h1e6 == btb_victim_ptr ? _btb_bht_T : btb_486_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5607 = 9'h1e7 == btb_victim_ptr ? _btb_bht_T : btb_487_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5608 = 9'h1e8 == btb_victim_ptr ? _btb_bht_T : btb_488_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5609 = 9'h1e9 == btb_victim_ptr ? _btb_bht_T : btb_489_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5610 = 9'h1ea == btb_victim_ptr ? _btb_bht_T : btb_490_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5611 = 9'h1eb == btb_victim_ptr ? _btb_bht_T : btb_491_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5612 = 9'h1ec == btb_victim_ptr ? _btb_bht_T : btb_492_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5613 = 9'h1ed == btb_victim_ptr ? _btb_bht_T : btb_493_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5614 = 9'h1ee == btb_victim_ptr ? _btb_bht_T : btb_494_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5615 = 9'h1ef == btb_victim_ptr ? _btb_bht_T : btb_495_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5616 = 9'h1f0 == btb_victim_ptr ? _btb_bht_T : btb_496_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5617 = 9'h1f1 == btb_victim_ptr ? _btb_bht_T : btb_497_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5618 = 9'h1f2 == btb_victim_ptr ? _btb_bht_T : btb_498_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5619 = 9'h1f3 == btb_victim_ptr ? _btb_bht_T : btb_499_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5620 = 9'h1f4 == btb_victim_ptr ? _btb_bht_T : btb_500_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5621 = 9'h1f5 == btb_victim_ptr ? _btb_bht_T : btb_501_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5622 = 9'h1f6 == btb_victim_ptr ? _btb_bht_T : btb_502_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5623 = 9'h1f7 == btb_victim_ptr ? _btb_bht_T : btb_503_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5624 = 9'h1f8 == btb_victim_ptr ? _btb_bht_T : btb_504_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5625 = 9'h1f9 == btb_victim_ptr ? _btb_bht_T : btb_505_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5626 = 9'h1fa == btb_victim_ptr ? _btb_bht_T : btb_506_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5627 = 9'h1fb == btb_victim_ptr ? _btb_bht_T : btb_507_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5628 = 9'h1fc == btb_victim_ptr ? _btb_bht_T : btb_508_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5629 = 9'h1fd == btb_victim_ptr ? _btb_bht_T : btb_509_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5630 = 9'h1fe == btb_victim_ptr ? _btb_bht_T : btb_510_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [1:0] _GEN_5631 = 9'h1ff == btb_victim_ptr ? _btb_bht_T : btb_511_bht; // @[branch_predictor.scala 30:22 68:{33,33}]
  wire [8:0] _btb_victim_ptr_T_1 = btb_victim_ptr + 9'h1; // @[branch_predictor.scala 71:42]
  wire  _GEN_5632 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2560 : btb_0_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5633 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2561 : btb_1_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5634 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2562 : btb_2_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5635 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2563 : btb_3_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5636 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2564 : btb_4_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5637 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2565 : btb_5_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5638 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2566 : btb_6_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5639 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2567 : btb_7_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5640 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2568 : btb_8_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5641 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2569 : btb_9_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5642 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2570 : btb_10_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5643 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2571 : btb_11_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5644 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2572 : btb_12_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5645 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2573 : btb_13_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5646 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2574 : btb_14_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5647 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2575 : btb_15_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5648 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2576 : btb_16_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5649 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2577 : btb_17_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5650 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2578 : btb_18_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5651 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2579 : btb_19_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5652 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2580 : btb_20_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5653 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2581 : btb_21_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5654 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2582 : btb_22_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5655 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2583 : btb_23_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5656 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2584 : btb_24_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5657 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2585 : btb_25_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5658 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2586 : btb_26_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5659 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2587 : btb_27_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5660 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2588 : btb_28_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5661 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2589 : btb_29_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5662 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2590 : btb_30_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5663 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2591 : btb_31_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5664 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2592 : btb_32_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5665 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2593 : btb_33_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5666 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2594 : btb_34_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5667 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2595 : btb_35_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5668 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2596 : btb_36_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5669 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2597 : btb_37_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5670 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2598 : btb_38_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5671 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2599 : btb_39_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5672 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2600 : btb_40_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5673 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2601 : btb_41_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5674 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2602 : btb_42_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5675 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2603 : btb_43_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5676 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2604 : btb_44_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5677 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2605 : btb_45_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5678 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2606 : btb_46_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5679 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2607 : btb_47_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5680 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2608 : btb_48_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5681 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2609 : btb_49_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5682 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2610 : btb_50_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5683 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2611 : btb_51_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5684 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2612 : btb_52_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5685 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2613 : btb_53_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5686 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2614 : btb_54_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5687 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2615 : btb_55_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5688 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2616 : btb_56_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5689 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2617 : btb_57_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5690 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2618 : btb_58_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5691 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2619 : btb_59_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5692 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2620 : btb_60_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5693 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2621 : btb_61_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5694 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2622 : btb_62_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5695 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2623 : btb_63_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5696 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2624 : btb_64_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5697 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2625 : btb_65_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5698 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2626 : btb_66_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5699 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2627 : btb_67_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5700 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2628 : btb_68_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5701 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2629 : btb_69_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5702 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2630 : btb_70_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5703 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2631 : btb_71_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5704 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2632 : btb_72_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5705 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2633 : btb_73_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5706 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2634 : btb_74_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5707 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2635 : btb_75_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5708 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2636 : btb_76_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5709 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2637 : btb_77_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5710 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2638 : btb_78_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5711 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2639 : btb_79_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5712 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2640 : btb_80_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5713 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2641 : btb_81_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5714 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2642 : btb_82_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5715 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2643 : btb_83_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5716 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2644 : btb_84_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5717 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2645 : btb_85_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5718 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2646 : btb_86_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5719 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2647 : btb_87_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5720 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2648 : btb_88_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5721 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2649 : btb_89_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5722 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2650 : btb_90_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5723 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2651 : btb_91_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5724 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2652 : btb_92_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5725 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2653 : btb_93_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5726 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2654 : btb_94_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5727 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2655 : btb_95_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5728 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2656 : btb_96_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5729 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2657 : btb_97_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5730 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2658 : btb_98_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5731 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2659 : btb_99_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5732 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2660 : btb_100_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5733 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2661 : btb_101_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5734 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2662 : btb_102_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5735 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2663 : btb_103_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5736 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2664 : btb_104_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5737 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2665 : btb_105_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5738 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2666 : btb_106_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5739 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2667 : btb_107_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5740 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2668 : btb_108_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5741 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2669 : btb_109_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5742 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2670 : btb_110_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5743 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2671 : btb_111_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5744 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2672 : btb_112_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5745 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2673 : btb_113_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5746 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2674 : btb_114_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5747 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2675 : btb_115_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5748 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2676 : btb_116_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5749 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2677 : btb_117_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5750 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2678 : btb_118_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5751 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2679 : btb_119_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5752 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2680 : btb_120_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5753 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2681 : btb_121_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5754 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2682 : btb_122_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5755 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2683 : btb_123_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5756 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2684 : btb_124_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5757 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2685 : btb_125_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5758 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2686 : btb_126_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5759 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2687 : btb_127_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5760 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2688 : btb_128_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5761 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2689 : btb_129_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5762 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2690 : btb_130_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5763 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2691 : btb_131_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5764 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2692 : btb_132_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5765 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2693 : btb_133_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5766 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2694 : btb_134_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5767 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2695 : btb_135_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5768 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2696 : btb_136_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5769 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2697 : btb_137_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5770 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2698 : btb_138_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5771 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2699 : btb_139_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5772 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2700 : btb_140_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5773 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2701 : btb_141_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5774 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2702 : btb_142_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5775 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2703 : btb_143_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5776 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2704 : btb_144_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5777 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2705 : btb_145_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5778 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2706 : btb_146_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5779 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2707 : btb_147_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5780 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2708 : btb_148_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5781 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2709 : btb_149_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5782 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2710 : btb_150_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5783 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2711 : btb_151_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5784 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2712 : btb_152_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5785 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2713 : btb_153_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5786 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2714 : btb_154_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5787 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2715 : btb_155_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5788 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2716 : btb_156_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5789 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2717 : btb_157_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5790 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2718 : btb_158_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5791 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2719 : btb_159_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5792 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2720 : btb_160_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5793 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2721 : btb_161_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5794 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2722 : btb_162_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5795 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2723 : btb_163_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5796 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2724 : btb_164_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5797 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2725 : btb_165_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5798 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2726 : btb_166_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5799 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2727 : btb_167_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5800 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2728 : btb_168_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5801 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2729 : btb_169_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5802 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2730 : btb_170_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5803 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2731 : btb_171_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5804 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2732 : btb_172_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5805 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2733 : btb_173_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5806 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2734 : btb_174_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5807 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2735 : btb_175_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5808 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2736 : btb_176_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5809 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2737 : btb_177_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5810 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2738 : btb_178_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5811 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2739 : btb_179_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5812 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2740 : btb_180_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5813 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2741 : btb_181_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5814 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2742 : btb_182_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5815 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2743 : btb_183_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5816 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2744 : btb_184_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5817 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2745 : btb_185_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5818 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2746 : btb_186_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5819 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2747 : btb_187_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5820 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2748 : btb_188_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5821 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2749 : btb_189_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5822 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2750 : btb_190_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5823 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2751 : btb_191_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5824 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2752 : btb_192_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5825 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2753 : btb_193_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5826 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2754 : btb_194_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5827 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2755 : btb_195_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5828 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2756 : btb_196_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5829 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2757 : btb_197_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5830 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2758 : btb_198_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5831 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2759 : btb_199_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5832 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2760 : btb_200_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5833 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2761 : btb_201_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5834 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2762 : btb_202_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5835 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2763 : btb_203_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5836 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2764 : btb_204_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5837 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2765 : btb_205_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5838 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2766 : btb_206_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5839 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2767 : btb_207_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5840 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2768 : btb_208_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5841 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2769 : btb_209_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5842 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2770 : btb_210_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5843 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2771 : btb_211_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5844 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2772 : btb_212_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5845 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2773 : btb_213_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5846 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2774 : btb_214_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5847 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2775 : btb_215_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5848 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2776 : btb_216_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5849 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2777 : btb_217_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5850 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2778 : btb_218_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5851 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2779 : btb_219_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5852 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2780 : btb_220_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5853 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2781 : btb_221_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5854 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2782 : btb_222_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5855 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2783 : btb_223_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5856 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2784 : btb_224_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5857 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2785 : btb_225_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5858 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2786 : btb_226_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5859 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2787 : btb_227_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5860 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2788 : btb_228_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5861 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2789 : btb_229_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5862 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2790 : btb_230_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5863 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2791 : btb_231_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5864 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2792 : btb_232_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5865 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2793 : btb_233_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5866 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2794 : btb_234_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5867 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2795 : btb_235_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5868 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2796 : btb_236_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5869 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2797 : btb_237_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5870 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2798 : btb_238_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5871 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2799 : btb_239_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5872 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2800 : btb_240_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5873 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2801 : btb_241_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5874 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2802 : btb_242_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5875 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2803 : btb_243_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5876 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2804 : btb_244_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5877 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2805 : btb_245_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5878 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2806 : btb_246_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5879 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2807 : btb_247_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5880 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2808 : btb_248_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5881 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2809 : btb_249_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5882 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2810 : btb_250_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5883 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2811 : btb_251_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5884 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2812 : btb_252_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5885 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2813 : btb_253_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5886 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2814 : btb_254_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5887 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2815 : btb_255_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5888 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2816 : btb_256_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5889 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2817 : btb_257_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5890 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2818 : btb_258_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5891 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2819 : btb_259_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5892 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2820 : btb_260_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5893 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2821 : btb_261_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5894 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2822 : btb_262_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5895 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2823 : btb_263_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5896 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2824 : btb_264_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5897 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2825 : btb_265_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5898 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2826 : btb_266_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5899 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2827 : btb_267_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5900 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2828 : btb_268_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5901 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2829 : btb_269_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5902 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2830 : btb_270_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5903 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2831 : btb_271_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5904 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2832 : btb_272_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5905 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2833 : btb_273_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5906 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2834 : btb_274_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5907 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2835 : btb_275_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5908 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2836 : btb_276_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5909 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2837 : btb_277_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5910 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2838 : btb_278_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5911 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2839 : btb_279_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5912 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2840 : btb_280_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5913 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2841 : btb_281_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5914 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2842 : btb_282_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5915 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2843 : btb_283_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5916 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2844 : btb_284_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5917 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2845 : btb_285_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5918 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2846 : btb_286_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5919 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2847 : btb_287_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5920 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2848 : btb_288_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5921 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2849 : btb_289_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5922 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2850 : btb_290_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5923 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2851 : btb_291_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5924 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2852 : btb_292_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5925 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2853 : btb_293_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5926 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2854 : btb_294_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5927 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2855 : btb_295_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5928 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2856 : btb_296_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5929 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2857 : btb_297_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5930 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2858 : btb_298_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5931 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2859 : btb_299_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5932 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2860 : btb_300_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5933 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2861 : btb_301_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5934 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2862 : btb_302_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5935 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2863 : btb_303_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5936 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2864 : btb_304_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5937 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2865 : btb_305_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5938 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2866 : btb_306_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5939 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2867 : btb_307_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5940 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2868 : btb_308_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5941 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2869 : btb_309_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5942 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2870 : btb_310_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5943 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2871 : btb_311_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5944 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2872 : btb_312_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5945 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2873 : btb_313_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5946 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2874 : btb_314_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5947 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2875 : btb_315_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5948 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2876 : btb_316_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5949 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2877 : btb_317_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5950 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2878 : btb_318_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5951 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2879 : btb_319_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5952 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2880 : btb_320_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5953 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2881 : btb_321_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5954 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2882 : btb_322_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5955 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2883 : btb_323_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5956 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2884 : btb_324_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5957 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2885 : btb_325_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5958 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2886 : btb_326_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5959 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2887 : btb_327_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5960 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2888 : btb_328_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5961 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2889 : btb_329_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5962 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2890 : btb_330_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5963 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2891 : btb_331_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5964 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2892 : btb_332_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5965 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2893 : btb_333_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5966 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2894 : btb_334_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5967 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2895 : btb_335_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5968 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2896 : btb_336_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5969 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2897 : btb_337_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5970 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2898 : btb_338_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5971 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2899 : btb_339_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5972 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2900 : btb_340_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5973 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2901 : btb_341_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5974 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2902 : btb_342_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5975 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2903 : btb_343_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5976 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2904 : btb_344_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5977 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2905 : btb_345_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5978 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2906 : btb_346_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5979 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2907 : btb_347_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5980 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2908 : btb_348_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5981 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2909 : btb_349_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5982 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2910 : btb_350_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5983 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2911 : btb_351_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5984 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2912 : btb_352_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5985 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2913 : btb_353_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5986 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2914 : btb_354_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5987 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2915 : btb_355_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5988 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2916 : btb_356_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5989 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2917 : btb_357_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5990 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2918 : btb_358_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5991 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2919 : btb_359_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5992 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2920 : btb_360_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5993 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2921 : btb_361_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5994 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2922 : btb_362_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5995 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2923 : btb_363_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5996 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2924 : btb_364_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5997 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2925 : btb_365_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5998 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2926 : btb_366_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_5999 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2927 : btb_367_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6000 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2928 : btb_368_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6001 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2929 : btb_369_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6002 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2930 : btb_370_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6003 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2931 : btb_371_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6004 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2932 : btb_372_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6005 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2933 : btb_373_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6006 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2934 : btb_374_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6007 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2935 : btb_375_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6008 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2936 : btb_376_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6009 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2937 : btb_377_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6010 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2938 : btb_378_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6011 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2939 : btb_379_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6012 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2940 : btb_380_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6013 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2941 : btb_381_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6014 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2942 : btb_382_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6015 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2943 : btb_383_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6016 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2944 : btb_384_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6017 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2945 : btb_385_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6018 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2946 : btb_386_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6019 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2947 : btb_387_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6020 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2948 : btb_388_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6021 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2949 : btb_389_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6022 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2950 : btb_390_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6023 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2951 : btb_391_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6024 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2952 : btb_392_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6025 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2953 : btb_393_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6026 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2954 : btb_394_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6027 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2955 : btb_395_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6028 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2956 : btb_396_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6029 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2957 : btb_397_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6030 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2958 : btb_398_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6031 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2959 : btb_399_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6032 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2960 : btb_400_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6033 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2961 : btb_401_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6034 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2962 : btb_402_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6035 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2963 : btb_403_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6036 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2964 : btb_404_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6037 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2965 : btb_405_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6038 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2966 : btb_406_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6039 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2967 : btb_407_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6040 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2968 : btb_408_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6041 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2969 : btb_409_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6042 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2970 : btb_410_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6043 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2971 : btb_411_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6044 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2972 : btb_412_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6045 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2973 : btb_413_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6046 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2974 : btb_414_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6047 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2975 : btb_415_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6048 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2976 : btb_416_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6049 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2977 : btb_417_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6050 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2978 : btb_418_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6051 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2979 : btb_419_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6052 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2980 : btb_420_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6053 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2981 : btb_421_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6054 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2982 : btb_422_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6055 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2983 : btb_423_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6056 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2984 : btb_424_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6057 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2985 : btb_425_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6058 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2986 : btb_426_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6059 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2987 : btb_427_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6060 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2988 : btb_428_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6061 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2989 : btb_429_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6062 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2990 : btb_430_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6063 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2991 : btb_431_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6064 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2992 : btb_432_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6065 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2993 : btb_433_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6066 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2994 : btb_434_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6067 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2995 : btb_435_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6068 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2996 : btb_436_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6069 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2997 : btb_437_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6070 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2998 : btb_438_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6071 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_2999 : btb_439_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6072 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3000 : btb_440_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6073 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3001 : btb_441_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6074 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3002 : btb_442_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6075 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3003 : btb_443_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6076 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3004 : btb_444_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6077 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3005 : btb_445_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6078 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3006 : btb_446_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6079 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3007 : btb_447_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6080 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3008 : btb_448_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6081 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3009 : btb_449_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6082 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3010 : btb_450_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6083 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3011 : btb_451_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6084 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3012 : btb_452_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6085 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3013 : btb_453_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6086 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3014 : btb_454_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6087 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3015 : btb_455_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6088 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3016 : btb_456_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6089 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3017 : btb_457_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6090 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3018 : btb_458_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6091 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3019 : btb_459_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6092 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3020 : btb_460_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6093 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3021 : btb_461_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6094 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3022 : btb_462_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6095 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3023 : btb_463_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6096 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3024 : btb_464_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6097 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3025 : btb_465_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6098 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3026 : btb_466_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6099 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3027 : btb_467_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6100 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3028 : btb_468_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6101 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3029 : btb_469_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6102 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3030 : btb_470_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6103 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3031 : btb_471_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6104 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3032 : btb_472_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6105 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3033 : btb_473_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6106 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3034 : btb_474_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6107 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3035 : btb_475_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6108 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3036 : btb_476_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6109 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3037 : btb_477_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6110 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3038 : btb_478_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6111 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3039 : btb_479_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6112 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3040 : btb_480_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6113 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3041 : btb_481_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6114 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3042 : btb_482_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6115 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3043 : btb_483_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6116 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3044 : btb_484_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6117 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3045 : btb_485_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6118 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3046 : btb_486_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6119 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3047 : btb_487_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6120 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3048 : btb_488_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6121 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3049 : btb_489_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6122 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3050 : btb_490_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6123 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3051 : btb_491_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6124 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3052 : btb_492_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6125 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3053 : btb_493_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6126 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3054 : btb_494_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6127 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3055 : btb_495_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6128 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3056 : btb_496_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6129 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3057 : btb_497_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6130 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3058 : btb_498_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6131 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3059 : btb_499_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6132 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3060 : btb_500_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6133 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3061 : btb_501_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6134 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3062 : btb_502_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6135 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3063 : btb_503_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6136 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3064 : btb_504_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6137 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3065 : btb_505_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6138 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3066 : btb_506_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6139 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3067 : btb_507_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6140 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3068 : btb_508_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6141 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3069 : btb_509_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6142 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3070 : btb_510_valid; // @[branch_predictor.scala 62:121 30:22]
  wire  _GEN_6143 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3071 : btb_511_valid; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6144 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3072 : btb_0_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6145 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3073 : btb_1_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6146 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3074 : btb_2_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6147 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3075 : btb_3_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6148 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3076 : btb_4_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6149 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3077 : btb_5_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6150 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3078 : btb_6_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6151 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3079 : btb_7_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6152 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3080 : btb_8_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6153 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3081 : btb_9_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6154 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3082 : btb_10_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6155 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3083 : btb_11_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6156 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3084 : btb_12_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6157 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3085 : btb_13_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6158 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3086 : btb_14_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6159 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3087 : btb_15_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6160 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3088 : btb_16_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6161 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3089 : btb_17_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6162 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3090 : btb_18_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6163 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3091 : btb_19_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6164 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3092 : btb_20_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6165 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3093 : btb_21_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6166 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3094 : btb_22_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6167 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3095 : btb_23_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6168 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3096 : btb_24_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6169 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3097 : btb_25_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6170 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3098 : btb_26_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6171 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3099 : btb_27_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6172 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3100 : btb_28_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6173 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3101 : btb_29_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6174 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3102 : btb_30_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6175 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3103 : btb_31_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6176 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3104 : btb_32_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6177 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3105 : btb_33_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6178 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3106 : btb_34_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6179 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3107 : btb_35_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6180 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3108 : btb_36_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6181 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3109 : btb_37_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6182 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3110 : btb_38_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6183 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3111 : btb_39_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6184 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3112 : btb_40_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6185 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3113 : btb_41_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6186 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3114 : btb_42_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6187 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3115 : btb_43_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6188 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3116 : btb_44_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6189 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3117 : btb_45_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6190 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3118 : btb_46_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6191 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3119 : btb_47_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6192 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3120 : btb_48_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6193 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3121 : btb_49_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6194 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3122 : btb_50_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6195 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3123 : btb_51_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6196 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3124 : btb_52_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6197 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3125 : btb_53_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6198 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3126 : btb_54_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6199 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3127 : btb_55_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6200 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3128 : btb_56_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6201 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3129 : btb_57_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6202 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3130 : btb_58_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6203 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3131 : btb_59_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6204 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3132 : btb_60_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6205 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3133 : btb_61_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6206 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3134 : btb_62_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6207 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3135 : btb_63_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6208 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3136 : btb_64_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6209 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3137 : btb_65_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6210 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3138 : btb_66_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6211 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3139 : btb_67_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6212 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3140 : btb_68_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6213 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3141 : btb_69_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6214 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3142 : btb_70_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6215 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3143 : btb_71_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6216 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3144 : btb_72_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6217 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3145 : btb_73_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6218 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3146 : btb_74_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6219 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3147 : btb_75_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6220 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3148 : btb_76_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6221 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3149 : btb_77_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6222 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3150 : btb_78_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6223 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3151 : btb_79_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6224 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3152 : btb_80_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6225 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3153 : btb_81_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6226 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3154 : btb_82_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6227 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3155 : btb_83_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6228 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3156 : btb_84_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6229 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3157 : btb_85_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6230 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3158 : btb_86_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6231 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3159 : btb_87_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6232 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3160 : btb_88_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6233 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3161 : btb_89_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6234 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3162 : btb_90_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6235 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3163 : btb_91_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6236 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3164 : btb_92_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6237 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3165 : btb_93_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6238 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3166 : btb_94_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6239 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3167 : btb_95_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6240 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3168 : btb_96_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6241 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3169 : btb_97_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6242 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3170 : btb_98_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6243 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3171 : btb_99_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6244 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3172 : btb_100_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6245 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3173 : btb_101_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6246 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3174 : btb_102_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6247 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3175 : btb_103_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6248 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3176 : btb_104_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6249 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3177 : btb_105_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6250 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3178 : btb_106_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6251 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3179 : btb_107_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6252 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3180 : btb_108_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6253 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3181 : btb_109_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6254 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3182 : btb_110_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6255 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3183 : btb_111_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6256 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3184 : btb_112_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6257 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3185 : btb_113_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6258 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3186 : btb_114_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6259 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3187 : btb_115_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6260 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3188 : btb_116_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6261 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3189 : btb_117_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6262 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3190 : btb_118_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6263 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3191 : btb_119_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6264 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3192 : btb_120_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6265 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3193 : btb_121_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6266 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3194 : btb_122_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6267 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3195 : btb_123_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6268 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3196 : btb_124_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6269 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3197 : btb_125_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6270 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3198 : btb_126_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6271 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3199 : btb_127_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6272 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3200 : btb_128_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6273 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3201 : btb_129_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6274 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3202 : btb_130_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6275 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3203 : btb_131_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6276 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3204 : btb_132_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6277 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3205 : btb_133_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6278 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3206 : btb_134_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6279 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3207 : btb_135_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6280 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3208 : btb_136_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6281 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3209 : btb_137_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6282 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3210 : btb_138_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6283 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3211 : btb_139_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6284 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3212 : btb_140_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6285 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3213 : btb_141_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6286 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3214 : btb_142_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6287 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3215 : btb_143_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6288 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3216 : btb_144_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6289 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3217 : btb_145_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6290 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3218 : btb_146_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6291 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3219 : btb_147_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6292 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3220 : btb_148_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6293 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3221 : btb_149_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6294 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3222 : btb_150_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6295 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3223 : btb_151_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6296 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3224 : btb_152_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6297 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3225 : btb_153_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6298 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3226 : btb_154_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6299 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3227 : btb_155_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6300 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3228 : btb_156_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6301 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3229 : btb_157_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6302 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3230 : btb_158_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6303 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3231 : btb_159_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6304 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3232 : btb_160_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6305 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3233 : btb_161_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6306 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3234 : btb_162_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6307 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3235 : btb_163_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6308 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3236 : btb_164_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6309 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3237 : btb_165_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6310 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3238 : btb_166_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6311 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3239 : btb_167_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6312 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3240 : btb_168_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6313 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3241 : btb_169_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6314 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3242 : btb_170_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6315 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3243 : btb_171_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6316 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3244 : btb_172_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6317 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3245 : btb_173_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6318 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3246 : btb_174_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6319 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3247 : btb_175_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6320 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3248 : btb_176_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6321 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3249 : btb_177_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6322 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3250 : btb_178_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6323 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3251 : btb_179_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6324 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3252 : btb_180_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6325 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3253 : btb_181_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6326 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3254 : btb_182_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6327 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3255 : btb_183_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6328 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3256 : btb_184_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6329 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3257 : btb_185_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6330 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3258 : btb_186_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6331 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3259 : btb_187_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6332 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3260 : btb_188_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6333 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3261 : btb_189_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6334 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3262 : btb_190_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6335 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3263 : btb_191_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6336 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3264 : btb_192_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6337 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3265 : btb_193_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6338 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3266 : btb_194_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6339 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3267 : btb_195_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6340 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3268 : btb_196_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6341 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3269 : btb_197_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6342 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3270 : btb_198_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6343 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3271 : btb_199_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6344 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3272 : btb_200_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6345 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3273 : btb_201_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6346 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3274 : btb_202_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6347 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3275 : btb_203_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6348 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3276 : btb_204_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6349 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3277 : btb_205_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6350 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3278 : btb_206_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6351 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3279 : btb_207_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6352 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3280 : btb_208_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6353 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3281 : btb_209_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6354 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3282 : btb_210_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6355 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3283 : btb_211_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6356 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3284 : btb_212_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6357 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3285 : btb_213_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6358 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3286 : btb_214_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6359 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3287 : btb_215_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6360 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3288 : btb_216_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6361 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3289 : btb_217_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6362 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3290 : btb_218_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6363 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3291 : btb_219_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6364 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3292 : btb_220_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6365 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3293 : btb_221_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6366 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3294 : btb_222_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6367 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3295 : btb_223_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6368 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3296 : btb_224_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6369 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3297 : btb_225_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6370 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3298 : btb_226_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6371 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3299 : btb_227_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6372 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3300 : btb_228_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6373 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3301 : btb_229_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6374 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3302 : btb_230_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6375 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3303 : btb_231_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6376 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3304 : btb_232_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6377 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3305 : btb_233_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6378 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3306 : btb_234_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6379 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3307 : btb_235_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6380 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3308 : btb_236_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6381 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3309 : btb_237_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6382 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3310 : btb_238_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6383 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3311 : btb_239_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6384 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3312 : btb_240_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6385 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3313 : btb_241_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6386 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3314 : btb_242_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6387 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3315 : btb_243_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6388 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3316 : btb_244_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6389 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3317 : btb_245_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6390 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3318 : btb_246_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6391 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3319 : btb_247_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6392 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3320 : btb_248_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6393 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3321 : btb_249_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6394 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3322 : btb_250_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6395 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3323 : btb_251_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6396 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3324 : btb_252_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6397 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3325 : btb_253_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6398 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3326 : btb_254_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6399 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3327 : btb_255_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6400 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3328 : btb_256_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6401 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3329 : btb_257_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6402 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3330 : btb_258_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6403 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3331 : btb_259_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6404 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3332 : btb_260_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6405 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3333 : btb_261_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6406 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3334 : btb_262_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6407 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3335 : btb_263_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6408 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3336 : btb_264_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6409 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3337 : btb_265_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6410 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3338 : btb_266_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6411 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3339 : btb_267_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6412 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3340 : btb_268_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6413 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3341 : btb_269_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6414 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3342 : btb_270_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6415 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3343 : btb_271_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6416 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3344 : btb_272_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6417 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3345 : btb_273_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6418 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3346 : btb_274_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6419 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3347 : btb_275_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6420 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3348 : btb_276_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6421 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3349 : btb_277_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6422 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3350 : btb_278_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6423 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3351 : btb_279_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6424 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3352 : btb_280_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6425 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3353 : btb_281_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6426 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3354 : btb_282_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6427 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3355 : btb_283_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6428 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3356 : btb_284_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6429 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3357 : btb_285_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6430 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3358 : btb_286_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6431 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3359 : btb_287_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6432 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3360 : btb_288_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6433 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3361 : btb_289_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6434 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3362 : btb_290_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6435 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3363 : btb_291_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6436 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3364 : btb_292_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6437 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3365 : btb_293_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6438 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3366 : btb_294_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6439 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3367 : btb_295_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6440 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3368 : btb_296_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6441 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3369 : btb_297_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6442 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3370 : btb_298_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6443 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3371 : btb_299_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6444 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3372 : btb_300_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6445 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3373 : btb_301_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6446 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3374 : btb_302_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6447 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3375 : btb_303_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6448 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3376 : btb_304_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6449 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3377 : btb_305_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6450 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3378 : btb_306_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6451 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3379 : btb_307_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6452 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3380 : btb_308_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6453 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3381 : btb_309_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6454 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3382 : btb_310_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6455 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3383 : btb_311_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6456 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3384 : btb_312_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6457 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3385 : btb_313_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6458 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3386 : btb_314_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6459 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3387 : btb_315_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6460 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3388 : btb_316_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6461 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3389 : btb_317_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6462 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3390 : btb_318_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6463 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3391 : btb_319_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6464 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3392 : btb_320_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6465 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3393 : btb_321_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6466 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3394 : btb_322_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6467 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3395 : btb_323_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6468 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3396 : btb_324_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6469 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3397 : btb_325_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6470 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3398 : btb_326_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6471 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3399 : btb_327_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6472 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3400 : btb_328_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6473 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3401 : btb_329_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6474 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3402 : btb_330_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6475 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3403 : btb_331_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6476 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3404 : btb_332_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6477 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3405 : btb_333_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6478 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3406 : btb_334_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6479 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3407 : btb_335_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6480 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3408 : btb_336_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6481 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3409 : btb_337_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6482 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3410 : btb_338_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6483 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3411 : btb_339_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6484 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3412 : btb_340_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6485 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3413 : btb_341_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6486 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3414 : btb_342_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6487 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3415 : btb_343_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6488 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3416 : btb_344_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6489 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3417 : btb_345_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6490 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3418 : btb_346_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6491 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3419 : btb_347_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6492 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3420 : btb_348_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6493 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3421 : btb_349_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6494 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3422 : btb_350_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6495 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3423 : btb_351_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6496 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3424 : btb_352_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6497 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3425 : btb_353_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6498 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3426 : btb_354_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6499 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3427 : btb_355_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6500 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3428 : btb_356_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6501 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3429 : btb_357_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6502 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3430 : btb_358_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6503 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3431 : btb_359_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6504 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3432 : btb_360_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6505 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3433 : btb_361_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6506 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3434 : btb_362_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6507 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3435 : btb_363_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6508 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3436 : btb_364_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6509 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3437 : btb_365_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6510 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3438 : btb_366_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6511 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3439 : btb_367_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6512 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3440 : btb_368_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6513 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3441 : btb_369_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6514 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3442 : btb_370_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6515 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3443 : btb_371_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6516 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3444 : btb_372_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6517 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3445 : btb_373_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6518 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3446 : btb_374_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6519 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3447 : btb_375_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6520 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3448 : btb_376_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6521 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3449 : btb_377_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6522 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3450 : btb_378_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6523 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3451 : btb_379_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6524 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3452 : btb_380_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6525 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3453 : btb_381_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6526 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3454 : btb_382_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6527 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3455 : btb_383_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6528 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3456 : btb_384_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6529 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3457 : btb_385_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6530 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3458 : btb_386_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6531 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3459 : btb_387_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6532 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3460 : btb_388_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6533 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3461 : btb_389_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6534 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3462 : btb_390_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6535 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3463 : btb_391_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6536 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3464 : btb_392_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6537 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3465 : btb_393_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6538 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3466 : btb_394_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6539 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3467 : btb_395_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6540 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3468 : btb_396_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6541 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3469 : btb_397_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6542 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3470 : btb_398_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6543 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3471 : btb_399_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6544 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3472 : btb_400_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6545 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3473 : btb_401_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6546 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3474 : btb_402_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6547 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3475 : btb_403_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6548 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3476 : btb_404_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6549 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3477 : btb_405_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6550 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3478 : btb_406_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6551 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3479 : btb_407_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6552 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3480 : btb_408_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6553 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3481 : btb_409_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6554 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3482 : btb_410_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6555 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3483 : btb_411_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6556 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3484 : btb_412_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6557 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3485 : btb_413_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6558 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3486 : btb_414_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6559 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3487 : btb_415_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6560 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3488 : btb_416_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6561 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3489 : btb_417_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6562 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3490 : btb_418_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6563 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3491 : btb_419_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6564 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3492 : btb_420_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6565 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3493 : btb_421_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6566 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3494 : btb_422_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6567 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3495 : btb_423_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6568 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3496 : btb_424_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6569 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3497 : btb_425_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6570 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3498 : btb_426_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6571 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3499 : btb_427_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6572 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3500 : btb_428_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6573 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3501 : btb_429_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6574 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3502 : btb_430_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6575 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3503 : btb_431_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6576 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3504 : btb_432_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6577 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3505 : btb_433_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6578 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3506 : btb_434_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6579 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3507 : btb_435_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6580 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3508 : btb_436_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6581 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3509 : btb_437_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6582 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3510 : btb_438_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6583 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3511 : btb_439_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6584 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3512 : btb_440_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6585 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3513 : btb_441_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6586 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3514 : btb_442_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6587 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3515 : btb_443_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6588 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3516 : btb_444_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6589 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3517 : btb_445_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6590 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3518 : btb_446_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6591 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3519 : btb_447_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6592 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3520 : btb_448_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6593 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3521 : btb_449_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6594 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3522 : btb_450_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6595 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3523 : btb_451_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6596 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3524 : btb_452_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6597 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3525 : btb_453_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6598 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3526 : btb_454_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6599 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3527 : btb_455_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6600 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3528 : btb_456_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6601 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3529 : btb_457_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6602 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3530 : btb_458_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6603 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3531 : btb_459_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6604 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3532 : btb_460_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6605 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3533 : btb_461_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6606 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3534 : btb_462_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6607 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3535 : btb_463_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6608 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3536 : btb_464_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6609 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3537 : btb_465_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6610 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3538 : btb_466_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6611 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3539 : btb_467_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6612 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3540 : btb_468_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6613 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3541 : btb_469_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6614 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3542 : btb_470_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6615 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3543 : btb_471_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6616 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3544 : btb_472_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6617 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3545 : btb_473_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6618 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3546 : btb_474_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6619 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3547 : btb_475_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6620 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3548 : btb_476_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6621 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3549 : btb_477_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6622 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3550 : btb_478_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6623 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3551 : btb_479_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6624 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3552 : btb_480_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6625 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3553 : btb_481_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6626 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3554 : btb_482_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6627 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3555 : btb_483_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6628 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3556 : btb_484_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6629 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3557 : btb_485_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6630 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3558 : btb_486_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6631 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3559 : btb_487_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6632 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3560 : btb_488_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6633 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3561 : btb_489_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6634 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3562 : btb_490_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6635 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3563 : btb_491_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6636 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3564 : btb_492_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6637 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3565 : btb_493_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6638 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3566 : btb_494_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6639 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3567 : btb_495_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6640 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3568 : btb_496_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6641 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3569 : btb_497_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6642 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3570 : btb_498_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6643 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3571 : btb_499_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6644 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3572 : btb_500_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6645 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3573 : btb_501_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6646 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3574 : btb_502_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6647 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3575 : btb_503_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6648 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3576 : btb_504_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6649 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3577 : btb_505_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6650 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3578 : btb_506_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6651 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3579 : btb_507_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6652 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3580 : btb_508_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6653 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3581 : btb_509_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6654 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3582 : btb_510_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [9:0] _GEN_6655 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3583 : btb_511_tag; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6656 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3584 : btb_0_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6657 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3585 : btb_1_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6658 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3586 : btb_2_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6659 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3587 : btb_3_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6660 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3588 : btb_4_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6661 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3589 : btb_5_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6662 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3590 : btb_6_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6663 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3591 : btb_7_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6664 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3592 : btb_8_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6665 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3593 : btb_9_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6666 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3594 : btb_10_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6667 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3595 : btb_11_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6668 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3596 : btb_12_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6669 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3597 : btb_13_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6670 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3598 : btb_14_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6671 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3599 : btb_15_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6672 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3600 : btb_16_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6673 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3601 : btb_17_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6674 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3602 : btb_18_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6675 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3603 : btb_19_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6676 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3604 : btb_20_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6677 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3605 : btb_21_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6678 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3606 : btb_22_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6679 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3607 : btb_23_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6680 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3608 : btb_24_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6681 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3609 : btb_25_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6682 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3610 : btb_26_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6683 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3611 : btb_27_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6684 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3612 : btb_28_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6685 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3613 : btb_29_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6686 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3614 : btb_30_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6687 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3615 : btb_31_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6688 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3616 : btb_32_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6689 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3617 : btb_33_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6690 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3618 : btb_34_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6691 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3619 : btb_35_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6692 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3620 : btb_36_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6693 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3621 : btb_37_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6694 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3622 : btb_38_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6695 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3623 : btb_39_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6696 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3624 : btb_40_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6697 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3625 : btb_41_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6698 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3626 : btb_42_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6699 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3627 : btb_43_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6700 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3628 : btb_44_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6701 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3629 : btb_45_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6702 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3630 : btb_46_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6703 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3631 : btb_47_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6704 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3632 : btb_48_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6705 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3633 : btb_49_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6706 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3634 : btb_50_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6707 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3635 : btb_51_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6708 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3636 : btb_52_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6709 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3637 : btb_53_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6710 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3638 : btb_54_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6711 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3639 : btb_55_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6712 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3640 : btb_56_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6713 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3641 : btb_57_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6714 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3642 : btb_58_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6715 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3643 : btb_59_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6716 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3644 : btb_60_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6717 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3645 : btb_61_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6718 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3646 : btb_62_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6719 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3647 : btb_63_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6720 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3648 : btb_64_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6721 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3649 : btb_65_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6722 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3650 : btb_66_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6723 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3651 : btb_67_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6724 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3652 : btb_68_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6725 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3653 : btb_69_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6726 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3654 : btb_70_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6727 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3655 : btb_71_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6728 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3656 : btb_72_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6729 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3657 : btb_73_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6730 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3658 : btb_74_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6731 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3659 : btb_75_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6732 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3660 : btb_76_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6733 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3661 : btb_77_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6734 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3662 : btb_78_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6735 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3663 : btb_79_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6736 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3664 : btb_80_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6737 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3665 : btb_81_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6738 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3666 : btb_82_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6739 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3667 : btb_83_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6740 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3668 : btb_84_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6741 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3669 : btb_85_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6742 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3670 : btb_86_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6743 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3671 : btb_87_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6744 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3672 : btb_88_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6745 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3673 : btb_89_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6746 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3674 : btb_90_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6747 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3675 : btb_91_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6748 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3676 : btb_92_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6749 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3677 : btb_93_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6750 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3678 : btb_94_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6751 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3679 : btb_95_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6752 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3680 : btb_96_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6753 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3681 : btb_97_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6754 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3682 : btb_98_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6755 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3683 : btb_99_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6756 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3684 : btb_100_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6757 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3685 : btb_101_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6758 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3686 : btb_102_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6759 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3687 : btb_103_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6760 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3688 : btb_104_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6761 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3689 : btb_105_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6762 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3690 : btb_106_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6763 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3691 : btb_107_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6764 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3692 : btb_108_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6765 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3693 : btb_109_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6766 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3694 : btb_110_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6767 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3695 : btb_111_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6768 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3696 : btb_112_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6769 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3697 : btb_113_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6770 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3698 : btb_114_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6771 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3699 : btb_115_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6772 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3700 : btb_116_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6773 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3701 : btb_117_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6774 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3702 : btb_118_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6775 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3703 : btb_119_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6776 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3704 : btb_120_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6777 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3705 : btb_121_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6778 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3706 : btb_122_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6779 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3707 : btb_123_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6780 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3708 : btb_124_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6781 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3709 : btb_125_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6782 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3710 : btb_126_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6783 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3711 : btb_127_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6784 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3712 : btb_128_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6785 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3713 : btb_129_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6786 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3714 : btb_130_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6787 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3715 : btb_131_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6788 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3716 : btb_132_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6789 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3717 : btb_133_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6790 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3718 : btb_134_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6791 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3719 : btb_135_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6792 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3720 : btb_136_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6793 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3721 : btb_137_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6794 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3722 : btb_138_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6795 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3723 : btb_139_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6796 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3724 : btb_140_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6797 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3725 : btb_141_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6798 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3726 : btb_142_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6799 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3727 : btb_143_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6800 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3728 : btb_144_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6801 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3729 : btb_145_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6802 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3730 : btb_146_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6803 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3731 : btb_147_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6804 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3732 : btb_148_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6805 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3733 : btb_149_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6806 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3734 : btb_150_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6807 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3735 : btb_151_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6808 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3736 : btb_152_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6809 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3737 : btb_153_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6810 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3738 : btb_154_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6811 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3739 : btb_155_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6812 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3740 : btb_156_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6813 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3741 : btb_157_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6814 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3742 : btb_158_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6815 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3743 : btb_159_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6816 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3744 : btb_160_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6817 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3745 : btb_161_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6818 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3746 : btb_162_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6819 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3747 : btb_163_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6820 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3748 : btb_164_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6821 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3749 : btb_165_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6822 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3750 : btb_166_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6823 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3751 : btb_167_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6824 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3752 : btb_168_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6825 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3753 : btb_169_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6826 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3754 : btb_170_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6827 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3755 : btb_171_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6828 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3756 : btb_172_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6829 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3757 : btb_173_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6830 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3758 : btb_174_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6831 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3759 : btb_175_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6832 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3760 : btb_176_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6833 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3761 : btb_177_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6834 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3762 : btb_178_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6835 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3763 : btb_179_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6836 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3764 : btb_180_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6837 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3765 : btb_181_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6838 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3766 : btb_182_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6839 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3767 : btb_183_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6840 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3768 : btb_184_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6841 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3769 : btb_185_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6842 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3770 : btb_186_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6843 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3771 : btb_187_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6844 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3772 : btb_188_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6845 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3773 : btb_189_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6846 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3774 : btb_190_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6847 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3775 : btb_191_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6848 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3776 : btb_192_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6849 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3777 : btb_193_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6850 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3778 : btb_194_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6851 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3779 : btb_195_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6852 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3780 : btb_196_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6853 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3781 : btb_197_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6854 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3782 : btb_198_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6855 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3783 : btb_199_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6856 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3784 : btb_200_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6857 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3785 : btb_201_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6858 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3786 : btb_202_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6859 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3787 : btb_203_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6860 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3788 : btb_204_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6861 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3789 : btb_205_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6862 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3790 : btb_206_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6863 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3791 : btb_207_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6864 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3792 : btb_208_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6865 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3793 : btb_209_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6866 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3794 : btb_210_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6867 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3795 : btb_211_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6868 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3796 : btb_212_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6869 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3797 : btb_213_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6870 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3798 : btb_214_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6871 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3799 : btb_215_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6872 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3800 : btb_216_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6873 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3801 : btb_217_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6874 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3802 : btb_218_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6875 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3803 : btb_219_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6876 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3804 : btb_220_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6877 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3805 : btb_221_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6878 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3806 : btb_222_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6879 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3807 : btb_223_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6880 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3808 : btb_224_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6881 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3809 : btb_225_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6882 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3810 : btb_226_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6883 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3811 : btb_227_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6884 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3812 : btb_228_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6885 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3813 : btb_229_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6886 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3814 : btb_230_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6887 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3815 : btb_231_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6888 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3816 : btb_232_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6889 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3817 : btb_233_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6890 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3818 : btb_234_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6891 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3819 : btb_235_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6892 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3820 : btb_236_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6893 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3821 : btb_237_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6894 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3822 : btb_238_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6895 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3823 : btb_239_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6896 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3824 : btb_240_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6897 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3825 : btb_241_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6898 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3826 : btb_242_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6899 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3827 : btb_243_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6900 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3828 : btb_244_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6901 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3829 : btb_245_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6902 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3830 : btb_246_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6903 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3831 : btb_247_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6904 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3832 : btb_248_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6905 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3833 : btb_249_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6906 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3834 : btb_250_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6907 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3835 : btb_251_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6908 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3836 : btb_252_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6909 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3837 : btb_253_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6910 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3838 : btb_254_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6911 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3839 : btb_255_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6912 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3840 : btb_256_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6913 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3841 : btb_257_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6914 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3842 : btb_258_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6915 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3843 : btb_259_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6916 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3844 : btb_260_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6917 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3845 : btb_261_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6918 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3846 : btb_262_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6919 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3847 : btb_263_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6920 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3848 : btb_264_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6921 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3849 : btb_265_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6922 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3850 : btb_266_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6923 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3851 : btb_267_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6924 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3852 : btb_268_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6925 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3853 : btb_269_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6926 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3854 : btb_270_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6927 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3855 : btb_271_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6928 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3856 : btb_272_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6929 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3857 : btb_273_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6930 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3858 : btb_274_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6931 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3859 : btb_275_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6932 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3860 : btb_276_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6933 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3861 : btb_277_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6934 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3862 : btb_278_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6935 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3863 : btb_279_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6936 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3864 : btb_280_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6937 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3865 : btb_281_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6938 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3866 : btb_282_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6939 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3867 : btb_283_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6940 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3868 : btb_284_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6941 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3869 : btb_285_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6942 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3870 : btb_286_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6943 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3871 : btb_287_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6944 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3872 : btb_288_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6945 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3873 : btb_289_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6946 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3874 : btb_290_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6947 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3875 : btb_291_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6948 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3876 : btb_292_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6949 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3877 : btb_293_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6950 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3878 : btb_294_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6951 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3879 : btb_295_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6952 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3880 : btb_296_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6953 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3881 : btb_297_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6954 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3882 : btb_298_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6955 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3883 : btb_299_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6956 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3884 : btb_300_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6957 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3885 : btb_301_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6958 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3886 : btb_302_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6959 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3887 : btb_303_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6960 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3888 : btb_304_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6961 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3889 : btb_305_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6962 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3890 : btb_306_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6963 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3891 : btb_307_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6964 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3892 : btb_308_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6965 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3893 : btb_309_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6966 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3894 : btb_310_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6967 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3895 : btb_311_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6968 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3896 : btb_312_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6969 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3897 : btb_313_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6970 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3898 : btb_314_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6971 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3899 : btb_315_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6972 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3900 : btb_316_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6973 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3901 : btb_317_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6974 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3902 : btb_318_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6975 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3903 : btb_319_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6976 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3904 : btb_320_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6977 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3905 : btb_321_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6978 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3906 : btb_322_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6979 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3907 : btb_323_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6980 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3908 : btb_324_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6981 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3909 : btb_325_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6982 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3910 : btb_326_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6983 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3911 : btb_327_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6984 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3912 : btb_328_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6985 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3913 : btb_329_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6986 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3914 : btb_330_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6987 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3915 : btb_331_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6988 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3916 : btb_332_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6989 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3917 : btb_333_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6990 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3918 : btb_334_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6991 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3919 : btb_335_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6992 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3920 : btb_336_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6993 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3921 : btb_337_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6994 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3922 : btb_338_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6995 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3923 : btb_339_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6996 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3924 : btb_340_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6997 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3925 : btb_341_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6998 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3926 : btb_342_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_6999 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3927 : btb_343_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7000 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3928 : btb_344_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7001 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3929 : btb_345_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7002 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3930 : btb_346_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7003 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3931 : btb_347_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7004 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3932 : btb_348_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7005 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3933 : btb_349_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7006 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3934 : btb_350_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7007 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3935 : btb_351_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7008 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3936 : btb_352_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7009 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3937 : btb_353_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7010 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3938 : btb_354_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7011 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3939 : btb_355_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7012 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3940 : btb_356_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7013 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3941 : btb_357_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7014 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3942 : btb_358_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7015 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3943 : btb_359_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7016 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3944 : btb_360_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7017 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3945 : btb_361_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7018 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3946 : btb_362_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7019 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3947 : btb_363_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7020 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3948 : btb_364_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7021 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3949 : btb_365_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7022 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3950 : btb_366_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7023 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3951 : btb_367_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7024 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3952 : btb_368_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7025 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3953 : btb_369_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7026 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3954 : btb_370_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7027 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3955 : btb_371_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7028 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3956 : btb_372_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7029 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3957 : btb_373_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7030 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3958 : btb_374_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7031 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3959 : btb_375_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7032 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3960 : btb_376_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7033 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3961 : btb_377_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7034 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3962 : btb_378_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7035 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3963 : btb_379_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7036 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3964 : btb_380_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7037 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3965 : btb_381_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7038 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3966 : btb_382_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7039 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3967 : btb_383_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7040 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3968 : btb_384_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7041 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3969 : btb_385_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7042 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3970 : btb_386_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7043 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3971 : btb_387_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7044 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3972 : btb_388_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7045 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3973 : btb_389_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7046 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3974 : btb_390_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7047 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3975 : btb_391_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7048 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3976 : btb_392_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7049 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3977 : btb_393_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7050 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3978 : btb_394_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7051 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3979 : btb_395_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7052 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3980 : btb_396_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7053 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3981 : btb_397_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7054 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3982 : btb_398_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7055 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3983 : btb_399_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7056 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3984 : btb_400_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7057 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3985 : btb_401_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7058 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3986 : btb_402_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7059 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3987 : btb_403_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7060 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3988 : btb_404_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7061 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3989 : btb_405_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7062 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3990 : btb_406_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7063 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3991 : btb_407_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7064 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3992 : btb_408_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7065 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3993 : btb_409_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7066 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3994 : btb_410_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7067 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3995 : btb_411_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7068 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3996 : btb_412_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7069 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3997 : btb_413_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7070 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3998 : btb_414_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7071 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_3999 : btb_415_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7072 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4000 : btb_416_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7073 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4001 : btb_417_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7074 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4002 : btb_418_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7075 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4003 : btb_419_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7076 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4004 : btb_420_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7077 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4005 : btb_421_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7078 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4006 : btb_422_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7079 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4007 : btb_423_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7080 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4008 : btb_424_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7081 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4009 : btb_425_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7082 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4010 : btb_426_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7083 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4011 : btb_427_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7084 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4012 : btb_428_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7085 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4013 : btb_429_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7086 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4014 : btb_430_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7087 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4015 : btb_431_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7088 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4016 : btb_432_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7089 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4017 : btb_433_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7090 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4018 : btb_434_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7091 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4019 : btb_435_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7092 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4020 : btb_436_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7093 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4021 : btb_437_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7094 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4022 : btb_438_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7095 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4023 : btb_439_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7096 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4024 : btb_440_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7097 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4025 : btb_441_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7098 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4026 : btb_442_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7099 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4027 : btb_443_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7100 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4028 : btb_444_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7101 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4029 : btb_445_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7102 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4030 : btb_446_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7103 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4031 : btb_447_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7104 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4032 : btb_448_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7105 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4033 : btb_449_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7106 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4034 : btb_450_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7107 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4035 : btb_451_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7108 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4036 : btb_452_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7109 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4037 : btb_453_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7110 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4038 : btb_454_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7111 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4039 : btb_455_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7112 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4040 : btb_456_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7113 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4041 : btb_457_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7114 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4042 : btb_458_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7115 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4043 : btb_459_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7116 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4044 : btb_460_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7117 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4045 : btb_461_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7118 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4046 : btb_462_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7119 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4047 : btb_463_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7120 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4048 : btb_464_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7121 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4049 : btb_465_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7122 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4050 : btb_466_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7123 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4051 : btb_467_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7124 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4052 : btb_468_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7125 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4053 : btb_469_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7126 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4054 : btb_470_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7127 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4055 : btb_471_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7128 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4056 : btb_472_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7129 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4057 : btb_473_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7130 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4058 : btb_474_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7131 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4059 : btb_475_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7132 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4060 : btb_476_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7133 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4061 : btb_477_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7134 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4062 : btb_478_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7135 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4063 : btb_479_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7136 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4064 : btb_480_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7137 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4065 : btb_481_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7138 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4066 : btb_482_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7139 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4067 : btb_483_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7140 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4068 : btb_484_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7141 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4069 : btb_485_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7142 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4070 : btb_486_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7143 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4071 : btb_487_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7144 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4072 : btb_488_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7145 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4073 : btb_489_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7146 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4074 : btb_490_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7147 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4075 : btb_491_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7148 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4076 : btb_492_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7149 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4077 : btb_493_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7150 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4078 : btb_494_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7151 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4079 : btb_495_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7152 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4080 : btb_496_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7153 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4081 : btb_497_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7154 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4082 : btb_498_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7155 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4083 : btb_499_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7156 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4084 : btb_500_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7157 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4085 : btb_501_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7158 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4086 : btb_502_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7159 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4087 : btb_503_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7160 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4088 : btb_504_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7161 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4089 : btb_505_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7162 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4090 : btb_506_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7163 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4091 : btb_507_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7164 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4092 : btb_508_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7165 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4093 : btb_509_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7166 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4094 : btb_510_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [63:0] _GEN_7167 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_4095 : btb_511_target_address; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8192 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5120 : btb_0_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8193 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5121 : btb_1_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8194 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5122 : btb_2_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8195 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5123 : btb_3_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8196 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5124 : btb_4_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8197 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5125 : btb_5_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8198 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5126 : btb_6_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8199 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5127 : btb_7_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8200 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5128 : btb_8_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8201 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5129 : btb_9_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8202 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5130 : btb_10_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8203 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5131 : btb_11_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8204 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5132 : btb_12_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8205 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5133 : btb_13_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8206 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5134 : btb_14_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8207 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5135 : btb_15_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8208 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5136 : btb_16_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8209 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5137 : btb_17_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8210 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5138 : btb_18_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8211 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5139 : btb_19_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8212 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5140 : btb_20_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8213 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5141 : btb_21_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8214 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5142 : btb_22_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8215 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5143 : btb_23_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8216 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5144 : btb_24_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8217 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5145 : btb_25_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8218 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5146 : btb_26_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8219 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5147 : btb_27_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8220 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5148 : btb_28_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8221 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5149 : btb_29_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8222 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5150 : btb_30_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8223 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5151 : btb_31_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8224 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5152 : btb_32_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8225 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5153 : btb_33_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8226 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5154 : btb_34_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8227 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5155 : btb_35_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8228 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5156 : btb_36_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8229 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5157 : btb_37_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8230 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5158 : btb_38_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8231 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5159 : btb_39_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8232 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5160 : btb_40_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8233 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5161 : btb_41_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8234 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5162 : btb_42_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8235 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5163 : btb_43_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8236 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5164 : btb_44_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8237 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5165 : btb_45_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8238 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5166 : btb_46_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8239 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5167 : btb_47_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8240 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5168 : btb_48_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8241 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5169 : btb_49_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8242 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5170 : btb_50_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8243 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5171 : btb_51_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8244 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5172 : btb_52_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8245 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5173 : btb_53_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8246 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5174 : btb_54_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8247 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5175 : btb_55_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8248 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5176 : btb_56_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8249 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5177 : btb_57_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8250 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5178 : btb_58_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8251 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5179 : btb_59_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8252 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5180 : btb_60_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8253 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5181 : btb_61_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8254 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5182 : btb_62_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8255 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5183 : btb_63_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8256 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5184 : btb_64_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8257 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5185 : btb_65_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8258 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5186 : btb_66_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8259 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5187 : btb_67_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8260 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5188 : btb_68_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8261 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5189 : btb_69_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8262 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5190 : btb_70_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8263 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5191 : btb_71_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8264 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5192 : btb_72_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8265 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5193 : btb_73_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8266 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5194 : btb_74_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8267 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5195 : btb_75_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8268 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5196 : btb_76_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8269 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5197 : btb_77_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8270 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5198 : btb_78_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8271 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5199 : btb_79_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8272 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5200 : btb_80_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8273 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5201 : btb_81_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8274 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5202 : btb_82_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8275 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5203 : btb_83_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8276 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5204 : btb_84_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8277 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5205 : btb_85_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8278 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5206 : btb_86_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8279 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5207 : btb_87_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8280 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5208 : btb_88_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8281 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5209 : btb_89_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8282 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5210 : btb_90_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8283 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5211 : btb_91_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8284 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5212 : btb_92_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8285 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5213 : btb_93_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8286 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5214 : btb_94_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8287 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5215 : btb_95_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8288 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5216 : btb_96_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8289 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5217 : btb_97_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8290 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5218 : btb_98_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8291 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5219 : btb_99_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8292 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5220 : btb_100_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8293 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5221 : btb_101_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8294 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5222 : btb_102_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8295 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5223 : btb_103_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8296 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5224 : btb_104_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8297 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5225 : btb_105_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8298 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5226 : btb_106_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8299 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5227 : btb_107_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8300 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5228 : btb_108_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8301 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5229 : btb_109_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8302 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5230 : btb_110_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8303 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5231 : btb_111_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8304 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5232 : btb_112_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8305 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5233 : btb_113_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8306 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5234 : btb_114_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8307 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5235 : btb_115_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8308 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5236 : btb_116_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8309 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5237 : btb_117_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8310 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5238 : btb_118_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8311 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5239 : btb_119_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8312 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5240 : btb_120_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8313 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5241 : btb_121_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8314 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5242 : btb_122_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8315 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5243 : btb_123_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8316 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5244 : btb_124_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8317 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5245 : btb_125_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8318 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5246 : btb_126_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8319 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5247 : btb_127_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8320 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5248 : btb_128_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8321 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5249 : btb_129_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8322 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5250 : btb_130_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8323 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5251 : btb_131_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8324 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5252 : btb_132_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8325 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5253 : btb_133_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8326 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5254 : btb_134_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8327 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5255 : btb_135_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8328 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5256 : btb_136_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8329 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5257 : btb_137_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8330 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5258 : btb_138_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8331 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5259 : btb_139_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8332 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5260 : btb_140_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8333 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5261 : btb_141_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8334 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5262 : btb_142_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8335 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5263 : btb_143_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8336 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5264 : btb_144_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8337 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5265 : btb_145_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8338 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5266 : btb_146_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8339 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5267 : btb_147_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8340 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5268 : btb_148_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8341 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5269 : btb_149_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8342 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5270 : btb_150_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8343 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5271 : btb_151_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8344 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5272 : btb_152_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8345 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5273 : btb_153_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8346 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5274 : btb_154_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8347 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5275 : btb_155_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8348 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5276 : btb_156_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8349 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5277 : btb_157_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8350 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5278 : btb_158_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8351 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5279 : btb_159_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8352 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5280 : btb_160_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8353 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5281 : btb_161_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8354 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5282 : btb_162_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8355 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5283 : btb_163_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8356 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5284 : btb_164_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8357 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5285 : btb_165_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8358 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5286 : btb_166_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8359 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5287 : btb_167_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8360 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5288 : btb_168_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8361 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5289 : btb_169_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8362 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5290 : btb_170_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8363 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5291 : btb_171_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8364 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5292 : btb_172_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8365 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5293 : btb_173_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8366 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5294 : btb_174_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8367 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5295 : btb_175_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8368 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5296 : btb_176_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8369 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5297 : btb_177_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8370 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5298 : btb_178_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8371 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5299 : btb_179_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8372 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5300 : btb_180_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8373 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5301 : btb_181_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8374 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5302 : btb_182_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8375 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5303 : btb_183_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8376 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5304 : btb_184_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8377 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5305 : btb_185_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8378 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5306 : btb_186_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8379 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5307 : btb_187_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8380 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5308 : btb_188_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8381 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5309 : btb_189_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8382 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5310 : btb_190_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8383 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5311 : btb_191_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8384 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5312 : btb_192_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8385 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5313 : btb_193_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8386 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5314 : btb_194_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8387 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5315 : btb_195_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8388 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5316 : btb_196_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8389 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5317 : btb_197_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8390 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5318 : btb_198_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8391 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5319 : btb_199_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8392 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5320 : btb_200_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8393 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5321 : btb_201_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8394 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5322 : btb_202_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8395 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5323 : btb_203_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8396 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5324 : btb_204_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8397 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5325 : btb_205_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8398 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5326 : btb_206_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8399 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5327 : btb_207_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8400 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5328 : btb_208_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8401 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5329 : btb_209_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8402 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5330 : btb_210_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8403 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5331 : btb_211_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8404 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5332 : btb_212_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8405 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5333 : btb_213_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8406 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5334 : btb_214_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8407 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5335 : btb_215_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8408 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5336 : btb_216_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8409 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5337 : btb_217_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8410 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5338 : btb_218_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8411 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5339 : btb_219_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8412 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5340 : btb_220_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8413 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5341 : btb_221_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8414 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5342 : btb_222_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8415 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5343 : btb_223_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8416 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5344 : btb_224_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8417 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5345 : btb_225_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8418 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5346 : btb_226_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8419 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5347 : btb_227_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8420 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5348 : btb_228_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8421 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5349 : btb_229_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8422 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5350 : btb_230_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8423 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5351 : btb_231_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8424 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5352 : btb_232_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8425 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5353 : btb_233_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8426 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5354 : btb_234_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8427 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5355 : btb_235_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8428 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5356 : btb_236_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8429 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5357 : btb_237_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8430 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5358 : btb_238_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8431 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5359 : btb_239_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8432 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5360 : btb_240_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8433 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5361 : btb_241_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8434 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5362 : btb_242_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8435 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5363 : btb_243_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8436 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5364 : btb_244_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8437 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5365 : btb_245_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8438 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5366 : btb_246_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8439 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5367 : btb_247_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8440 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5368 : btb_248_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8441 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5369 : btb_249_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8442 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5370 : btb_250_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8443 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5371 : btb_251_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8444 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5372 : btb_252_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8445 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5373 : btb_253_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8446 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5374 : btb_254_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8447 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5375 : btb_255_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8448 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5376 : btb_256_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8449 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5377 : btb_257_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8450 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5378 : btb_258_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8451 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5379 : btb_259_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8452 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5380 : btb_260_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8453 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5381 : btb_261_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8454 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5382 : btb_262_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8455 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5383 : btb_263_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8456 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5384 : btb_264_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8457 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5385 : btb_265_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8458 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5386 : btb_266_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8459 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5387 : btb_267_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8460 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5388 : btb_268_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8461 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5389 : btb_269_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8462 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5390 : btb_270_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8463 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5391 : btb_271_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8464 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5392 : btb_272_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8465 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5393 : btb_273_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8466 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5394 : btb_274_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8467 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5395 : btb_275_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8468 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5396 : btb_276_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8469 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5397 : btb_277_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8470 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5398 : btb_278_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8471 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5399 : btb_279_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8472 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5400 : btb_280_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8473 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5401 : btb_281_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8474 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5402 : btb_282_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8475 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5403 : btb_283_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8476 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5404 : btb_284_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8477 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5405 : btb_285_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8478 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5406 : btb_286_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8479 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5407 : btb_287_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8480 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5408 : btb_288_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8481 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5409 : btb_289_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8482 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5410 : btb_290_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8483 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5411 : btb_291_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8484 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5412 : btb_292_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8485 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5413 : btb_293_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8486 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5414 : btb_294_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8487 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5415 : btb_295_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8488 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5416 : btb_296_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8489 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5417 : btb_297_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8490 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5418 : btb_298_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8491 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5419 : btb_299_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8492 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5420 : btb_300_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8493 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5421 : btb_301_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8494 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5422 : btb_302_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8495 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5423 : btb_303_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8496 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5424 : btb_304_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8497 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5425 : btb_305_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8498 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5426 : btb_306_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8499 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5427 : btb_307_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8500 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5428 : btb_308_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8501 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5429 : btb_309_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8502 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5430 : btb_310_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8503 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5431 : btb_311_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8504 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5432 : btb_312_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8505 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5433 : btb_313_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8506 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5434 : btb_314_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8507 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5435 : btb_315_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8508 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5436 : btb_316_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8509 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5437 : btb_317_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8510 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5438 : btb_318_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8511 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5439 : btb_319_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8512 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5440 : btb_320_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8513 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5441 : btb_321_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8514 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5442 : btb_322_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8515 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5443 : btb_323_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8516 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5444 : btb_324_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8517 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5445 : btb_325_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8518 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5446 : btb_326_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8519 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5447 : btb_327_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8520 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5448 : btb_328_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8521 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5449 : btb_329_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8522 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5450 : btb_330_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8523 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5451 : btb_331_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8524 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5452 : btb_332_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8525 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5453 : btb_333_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8526 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5454 : btb_334_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8527 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5455 : btb_335_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8528 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5456 : btb_336_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8529 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5457 : btb_337_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8530 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5458 : btb_338_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8531 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5459 : btb_339_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8532 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5460 : btb_340_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8533 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5461 : btb_341_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8534 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5462 : btb_342_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8535 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5463 : btb_343_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8536 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5464 : btb_344_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8537 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5465 : btb_345_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8538 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5466 : btb_346_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8539 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5467 : btb_347_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8540 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5468 : btb_348_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8541 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5469 : btb_349_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8542 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5470 : btb_350_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8543 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5471 : btb_351_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8544 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5472 : btb_352_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8545 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5473 : btb_353_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8546 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5474 : btb_354_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8547 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5475 : btb_355_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8548 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5476 : btb_356_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8549 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5477 : btb_357_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8550 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5478 : btb_358_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8551 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5479 : btb_359_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8552 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5480 : btb_360_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8553 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5481 : btb_361_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8554 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5482 : btb_362_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8555 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5483 : btb_363_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8556 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5484 : btb_364_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8557 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5485 : btb_365_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8558 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5486 : btb_366_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8559 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5487 : btb_367_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8560 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5488 : btb_368_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8561 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5489 : btb_369_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8562 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5490 : btb_370_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8563 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5491 : btb_371_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8564 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5492 : btb_372_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8565 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5493 : btb_373_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8566 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5494 : btb_374_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8567 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5495 : btb_375_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8568 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5496 : btb_376_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8569 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5497 : btb_377_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8570 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5498 : btb_378_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8571 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5499 : btb_379_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8572 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5500 : btb_380_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8573 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5501 : btb_381_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8574 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5502 : btb_382_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8575 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5503 : btb_383_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8576 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5504 : btb_384_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8577 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5505 : btb_385_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8578 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5506 : btb_386_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8579 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5507 : btb_387_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8580 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5508 : btb_388_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8581 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5509 : btb_389_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8582 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5510 : btb_390_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8583 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5511 : btb_391_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8584 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5512 : btb_392_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8585 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5513 : btb_393_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8586 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5514 : btb_394_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8587 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5515 : btb_395_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8588 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5516 : btb_396_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8589 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5517 : btb_397_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8590 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5518 : btb_398_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8591 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5519 : btb_399_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8592 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5520 : btb_400_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8593 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5521 : btb_401_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8594 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5522 : btb_402_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8595 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5523 : btb_403_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8596 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5524 : btb_404_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8597 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5525 : btb_405_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8598 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5526 : btb_406_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8599 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5527 : btb_407_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8600 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5528 : btb_408_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8601 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5529 : btb_409_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8602 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5530 : btb_410_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8603 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5531 : btb_411_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8604 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5532 : btb_412_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8605 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5533 : btb_413_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8606 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5534 : btb_414_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8607 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5535 : btb_415_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8608 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5536 : btb_416_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8609 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5537 : btb_417_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8610 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5538 : btb_418_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8611 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5539 : btb_419_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8612 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5540 : btb_420_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8613 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5541 : btb_421_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8614 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5542 : btb_422_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8615 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5543 : btb_423_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8616 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5544 : btb_424_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8617 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5545 : btb_425_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8618 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5546 : btb_426_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8619 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5547 : btb_427_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8620 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5548 : btb_428_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8621 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5549 : btb_429_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8622 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5550 : btb_430_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8623 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5551 : btb_431_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8624 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5552 : btb_432_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8625 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5553 : btb_433_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8626 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5554 : btb_434_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8627 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5555 : btb_435_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8628 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5556 : btb_436_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8629 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5557 : btb_437_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8630 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5558 : btb_438_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8631 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5559 : btb_439_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8632 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5560 : btb_440_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8633 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5561 : btb_441_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8634 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5562 : btb_442_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8635 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5563 : btb_443_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8636 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5564 : btb_444_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8637 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5565 : btb_445_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8638 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5566 : btb_446_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8639 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5567 : btb_447_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8640 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5568 : btb_448_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8641 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5569 : btb_449_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8642 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5570 : btb_450_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8643 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5571 : btb_451_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8644 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5572 : btb_452_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8645 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5573 : btb_453_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8646 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5574 : btb_454_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8647 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5575 : btb_455_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8648 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5576 : btb_456_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8649 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5577 : btb_457_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8650 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5578 : btb_458_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8651 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5579 : btb_459_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8652 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5580 : btb_460_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8653 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5581 : btb_461_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8654 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5582 : btb_462_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8655 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5583 : btb_463_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8656 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5584 : btb_464_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8657 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5585 : btb_465_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8658 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5586 : btb_466_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8659 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5587 : btb_467_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8660 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5588 : btb_468_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8661 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5589 : btb_469_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8662 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5590 : btb_470_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8663 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5591 : btb_471_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8664 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5592 : btb_472_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8665 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5593 : btb_473_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8666 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5594 : btb_474_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8667 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5595 : btb_475_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8668 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5596 : btb_476_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8669 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5597 : btb_477_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8670 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5598 : btb_478_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8671 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5599 : btb_479_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8672 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5600 : btb_480_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8673 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5601 : btb_481_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8674 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5602 : btb_482_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8675 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5603 : btb_483_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8676 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5604 : btb_484_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8677 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5605 : btb_485_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8678 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5606 : btb_486_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8679 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5607 : btb_487_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8680 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5608 : btb_488_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8681 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5609 : btb_489_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8682 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5610 : btb_490_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8683 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5611 : btb_491_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8684 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5612 : btb_492_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8685 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5613 : btb_493_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8686 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5614 : btb_494_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8687 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5615 : btb_495_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8688 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5616 : btb_496_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8689 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5617 : btb_497_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8690 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5618 : btb_498_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8691 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5619 : btb_499_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8692 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5620 : btb_500_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8693 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5621 : btb_501_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8694 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5622 : btb_502_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8695 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5623 : btb_503_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8696 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5624 : btb_504_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8697 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5625 : btb_505_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8698 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5626 : btb_506_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8699 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5627 : btb_507_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8700 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5628 : btb_508_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8701 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5629 : btb_509_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8702 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5630 : btb_510_bht; // @[branch_predictor.scala 62:121 30:22]
  wire [1:0] _GEN_8703 = io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
    io_i_branch_resolve_pack_taken ? _GEN_5631 : btb_511_bht; // @[branch_predictor.scala 62:121 30:22]
  wire  _T_1027 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid; // @[branch_predictor.scala 77:42]
  wire  _btb_0_bht_T = btb_0_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_0_bht_T_1 = io_i_branch_resolve_pack_taken & btb_0_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_0_bht_T_2 = btb_0_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_0_bht_T_3 = io_i_branch_resolve_pack_taken & btb_0_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_0_bht_T_4 = btb_0_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_0_bht_T_5 = io_i_branch_resolve_pack_taken & btb_0_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_0_bht_T_6 = btb_0_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_0_bht_T_7 = io_i_branch_resolve_pack_taken & btb_0_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_0_bht_T_8 = ~io_i_branch_resolve_pack_taken; // @[branch_predictor.scala 89:22]
  wire  _btb_0_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_0_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_0_bht_T_13 = _btb_0_bht_T_8 & _btb_0_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_0_bht_T_16 = _btb_0_bht_T_8 & _btb_0_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_0_bht_T_19 = _btb_0_bht_T_8 & _btb_0_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_0_bht_T_20 = _btb_0_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_21 = _btb_0_bht_T_16 ? 2'h0 : _btb_0_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_22 = _btb_0_bht_T_13 ? 2'h0 : _btb_0_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_23 = _btb_0_bht_T_10 ? 2'h0 : _btb_0_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_24 = _btb_0_bht_T_7 ? 2'h3 : _btb_0_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_25 = _btb_0_bht_T_5 ? 2'h3 : _btb_0_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_26 = _btb_0_bht_T_3 ? 2'h3 : _btb_0_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_0_bht_T_27 = _btb_0_bht_T_1 ? 2'h1 : _btb_0_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8706 = btb_0_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6656; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8708 = btb_0_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_0_bht_T_27 : _GEN_8192; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_1_bht_T = btb_1_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_1_bht_T_1 = io_i_branch_resolve_pack_taken & btb_1_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_1_bht_T_2 = btb_1_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_1_bht_T_3 = io_i_branch_resolve_pack_taken & btb_1_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_1_bht_T_4 = btb_1_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_1_bht_T_5 = io_i_branch_resolve_pack_taken & btb_1_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_1_bht_T_6 = btb_1_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_1_bht_T_7 = io_i_branch_resolve_pack_taken & btb_1_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_1_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_1_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_1_bht_T_13 = _btb_0_bht_T_8 & _btb_1_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_1_bht_T_16 = _btb_0_bht_T_8 & _btb_1_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_1_bht_T_19 = _btb_0_bht_T_8 & _btb_1_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_1_bht_T_20 = _btb_1_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_21 = _btb_1_bht_T_16 ? 2'h0 : _btb_1_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_22 = _btb_1_bht_T_13 ? 2'h0 : _btb_1_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_23 = _btb_1_bht_T_10 ? 2'h0 : _btb_1_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_24 = _btb_1_bht_T_7 ? 2'h3 : _btb_1_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_25 = _btb_1_bht_T_5 ? 2'h3 : _btb_1_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_26 = _btb_1_bht_T_3 ? 2'h3 : _btb_1_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_1_bht_T_27 = _btb_1_bht_T_1 ? 2'h1 : _btb_1_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8710 = btb_1_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6657; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8712 = btb_1_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_1_bht_T_27 : _GEN_8193; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_2_bht_T = btb_2_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_2_bht_T_1 = io_i_branch_resolve_pack_taken & btb_2_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_2_bht_T_2 = btb_2_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_2_bht_T_3 = io_i_branch_resolve_pack_taken & btb_2_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_2_bht_T_4 = btb_2_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_2_bht_T_5 = io_i_branch_resolve_pack_taken & btb_2_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_2_bht_T_6 = btb_2_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_2_bht_T_7 = io_i_branch_resolve_pack_taken & btb_2_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_2_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_2_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_2_bht_T_13 = _btb_0_bht_T_8 & _btb_2_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_2_bht_T_16 = _btb_0_bht_T_8 & _btb_2_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_2_bht_T_19 = _btb_0_bht_T_8 & _btb_2_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_2_bht_T_20 = _btb_2_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_21 = _btb_2_bht_T_16 ? 2'h0 : _btb_2_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_22 = _btb_2_bht_T_13 ? 2'h0 : _btb_2_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_23 = _btb_2_bht_T_10 ? 2'h0 : _btb_2_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_24 = _btb_2_bht_T_7 ? 2'h3 : _btb_2_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_25 = _btb_2_bht_T_5 ? 2'h3 : _btb_2_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_26 = _btb_2_bht_T_3 ? 2'h3 : _btb_2_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_2_bht_T_27 = _btb_2_bht_T_1 ? 2'h1 : _btb_2_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8714 = btb_2_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6658; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8716 = btb_2_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_2_bht_T_27 : _GEN_8194; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_3_bht_T = btb_3_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_3_bht_T_1 = io_i_branch_resolve_pack_taken & btb_3_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_3_bht_T_2 = btb_3_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_3_bht_T_3 = io_i_branch_resolve_pack_taken & btb_3_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_3_bht_T_4 = btb_3_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_3_bht_T_5 = io_i_branch_resolve_pack_taken & btb_3_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_3_bht_T_6 = btb_3_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_3_bht_T_7 = io_i_branch_resolve_pack_taken & btb_3_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_3_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_3_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_3_bht_T_13 = _btb_0_bht_T_8 & _btb_3_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_3_bht_T_16 = _btb_0_bht_T_8 & _btb_3_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_3_bht_T_19 = _btb_0_bht_T_8 & _btb_3_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_3_bht_T_20 = _btb_3_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_21 = _btb_3_bht_T_16 ? 2'h0 : _btb_3_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_22 = _btb_3_bht_T_13 ? 2'h0 : _btb_3_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_23 = _btb_3_bht_T_10 ? 2'h0 : _btb_3_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_24 = _btb_3_bht_T_7 ? 2'h3 : _btb_3_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_25 = _btb_3_bht_T_5 ? 2'h3 : _btb_3_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_26 = _btb_3_bht_T_3 ? 2'h3 : _btb_3_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_3_bht_T_27 = _btb_3_bht_T_1 ? 2'h1 : _btb_3_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8718 = btb_3_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6659; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8720 = btb_3_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_3_bht_T_27 : _GEN_8195; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_4_bht_T = btb_4_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_4_bht_T_1 = io_i_branch_resolve_pack_taken & btb_4_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_4_bht_T_2 = btb_4_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_4_bht_T_3 = io_i_branch_resolve_pack_taken & btb_4_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_4_bht_T_4 = btb_4_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_4_bht_T_5 = io_i_branch_resolve_pack_taken & btb_4_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_4_bht_T_6 = btb_4_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_4_bht_T_7 = io_i_branch_resolve_pack_taken & btb_4_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_4_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_4_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_4_bht_T_13 = _btb_0_bht_T_8 & _btb_4_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_4_bht_T_16 = _btb_0_bht_T_8 & _btb_4_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_4_bht_T_19 = _btb_0_bht_T_8 & _btb_4_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_4_bht_T_20 = _btb_4_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_21 = _btb_4_bht_T_16 ? 2'h0 : _btb_4_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_22 = _btb_4_bht_T_13 ? 2'h0 : _btb_4_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_23 = _btb_4_bht_T_10 ? 2'h0 : _btb_4_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_24 = _btb_4_bht_T_7 ? 2'h3 : _btb_4_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_25 = _btb_4_bht_T_5 ? 2'h3 : _btb_4_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_26 = _btb_4_bht_T_3 ? 2'h3 : _btb_4_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_4_bht_T_27 = _btb_4_bht_T_1 ? 2'h1 : _btb_4_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8722 = btb_4_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6660; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8724 = btb_4_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_4_bht_T_27 : _GEN_8196; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_5_bht_T = btb_5_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_5_bht_T_1 = io_i_branch_resolve_pack_taken & btb_5_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_5_bht_T_2 = btb_5_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_5_bht_T_3 = io_i_branch_resolve_pack_taken & btb_5_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_5_bht_T_4 = btb_5_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_5_bht_T_5 = io_i_branch_resolve_pack_taken & btb_5_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_5_bht_T_6 = btb_5_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_5_bht_T_7 = io_i_branch_resolve_pack_taken & btb_5_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_5_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_5_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_5_bht_T_13 = _btb_0_bht_T_8 & _btb_5_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_5_bht_T_16 = _btb_0_bht_T_8 & _btb_5_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_5_bht_T_19 = _btb_0_bht_T_8 & _btb_5_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_5_bht_T_20 = _btb_5_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_21 = _btb_5_bht_T_16 ? 2'h0 : _btb_5_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_22 = _btb_5_bht_T_13 ? 2'h0 : _btb_5_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_23 = _btb_5_bht_T_10 ? 2'h0 : _btb_5_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_24 = _btb_5_bht_T_7 ? 2'h3 : _btb_5_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_25 = _btb_5_bht_T_5 ? 2'h3 : _btb_5_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_26 = _btb_5_bht_T_3 ? 2'h3 : _btb_5_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_5_bht_T_27 = _btb_5_bht_T_1 ? 2'h1 : _btb_5_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8726 = btb_5_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6661; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8728 = btb_5_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_5_bht_T_27 : _GEN_8197; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_6_bht_T = btb_6_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_6_bht_T_1 = io_i_branch_resolve_pack_taken & btb_6_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_6_bht_T_2 = btb_6_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_6_bht_T_3 = io_i_branch_resolve_pack_taken & btb_6_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_6_bht_T_4 = btb_6_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_6_bht_T_5 = io_i_branch_resolve_pack_taken & btb_6_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_6_bht_T_6 = btb_6_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_6_bht_T_7 = io_i_branch_resolve_pack_taken & btb_6_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_6_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_6_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_6_bht_T_13 = _btb_0_bht_T_8 & _btb_6_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_6_bht_T_16 = _btb_0_bht_T_8 & _btb_6_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_6_bht_T_19 = _btb_0_bht_T_8 & _btb_6_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_6_bht_T_20 = _btb_6_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_21 = _btb_6_bht_T_16 ? 2'h0 : _btb_6_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_22 = _btb_6_bht_T_13 ? 2'h0 : _btb_6_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_23 = _btb_6_bht_T_10 ? 2'h0 : _btb_6_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_24 = _btb_6_bht_T_7 ? 2'h3 : _btb_6_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_25 = _btb_6_bht_T_5 ? 2'h3 : _btb_6_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_26 = _btb_6_bht_T_3 ? 2'h3 : _btb_6_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_6_bht_T_27 = _btb_6_bht_T_1 ? 2'h1 : _btb_6_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8730 = btb_6_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6662; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8732 = btb_6_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_6_bht_T_27 : _GEN_8198; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_7_bht_T = btb_7_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_7_bht_T_1 = io_i_branch_resolve_pack_taken & btb_7_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_7_bht_T_2 = btb_7_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_7_bht_T_3 = io_i_branch_resolve_pack_taken & btb_7_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_7_bht_T_4 = btb_7_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_7_bht_T_5 = io_i_branch_resolve_pack_taken & btb_7_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_7_bht_T_6 = btb_7_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_7_bht_T_7 = io_i_branch_resolve_pack_taken & btb_7_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_7_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_7_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_7_bht_T_13 = _btb_0_bht_T_8 & _btb_7_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_7_bht_T_16 = _btb_0_bht_T_8 & _btb_7_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_7_bht_T_19 = _btb_0_bht_T_8 & _btb_7_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_7_bht_T_20 = _btb_7_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_21 = _btb_7_bht_T_16 ? 2'h0 : _btb_7_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_22 = _btb_7_bht_T_13 ? 2'h0 : _btb_7_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_23 = _btb_7_bht_T_10 ? 2'h0 : _btb_7_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_24 = _btb_7_bht_T_7 ? 2'h3 : _btb_7_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_25 = _btb_7_bht_T_5 ? 2'h3 : _btb_7_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_26 = _btb_7_bht_T_3 ? 2'h3 : _btb_7_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_7_bht_T_27 = _btb_7_bht_T_1 ? 2'h1 : _btb_7_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8734 = btb_7_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6663; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8736 = btb_7_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_7_bht_T_27 : _GEN_8199; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_8_bht_T = btb_8_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_8_bht_T_1 = io_i_branch_resolve_pack_taken & btb_8_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_8_bht_T_2 = btb_8_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_8_bht_T_3 = io_i_branch_resolve_pack_taken & btb_8_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_8_bht_T_4 = btb_8_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_8_bht_T_5 = io_i_branch_resolve_pack_taken & btb_8_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_8_bht_T_6 = btb_8_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_8_bht_T_7 = io_i_branch_resolve_pack_taken & btb_8_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_8_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_8_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_8_bht_T_13 = _btb_0_bht_T_8 & _btb_8_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_8_bht_T_16 = _btb_0_bht_T_8 & _btb_8_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_8_bht_T_19 = _btb_0_bht_T_8 & _btb_8_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_8_bht_T_20 = _btb_8_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_21 = _btb_8_bht_T_16 ? 2'h0 : _btb_8_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_22 = _btb_8_bht_T_13 ? 2'h0 : _btb_8_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_23 = _btb_8_bht_T_10 ? 2'h0 : _btb_8_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_24 = _btb_8_bht_T_7 ? 2'h3 : _btb_8_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_25 = _btb_8_bht_T_5 ? 2'h3 : _btb_8_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_26 = _btb_8_bht_T_3 ? 2'h3 : _btb_8_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_8_bht_T_27 = _btb_8_bht_T_1 ? 2'h1 : _btb_8_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8738 = btb_8_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6664; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8740 = btb_8_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_8_bht_T_27 : _GEN_8200; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_9_bht_T = btb_9_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_9_bht_T_1 = io_i_branch_resolve_pack_taken & btb_9_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_9_bht_T_2 = btb_9_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_9_bht_T_3 = io_i_branch_resolve_pack_taken & btb_9_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_9_bht_T_4 = btb_9_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_9_bht_T_5 = io_i_branch_resolve_pack_taken & btb_9_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_9_bht_T_6 = btb_9_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_9_bht_T_7 = io_i_branch_resolve_pack_taken & btb_9_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_9_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_9_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_9_bht_T_13 = _btb_0_bht_T_8 & _btb_9_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_9_bht_T_16 = _btb_0_bht_T_8 & _btb_9_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_9_bht_T_19 = _btb_0_bht_T_8 & _btb_9_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_9_bht_T_20 = _btb_9_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_21 = _btb_9_bht_T_16 ? 2'h0 : _btb_9_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_22 = _btb_9_bht_T_13 ? 2'h0 : _btb_9_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_23 = _btb_9_bht_T_10 ? 2'h0 : _btb_9_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_24 = _btb_9_bht_T_7 ? 2'h3 : _btb_9_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_25 = _btb_9_bht_T_5 ? 2'h3 : _btb_9_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_26 = _btb_9_bht_T_3 ? 2'h3 : _btb_9_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_9_bht_T_27 = _btb_9_bht_T_1 ? 2'h1 : _btb_9_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8742 = btb_9_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6665; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8744 = btb_9_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_9_bht_T_27 : _GEN_8201; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_10_bht_T = btb_10_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_10_bht_T_1 = io_i_branch_resolve_pack_taken & btb_10_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_10_bht_T_2 = btb_10_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_10_bht_T_3 = io_i_branch_resolve_pack_taken & btb_10_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_10_bht_T_4 = btb_10_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_10_bht_T_5 = io_i_branch_resolve_pack_taken & btb_10_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_10_bht_T_6 = btb_10_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_10_bht_T_7 = io_i_branch_resolve_pack_taken & btb_10_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_10_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_10_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_10_bht_T_13 = _btb_0_bht_T_8 & _btb_10_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_10_bht_T_16 = _btb_0_bht_T_8 & _btb_10_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_10_bht_T_19 = _btb_0_bht_T_8 & _btb_10_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_10_bht_T_20 = _btb_10_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_21 = _btb_10_bht_T_16 ? 2'h0 : _btb_10_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_22 = _btb_10_bht_T_13 ? 2'h0 : _btb_10_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_23 = _btb_10_bht_T_10 ? 2'h0 : _btb_10_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_24 = _btb_10_bht_T_7 ? 2'h3 : _btb_10_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_25 = _btb_10_bht_T_5 ? 2'h3 : _btb_10_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_26 = _btb_10_bht_T_3 ? 2'h3 : _btb_10_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_10_bht_T_27 = _btb_10_bht_T_1 ? 2'h1 : _btb_10_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8746 = btb_10_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6666; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8748 = btb_10_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_10_bht_T_27 : _GEN_8202; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_11_bht_T = btb_11_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_11_bht_T_1 = io_i_branch_resolve_pack_taken & btb_11_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_11_bht_T_2 = btb_11_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_11_bht_T_3 = io_i_branch_resolve_pack_taken & btb_11_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_11_bht_T_4 = btb_11_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_11_bht_T_5 = io_i_branch_resolve_pack_taken & btb_11_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_11_bht_T_6 = btb_11_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_11_bht_T_7 = io_i_branch_resolve_pack_taken & btb_11_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_11_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_11_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_11_bht_T_13 = _btb_0_bht_T_8 & _btb_11_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_11_bht_T_16 = _btb_0_bht_T_8 & _btb_11_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_11_bht_T_19 = _btb_0_bht_T_8 & _btb_11_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_11_bht_T_20 = _btb_11_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_21 = _btb_11_bht_T_16 ? 2'h0 : _btb_11_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_22 = _btb_11_bht_T_13 ? 2'h0 : _btb_11_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_23 = _btb_11_bht_T_10 ? 2'h0 : _btb_11_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_24 = _btb_11_bht_T_7 ? 2'h3 : _btb_11_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_25 = _btb_11_bht_T_5 ? 2'h3 : _btb_11_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_26 = _btb_11_bht_T_3 ? 2'h3 : _btb_11_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_11_bht_T_27 = _btb_11_bht_T_1 ? 2'h1 : _btb_11_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8750 = btb_11_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6667; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8752 = btb_11_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_11_bht_T_27 : _GEN_8203; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_12_bht_T = btb_12_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_12_bht_T_1 = io_i_branch_resolve_pack_taken & btb_12_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_12_bht_T_2 = btb_12_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_12_bht_T_3 = io_i_branch_resolve_pack_taken & btb_12_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_12_bht_T_4 = btb_12_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_12_bht_T_5 = io_i_branch_resolve_pack_taken & btb_12_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_12_bht_T_6 = btb_12_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_12_bht_T_7 = io_i_branch_resolve_pack_taken & btb_12_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_12_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_12_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_12_bht_T_13 = _btb_0_bht_T_8 & _btb_12_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_12_bht_T_16 = _btb_0_bht_T_8 & _btb_12_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_12_bht_T_19 = _btb_0_bht_T_8 & _btb_12_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_12_bht_T_20 = _btb_12_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_21 = _btb_12_bht_T_16 ? 2'h0 : _btb_12_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_22 = _btb_12_bht_T_13 ? 2'h0 : _btb_12_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_23 = _btb_12_bht_T_10 ? 2'h0 : _btb_12_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_24 = _btb_12_bht_T_7 ? 2'h3 : _btb_12_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_25 = _btb_12_bht_T_5 ? 2'h3 : _btb_12_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_26 = _btb_12_bht_T_3 ? 2'h3 : _btb_12_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_12_bht_T_27 = _btb_12_bht_T_1 ? 2'h1 : _btb_12_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8754 = btb_12_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6668; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8756 = btb_12_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_12_bht_T_27 : _GEN_8204; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_13_bht_T = btb_13_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_13_bht_T_1 = io_i_branch_resolve_pack_taken & btb_13_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_13_bht_T_2 = btb_13_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_13_bht_T_3 = io_i_branch_resolve_pack_taken & btb_13_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_13_bht_T_4 = btb_13_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_13_bht_T_5 = io_i_branch_resolve_pack_taken & btb_13_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_13_bht_T_6 = btb_13_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_13_bht_T_7 = io_i_branch_resolve_pack_taken & btb_13_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_13_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_13_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_13_bht_T_13 = _btb_0_bht_T_8 & _btb_13_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_13_bht_T_16 = _btb_0_bht_T_8 & _btb_13_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_13_bht_T_19 = _btb_0_bht_T_8 & _btb_13_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_13_bht_T_20 = _btb_13_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_21 = _btb_13_bht_T_16 ? 2'h0 : _btb_13_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_22 = _btb_13_bht_T_13 ? 2'h0 : _btb_13_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_23 = _btb_13_bht_T_10 ? 2'h0 : _btb_13_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_24 = _btb_13_bht_T_7 ? 2'h3 : _btb_13_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_25 = _btb_13_bht_T_5 ? 2'h3 : _btb_13_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_26 = _btb_13_bht_T_3 ? 2'h3 : _btb_13_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_13_bht_T_27 = _btb_13_bht_T_1 ? 2'h1 : _btb_13_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8758 = btb_13_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6669; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8760 = btb_13_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_13_bht_T_27 : _GEN_8205; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_14_bht_T = btb_14_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_14_bht_T_1 = io_i_branch_resolve_pack_taken & btb_14_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_14_bht_T_2 = btb_14_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_14_bht_T_3 = io_i_branch_resolve_pack_taken & btb_14_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_14_bht_T_4 = btb_14_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_14_bht_T_5 = io_i_branch_resolve_pack_taken & btb_14_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_14_bht_T_6 = btb_14_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_14_bht_T_7 = io_i_branch_resolve_pack_taken & btb_14_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_14_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_14_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_14_bht_T_13 = _btb_0_bht_T_8 & _btb_14_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_14_bht_T_16 = _btb_0_bht_T_8 & _btb_14_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_14_bht_T_19 = _btb_0_bht_T_8 & _btb_14_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_14_bht_T_20 = _btb_14_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_21 = _btb_14_bht_T_16 ? 2'h0 : _btb_14_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_22 = _btb_14_bht_T_13 ? 2'h0 : _btb_14_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_23 = _btb_14_bht_T_10 ? 2'h0 : _btb_14_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_24 = _btb_14_bht_T_7 ? 2'h3 : _btb_14_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_25 = _btb_14_bht_T_5 ? 2'h3 : _btb_14_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_26 = _btb_14_bht_T_3 ? 2'h3 : _btb_14_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_14_bht_T_27 = _btb_14_bht_T_1 ? 2'h1 : _btb_14_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_8761 = btb_14_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_13_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_12_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_11_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_10_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_9_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_8_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_7_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_6_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_5_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_4_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_3_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_2_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_1_tag == io_i_branch_resolve_pack_pc[12:3] | btb_0_tag ==
    io_i_branch_resolve_pack_pc[12:3]))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_8762 = btb_14_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6670; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8764 = btb_14_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_14_bht_T_27 : _GEN_8206; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_15_bht_T = btb_15_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_15_bht_T_1 = io_i_branch_resolve_pack_taken & btb_15_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_15_bht_T_2 = btb_15_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_15_bht_T_3 = io_i_branch_resolve_pack_taken & btb_15_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_15_bht_T_4 = btb_15_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_15_bht_T_5 = io_i_branch_resolve_pack_taken & btb_15_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_15_bht_T_6 = btb_15_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_15_bht_T_7 = io_i_branch_resolve_pack_taken & btb_15_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_15_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_15_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_15_bht_T_13 = _btb_0_bht_T_8 & _btb_15_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_15_bht_T_16 = _btb_0_bht_T_8 & _btb_15_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_15_bht_T_19 = _btb_0_bht_T_8 & _btb_15_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_15_bht_T_20 = _btb_15_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_21 = _btb_15_bht_T_16 ? 2'h0 : _btb_15_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_22 = _btb_15_bht_T_13 ? 2'h0 : _btb_15_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_23 = _btb_15_bht_T_10 ? 2'h0 : _btb_15_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_24 = _btb_15_bht_T_7 ? 2'h3 : _btb_15_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_25 = _btb_15_bht_T_5 ? 2'h3 : _btb_15_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_26 = _btb_15_bht_T_3 ? 2'h3 : _btb_15_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_15_bht_T_27 = _btb_15_bht_T_1 ? 2'h1 : _btb_15_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8766 = btb_15_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6671; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8768 = btb_15_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_15_bht_T_27 : _GEN_8207; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_16_bht_T = btb_16_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_16_bht_T_1 = io_i_branch_resolve_pack_taken & btb_16_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_16_bht_T_2 = btb_16_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_16_bht_T_3 = io_i_branch_resolve_pack_taken & btb_16_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_16_bht_T_4 = btb_16_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_16_bht_T_5 = io_i_branch_resolve_pack_taken & btb_16_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_16_bht_T_6 = btb_16_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_16_bht_T_7 = io_i_branch_resolve_pack_taken & btb_16_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_16_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_16_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_16_bht_T_13 = _btb_0_bht_T_8 & _btb_16_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_16_bht_T_16 = _btb_0_bht_T_8 & _btb_16_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_16_bht_T_19 = _btb_0_bht_T_8 & _btb_16_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_16_bht_T_20 = _btb_16_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_21 = _btb_16_bht_T_16 ? 2'h0 : _btb_16_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_22 = _btb_16_bht_T_13 ? 2'h0 : _btb_16_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_23 = _btb_16_bht_T_10 ? 2'h0 : _btb_16_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_24 = _btb_16_bht_T_7 ? 2'h3 : _btb_16_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_25 = _btb_16_bht_T_5 ? 2'h3 : _btb_16_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_26 = _btb_16_bht_T_3 ? 2'h3 : _btb_16_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_16_bht_T_27 = _btb_16_bht_T_1 ? 2'h1 : _btb_16_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8770 = btb_16_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6672; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8772 = btb_16_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_16_bht_T_27 : _GEN_8208; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_17_bht_T = btb_17_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_17_bht_T_1 = io_i_branch_resolve_pack_taken & btb_17_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_17_bht_T_2 = btb_17_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_17_bht_T_3 = io_i_branch_resolve_pack_taken & btb_17_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_17_bht_T_4 = btb_17_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_17_bht_T_5 = io_i_branch_resolve_pack_taken & btb_17_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_17_bht_T_6 = btb_17_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_17_bht_T_7 = io_i_branch_resolve_pack_taken & btb_17_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_17_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_17_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_17_bht_T_13 = _btb_0_bht_T_8 & _btb_17_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_17_bht_T_16 = _btb_0_bht_T_8 & _btb_17_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_17_bht_T_19 = _btb_0_bht_T_8 & _btb_17_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_17_bht_T_20 = _btb_17_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_21 = _btb_17_bht_T_16 ? 2'h0 : _btb_17_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_22 = _btb_17_bht_T_13 ? 2'h0 : _btb_17_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_23 = _btb_17_bht_T_10 ? 2'h0 : _btb_17_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_24 = _btb_17_bht_T_7 ? 2'h3 : _btb_17_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_25 = _btb_17_bht_T_5 ? 2'h3 : _btb_17_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_26 = _btb_17_bht_T_3 ? 2'h3 : _btb_17_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_17_bht_T_27 = _btb_17_bht_T_1 ? 2'h1 : _btb_17_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8774 = btb_17_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6673; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8776 = btb_17_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_17_bht_T_27 : _GEN_8209; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_18_bht_T = btb_18_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_18_bht_T_1 = io_i_branch_resolve_pack_taken & btb_18_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_18_bht_T_2 = btb_18_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_18_bht_T_3 = io_i_branch_resolve_pack_taken & btb_18_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_18_bht_T_4 = btb_18_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_18_bht_T_5 = io_i_branch_resolve_pack_taken & btb_18_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_18_bht_T_6 = btb_18_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_18_bht_T_7 = io_i_branch_resolve_pack_taken & btb_18_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_18_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_18_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_18_bht_T_13 = _btb_0_bht_T_8 & _btb_18_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_18_bht_T_16 = _btb_0_bht_T_8 & _btb_18_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_18_bht_T_19 = _btb_0_bht_T_8 & _btb_18_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_18_bht_T_20 = _btb_18_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_21 = _btb_18_bht_T_16 ? 2'h0 : _btb_18_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_22 = _btb_18_bht_T_13 ? 2'h0 : _btb_18_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_23 = _btb_18_bht_T_10 ? 2'h0 : _btb_18_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_24 = _btb_18_bht_T_7 ? 2'h3 : _btb_18_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_25 = _btb_18_bht_T_5 ? 2'h3 : _btb_18_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_26 = _btb_18_bht_T_3 ? 2'h3 : _btb_18_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_18_bht_T_27 = _btb_18_bht_T_1 ? 2'h1 : _btb_18_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8778 = btb_18_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6674; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8780 = btb_18_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_18_bht_T_27 : _GEN_8210; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_19_bht_T = btb_19_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_19_bht_T_1 = io_i_branch_resolve_pack_taken & btb_19_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_19_bht_T_2 = btb_19_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_19_bht_T_3 = io_i_branch_resolve_pack_taken & btb_19_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_19_bht_T_4 = btb_19_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_19_bht_T_5 = io_i_branch_resolve_pack_taken & btb_19_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_19_bht_T_6 = btb_19_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_19_bht_T_7 = io_i_branch_resolve_pack_taken & btb_19_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_19_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_19_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_19_bht_T_13 = _btb_0_bht_T_8 & _btb_19_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_19_bht_T_16 = _btb_0_bht_T_8 & _btb_19_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_19_bht_T_19 = _btb_0_bht_T_8 & _btb_19_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_19_bht_T_20 = _btb_19_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_21 = _btb_19_bht_T_16 ? 2'h0 : _btb_19_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_22 = _btb_19_bht_T_13 ? 2'h0 : _btb_19_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_23 = _btb_19_bht_T_10 ? 2'h0 : _btb_19_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_24 = _btb_19_bht_T_7 ? 2'h3 : _btb_19_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_25 = _btb_19_bht_T_5 ? 2'h3 : _btb_19_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_26 = _btb_19_bht_T_3 ? 2'h3 : _btb_19_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_19_bht_T_27 = _btb_19_bht_T_1 ? 2'h1 : _btb_19_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8782 = btb_19_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6675; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8784 = btb_19_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_19_bht_T_27 : _GEN_8211; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_20_bht_T = btb_20_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_20_bht_T_1 = io_i_branch_resolve_pack_taken & btb_20_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_20_bht_T_2 = btb_20_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_20_bht_T_3 = io_i_branch_resolve_pack_taken & btb_20_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_20_bht_T_4 = btb_20_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_20_bht_T_5 = io_i_branch_resolve_pack_taken & btb_20_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_20_bht_T_6 = btb_20_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_20_bht_T_7 = io_i_branch_resolve_pack_taken & btb_20_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_20_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_20_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_20_bht_T_13 = _btb_0_bht_T_8 & _btb_20_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_20_bht_T_16 = _btb_0_bht_T_8 & _btb_20_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_20_bht_T_19 = _btb_0_bht_T_8 & _btb_20_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_20_bht_T_20 = _btb_20_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_21 = _btb_20_bht_T_16 ? 2'h0 : _btb_20_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_22 = _btb_20_bht_T_13 ? 2'h0 : _btb_20_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_23 = _btb_20_bht_T_10 ? 2'h0 : _btb_20_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_24 = _btb_20_bht_T_7 ? 2'h3 : _btb_20_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_25 = _btb_20_bht_T_5 ? 2'h3 : _btb_20_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_26 = _btb_20_bht_T_3 ? 2'h3 : _btb_20_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_20_bht_T_27 = _btb_20_bht_T_1 ? 2'h1 : _btb_20_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8786 = btb_20_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6676; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8788 = btb_20_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_20_bht_T_27 : _GEN_8212; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_21_bht_T = btb_21_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_21_bht_T_1 = io_i_branch_resolve_pack_taken & btb_21_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_21_bht_T_2 = btb_21_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_21_bht_T_3 = io_i_branch_resolve_pack_taken & btb_21_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_21_bht_T_4 = btb_21_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_21_bht_T_5 = io_i_branch_resolve_pack_taken & btb_21_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_21_bht_T_6 = btb_21_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_21_bht_T_7 = io_i_branch_resolve_pack_taken & btb_21_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_21_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_21_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_21_bht_T_13 = _btb_0_bht_T_8 & _btb_21_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_21_bht_T_16 = _btb_0_bht_T_8 & _btb_21_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_21_bht_T_19 = _btb_0_bht_T_8 & _btb_21_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_21_bht_T_20 = _btb_21_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_21 = _btb_21_bht_T_16 ? 2'h0 : _btb_21_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_22 = _btb_21_bht_T_13 ? 2'h0 : _btb_21_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_23 = _btb_21_bht_T_10 ? 2'h0 : _btb_21_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_24 = _btb_21_bht_T_7 ? 2'h3 : _btb_21_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_25 = _btb_21_bht_T_5 ? 2'h3 : _btb_21_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_26 = _btb_21_bht_T_3 ? 2'h3 : _btb_21_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_21_bht_T_27 = _btb_21_bht_T_1 ? 2'h1 : _btb_21_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8790 = btb_21_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6677; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8792 = btb_21_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_21_bht_T_27 : _GEN_8213; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_22_bht_T = btb_22_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_22_bht_T_1 = io_i_branch_resolve_pack_taken & btb_22_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_22_bht_T_2 = btb_22_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_22_bht_T_3 = io_i_branch_resolve_pack_taken & btb_22_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_22_bht_T_4 = btb_22_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_22_bht_T_5 = io_i_branch_resolve_pack_taken & btb_22_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_22_bht_T_6 = btb_22_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_22_bht_T_7 = io_i_branch_resolve_pack_taken & btb_22_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_22_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_22_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_22_bht_T_13 = _btb_0_bht_T_8 & _btb_22_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_22_bht_T_16 = _btb_0_bht_T_8 & _btb_22_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_22_bht_T_19 = _btb_0_bht_T_8 & _btb_22_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_22_bht_T_20 = _btb_22_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_21 = _btb_22_bht_T_16 ? 2'h0 : _btb_22_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_22 = _btb_22_bht_T_13 ? 2'h0 : _btb_22_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_23 = _btb_22_bht_T_10 ? 2'h0 : _btb_22_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_24 = _btb_22_bht_T_7 ? 2'h3 : _btb_22_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_25 = _btb_22_bht_T_5 ? 2'h3 : _btb_22_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_26 = _btb_22_bht_T_3 ? 2'h3 : _btb_22_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_22_bht_T_27 = _btb_22_bht_T_1 ? 2'h1 : _btb_22_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8794 = btb_22_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6678; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8796 = btb_22_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_22_bht_T_27 : _GEN_8214; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_23_bht_T = btb_23_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_23_bht_T_1 = io_i_branch_resolve_pack_taken & btb_23_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_23_bht_T_2 = btb_23_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_23_bht_T_3 = io_i_branch_resolve_pack_taken & btb_23_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_23_bht_T_4 = btb_23_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_23_bht_T_5 = io_i_branch_resolve_pack_taken & btb_23_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_23_bht_T_6 = btb_23_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_23_bht_T_7 = io_i_branch_resolve_pack_taken & btb_23_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_23_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_23_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_23_bht_T_13 = _btb_0_bht_T_8 & _btb_23_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_23_bht_T_16 = _btb_0_bht_T_8 & _btb_23_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_23_bht_T_19 = _btb_0_bht_T_8 & _btb_23_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_23_bht_T_20 = _btb_23_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_21 = _btb_23_bht_T_16 ? 2'h0 : _btb_23_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_22 = _btb_23_bht_T_13 ? 2'h0 : _btb_23_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_23 = _btb_23_bht_T_10 ? 2'h0 : _btb_23_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_24 = _btb_23_bht_T_7 ? 2'h3 : _btb_23_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_25 = _btb_23_bht_T_5 ? 2'h3 : _btb_23_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_26 = _btb_23_bht_T_3 ? 2'h3 : _btb_23_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_23_bht_T_27 = _btb_23_bht_T_1 ? 2'h1 : _btb_23_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8798 = btb_23_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6679; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8800 = btb_23_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_23_bht_T_27 : _GEN_8215; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_24_bht_T = btb_24_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_24_bht_T_1 = io_i_branch_resolve_pack_taken & btb_24_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_24_bht_T_2 = btb_24_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_24_bht_T_3 = io_i_branch_resolve_pack_taken & btb_24_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_24_bht_T_4 = btb_24_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_24_bht_T_5 = io_i_branch_resolve_pack_taken & btb_24_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_24_bht_T_6 = btb_24_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_24_bht_T_7 = io_i_branch_resolve_pack_taken & btb_24_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_24_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_24_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_24_bht_T_13 = _btb_0_bht_T_8 & _btb_24_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_24_bht_T_16 = _btb_0_bht_T_8 & _btb_24_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_24_bht_T_19 = _btb_0_bht_T_8 & _btb_24_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_24_bht_T_20 = _btb_24_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_21 = _btb_24_bht_T_16 ? 2'h0 : _btb_24_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_22 = _btb_24_bht_T_13 ? 2'h0 : _btb_24_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_23 = _btb_24_bht_T_10 ? 2'h0 : _btb_24_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_24 = _btb_24_bht_T_7 ? 2'h3 : _btb_24_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_25 = _btb_24_bht_T_5 ? 2'h3 : _btb_24_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_26 = _btb_24_bht_T_3 ? 2'h3 : _btb_24_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_24_bht_T_27 = _btb_24_bht_T_1 ? 2'h1 : _btb_24_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8802 = btb_24_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6680; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8804 = btb_24_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_24_bht_T_27 : _GEN_8216; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_25_bht_T = btb_25_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_25_bht_T_1 = io_i_branch_resolve_pack_taken & btb_25_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_25_bht_T_2 = btb_25_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_25_bht_T_3 = io_i_branch_resolve_pack_taken & btb_25_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_25_bht_T_4 = btb_25_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_25_bht_T_5 = io_i_branch_resolve_pack_taken & btb_25_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_25_bht_T_6 = btb_25_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_25_bht_T_7 = io_i_branch_resolve_pack_taken & btb_25_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_25_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_25_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_25_bht_T_13 = _btb_0_bht_T_8 & _btb_25_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_25_bht_T_16 = _btb_0_bht_T_8 & _btb_25_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_25_bht_T_19 = _btb_0_bht_T_8 & _btb_25_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_25_bht_T_20 = _btb_25_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_21 = _btb_25_bht_T_16 ? 2'h0 : _btb_25_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_22 = _btb_25_bht_T_13 ? 2'h0 : _btb_25_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_23 = _btb_25_bht_T_10 ? 2'h0 : _btb_25_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_24 = _btb_25_bht_T_7 ? 2'h3 : _btb_25_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_25 = _btb_25_bht_T_5 ? 2'h3 : _btb_25_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_26 = _btb_25_bht_T_3 ? 2'h3 : _btb_25_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_25_bht_T_27 = _btb_25_bht_T_1 ? 2'h1 : _btb_25_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8806 = btb_25_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6681; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8808 = btb_25_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_25_bht_T_27 : _GEN_8217; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_26_bht_T = btb_26_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_26_bht_T_1 = io_i_branch_resolve_pack_taken & btb_26_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_26_bht_T_2 = btb_26_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_26_bht_T_3 = io_i_branch_resolve_pack_taken & btb_26_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_26_bht_T_4 = btb_26_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_26_bht_T_5 = io_i_branch_resolve_pack_taken & btb_26_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_26_bht_T_6 = btb_26_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_26_bht_T_7 = io_i_branch_resolve_pack_taken & btb_26_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_26_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_26_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_26_bht_T_13 = _btb_0_bht_T_8 & _btb_26_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_26_bht_T_16 = _btb_0_bht_T_8 & _btb_26_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_26_bht_T_19 = _btb_0_bht_T_8 & _btb_26_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_26_bht_T_20 = _btb_26_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_21 = _btb_26_bht_T_16 ? 2'h0 : _btb_26_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_22 = _btb_26_bht_T_13 ? 2'h0 : _btb_26_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_23 = _btb_26_bht_T_10 ? 2'h0 : _btb_26_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_24 = _btb_26_bht_T_7 ? 2'h3 : _btb_26_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_25 = _btb_26_bht_T_5 ? 2'h3 : _btb_26_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_26 = _btb_26_bht_T_3 ? 2'h3 : _btb_26_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_26_bht_T_27 = _btb_26_bht_T_1 ? 2'h1 : _btb_26_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8810 = btb_26_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6682; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8812 = btb_26_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_26_bht_T_27 : _GEN_8218; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_27_bht_T = btb_27_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_27_bht_T_1 = io_i_branch_resolve_pack_taken & btb_27_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_27_bht_T_2 = btb_27_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_27_bht_T_3 = io_i_branch_resolve_pack_taken & btb_27_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_27_bht_T_4 = btb_27_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_27_bht_T_5 = io_i_branch_resolve_pack_taken & btb_27_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_27_bht_T_6 = btb_27_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_27_bht_T_7 = io_i_branch_resolve_pack_taken & btb_27_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_27_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_27_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_27_bht_T_13 = _btb_0_bht_T_8 & _btb_27_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_27_bht_T_16 = _btb_0_bht_T_8 & _btb_27_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_27_bht_T_19 = _btb_0_bht_T_8 & _btb_27_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_27_bht_T_20 = _btb_27_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_21 = _btb_27_bht_T_16 ? 2'h0 : _btb_27_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_22 = _btb_27_bht_T_13 ? 2'h0 : _btb_27_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_23 = _btb_27_bht_T_10 ? 2'h0 : _btb_27_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_24 = _btb_27_bht_T_7 ? 2'h3 : _btb_27_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_25 = _btb_27_bht_T_5 ? 2'h3 : _btb_27_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_26 = _btb_27_bht_T_3 ? 2'h3 : _btb_27_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_27_bht_T_27 = _btb_27_bht_T_1 ? 2'h1 : _btb_27_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8814 = btb_27_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6683; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8816 = btb_27_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_27_bht_T_27 : _GEN_8219; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_28_bht_T = btb_28_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_28_bht_T_1 = io_i_branch_resolve_pack_taken & btb_28_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_28_bht_T_2 = btb_28_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_28_bht_T_3 = io_i_branch_resolve_pack_taken & btb_28_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_28_bht_T_4 = btb_28_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_28_bht_T_5 = io_i_branch_resolve_pack_taken & btb_28_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_28_bht_T_6 = btb_28_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_28_bht_T_7 = io_i_branch_resolve_pack_taken & btb_28_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_28_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_28_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_28_bht_T_13 = _btb_0_bht_T_8 & _btb_28_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_28_bht_T_16 = _btb_0_bht_T_8 & _btb_28_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_28_bht_T_19 = _btb_0_bht_T_8 & _btb_28_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_28_bht_T_20 = _btb_28_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_21 = _btb_28_bht_T_16 ? 2'h0 : _btb_28_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_22 = _btb_28_bht_T_13 ? 2'h0 : _btb_28_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_23 = _btb_28_bht_T_10 ? 2'h0 : _btb_28_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_24 = _btb_28_bht_T_7 ? 2'h3 : _btb_28_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_25 = _btb_28_bht_T_5 ? 2'h3 : _btb_28_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_26 = _btb_28_bht_T_3 ? 2'h3 : _btb_28_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_28_bht_T_27 = _btb_28_bht_T_1 ? 2'h1 : _btb_28_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8818 = btb_28_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6684; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8820 = btb_28_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_28_bht_T_27 : _GEN_8220; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_29_bht_T = btb_29_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_29_bht_T_1 = io_i_branch_resolve_pack_taken & btb_29_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_29_bht_T_2 = btb_29_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_29_bht_T_3 = io_i_branch_resolve_pack_taken & btb_29_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_29_bht_T_4 = btb_29_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_29_bht_T_5 = io_i_branch_resolve_pack_taken & btb_29_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_29_bht_T_6 = btb_29_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_29_bht_T_7 = io_i_branch_resolve_pack_taken & btb_29_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_29_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_29_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_29_bht_T_13 = _btb_0_bht_T_8 & _btb_29_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_29_bht_T_16 = _btb_0_bht_T_8 & _btb_29_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_29_bht_T_19 = _btb_0_bht_T_8 & _btb_29_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_29_bht_T_20 = _btb_29_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_21 = _btb_29_bht_T_16 ? 2'h0 : _btb_29_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_22 = _btb_29_bht_T_13 ? 2'h0 : _btb_29_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_23 = _btb_29_bht_T_10 ? 2'h0 : _btb_29_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_24 = _btb_29_bht_T_7 ? 2'h3 : _btb_29_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_25 = _btb_29_bht_T_5 ? 2'h3 : _btb_29_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_26 = _btb_29_bht_T_3 ? 2'h3 : _btb_29_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_29_bht_T_27 = _btb_29_bht_T_1 ? 2'h1 : _btb_29_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_8821 = btb_29_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_28_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_27_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_26_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_25_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_24_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_23_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_22_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_21_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_20_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_19_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_18_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_17_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_16_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_15_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_8761)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_8822 = btb_29_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6685; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8824 = btb_29_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_29_bht_T_27 : _GEN_8221; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_30_bht_T = btb_30_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_30_bht_T_1 = io_i_branch_resolve_pack_taken & btb_30_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_30_bht_T_2 = btb_30_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_30_bht_T_3 = io_i_branch_resolve_pack_taken & btb_30_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_30_bht_T_4 = btb_30_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_30_bht_T_5 = io_i_branch_resolve_pack_taken & btb_30_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_30_bht_T_6 = btb_30_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_30_bht_T_7 = io_i_branch_resolve_pack_taken & btb_30_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_30_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_30_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_30_bht_T_13 = _btb_0_bht_T_8 & _btb_30_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_30_bht_T_16 = _btb_0_bht_T_8 & _btb_30_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_30_bht_T_19 = _btb_0_bht_T_8 & _btb_30_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_30_bht_T_20 = _btb_30_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_21 = _btb_30_bht_T_16 ? 2'h0 : _btb_30_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_22 = _btb_30_bht_T_13 ? 2'h0 : _btb_30_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_23 = _btb_30_bht_T_10 ? 2'h0 : _btb_30_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_24 = _btb_30_bht_T_7 ? 2'h3 : _btb_30_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_25 = _btb_30_bht_T_5 ? 2'h3 : _btb_30_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_26 = _btb_30_bht_T_3 ? 2'h3 : _btb_30_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_30_bht_T_27 = _btb_30_bht_T_1 ? 2'h1 : _btb_30_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8826 = btb_30_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6686; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8828 = btb_30_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_30_bht_T_27 : _GEN_8222; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_31_bht_T = btb_31_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_31_bht_T_1 = io_i_branch_resolve_pack_taken & btb_31_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_31_bht_T_2 = btb_31_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_31_bht_T_3 = io_i_branch_resolve_pack_taken & btb_31_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_31_bht_T_4 = btb_31_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_31_bht_T_5 = io_i_branch_resolve_pack_taken & btb_31_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_31_bht_T_6 = btb_31_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_31_bht_T_7 = io_i_branch_resolve_pack_taken & btb_31_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_31_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_31_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_31_bht_T_13 = _btb_0_bht_T_8 & _btb_31_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_31_bht_T_16 = _btb_0_bht_T_8 & _btb_31_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_31_bht_T_19 = _btb_0_bht_T_8 & _btb_31_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_31_bht_T_20 = _btb_31_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_21 = _btb_31_bht_T_16 ? 2'h0 : _btb_31_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_22 = _btb_31_bht_T_13 ? 2'h0 : _btb_31_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_23 = _btb_31_bht_T_10 ? 2'h0 : _btb_31_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_24 = _btb_31_bht_T_7 ? 2'h3 : _btb_31_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_25 = _btb_31_bht_T_5 ? 2'h3 : _btb_31_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_26 = _btb_31_bht_T_3 ? 2'h3 : _btb_31_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_31_bht_T_27 = _btb_31_bht_T_1 ? 2'h1 : _btb_31_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8830 = btb_31_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6687; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8832 = btb_31_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_31_bht_T_27 : _GEN_8223; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_32_bht_T = btb_32_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_32_bht_T_1 = io_i_branch_resolve_pack_taken & btb_32_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_32_bht_T_2 = btb_32_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_32_bht_T_3 = io_i_branch_resolve_pack_taken & btb_32_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_32_bht_T_4 = btb_32_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_32_bht_T_5 = io_i_branch_resolve_pack_taken & btb_32_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_32_bht_T_6 = btb_32_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_32_bht_T_7 = io_i_branch_resolve_pack_taken & btb_32_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_32_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_32_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_32_bht_T_13 = _btb_0_bht_T_8 & _btb_32_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_32_bht_T_16 = _btb_0_bht_T_8 & _btb_32_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_32_bht_T_19 = _btb_0_bht_T_8 & _btb_32_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_32_bht_T_20 = _btb_32_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_21 = _btb_32_bht_T_16 ? 2'h0 : _btb_32_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_22 = _btb_32_bht_T_13 ? 2'h0 : _btb_32_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_23 = _btb_32_bht_T_10 ? 2'h0 : _btb_32_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_24 = _btb_32_bht_T_7 ? 2'h3 : _btb_32_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_25 = _btb_32_bht_T_5 ? 2'h3 : _btb_32_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_26 = _btb_32_bht_T_3 ? 2'h3 : _btb_32_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_32_bht_T_27 = _btb_32_bht_T_1 ? 2'h1 : _btb_32_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8834 = btb_32_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6688; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8836 = btb_32_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_32_bht_T_27 : _GEN_8224; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_33_bht_T = btb_33_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_33_bht_T_1 = io_i_branch_resolve_pack_taken & btb_33_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_33_bht_T_2 = btb_33_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_33_bht_T_3 = io_i_branch_resolve_pack_taken & btb_33_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_33_bht_T_4 = btb_33_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_33_bht_T_5 = io_i_branch_resolve_pack_taken & btb_33_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_33_bht_T_6 = btb_33_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_33_bht_T_7 = io_i_branch_resolve_pack_taken & btb_33_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_33_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_33_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_33_bht_T_13 = _btb_0_bht_T_8 & _btb_33_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_33_bht_T_16 = _btb_0_bht_T_8 & _btb_33_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_33_bht_T_19 = _btb_0_bht_T_8 & _btb_33_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_33_bht_T_20 = _btb_33_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_21 = _btb_33_bht_T_16 ? 2'h0 : _btb_33_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_22 = _btb_33_bht_T_13 ? 2'h0 : _btb_33_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_23 = _btb_33_bht_T_10 ? 2'h0 : _btb_33_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_24 = _btb_33_bht_T_7 ? 2'h3 : _btb_33_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_25 = _btb_33_bht_T_5 ? 2'h3 : _btb_33_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_26 = _btb_33_bht_T_3 ? 2'h3 : _btb_33_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_33_bht_T_27 = _btb_33_bht_T_1 ? 2'h1 : _btb_33_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8838 = btb_33_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6689; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8840 = btb_33_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_33_bht_T_27 : _GEN_8225; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_34_bht_T = btb_34_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_34_bht_T_1 = io_i_branch_resolve_pack_taken & btb_34_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_34_bht_T_2 = btb_34_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_34_bht_T_3 = io_i_branch_resolve_pack_taken & btb_34_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_34_bht_T_4 = btb_34_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_34_bht_T_5 = io_i_branch_resolve_pack_taken & btb_34_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_34_bht_T_6 = btb_34_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_34_bht_T_7 = io_i_branch_resolve_pack_taken & btb_34_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_34_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_34_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_34_bht_T_13 = _btb_0_bht_T_8 & _btb_34_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_34_bht_T_16 = _btb_0_bht_T_8 & _btb_34_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_34_bht_T_19 = _btb_0_bht_T_8 & _btb_34_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_34_bht_T_20 = _btb_34_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_21 = _btb_34_bht_T_16 ? 2'h0 : _btb_34_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_22 = _btb_34_bht_T_13 ? 2'h0 : _btb_34_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_23 = _btb_34_bht_T_10 ? 2'h0 : _btb_34_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_24 = _btb_34_bht_T_7 ? 2'h3 : _btb_34_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_25 = _btb_34_bht_T_5 ? 2'h3 : _btb_34_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_26 = _btb_34_bht_T_3 ? 2'h3 : _btb_34_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_34_bht_T_27 = _btb_34_bht_T_1 ? 2'h1 : _btb_34_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8842 = btb_34_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6690; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8844 = btb_34_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_34_bht_T_27 : _GEN_8226; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_35_bht_T = btb_35_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_35_bht_T_1 = io_i_branch_resolve_pack_taken & btb_35_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_35_bht_T_2 = btb_35_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_35_bht_T_3 = io_i_branch_resolve_pack_taken & btb_35_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_35_bht_T_4 = btb_35_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_35_bht_T_5 = io_i_branch_resolve_pack_taken & btb_35_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_35_bht_T_6 = btb_35_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_35_bht_T_7 = io_i_branch_resolve_pack_taken & btb_35_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_35_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_35_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_35_bht_T_13 = _btb_0_bht_T_8 & _btb_35_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_35_bht_T_16 = _btb_0_bht_T_8 & _btb_35_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_35_bht_T_19 = _btb_0_bht_T_8 & _btb_35_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_35_bht_T_20 = _btb_35_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_21 = _btb_35_bht_T_16 ? 2'h0 : _btb_35_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_22 = _btb_35_bht_T_13 ? 2'h0 : _btb_35_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_23 = _btb_35_bht_T_10 ? 2'h0 : _btb_35_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_24 = _btb_35_bht_T_7 ? 2'h3 : _btb_35_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_25 = _btb_35_bht_T_5 ? 2'h3 : _btb_35_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_26 = _btb_35_bht_T_3 ? 2'h3 : _btb_35_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_35_bht_T_27 = _btb_35_bht_T_1 ? 2'h1 : _btb_35_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8846 = btb_35_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6691; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8848 = btb_35_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_35_bht_T_27 : _GEN_8227; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_36_bht_T = btb_36_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_36_bht_T_1 = io_i_branch_resolve_pack_taken & btb_36_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_36_bht_T_2 = btb_36_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_36_bht_T_3 = io_i_branch_resolve_pack_taken & btb_36_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_36_bht_T_4 = btb_36_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_36_bht_T_5 = io_i_branch_resolve_pack_taken & btb_36_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_36_bht_T_6 = btb_36_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_36_bht_T_7 = io_i_branch_resolve_pack_taken & btb_36_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_36_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_36_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_36_bht_T_13 = _btb_0_bht_T_8 & _btb_36_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_36_bht_T_16 = _btb_0_bht_T_8 & _btb_36_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_36_bht_T_19 = _btb_0_bht_T_8 & _btb_36_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_36_bht_T_20 = _btb_36_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_21 = _btb_36_bht_T_16 ? 2'h0 : _btb_36_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_22 = _btb_36_bht_T_13 ? 2'h0 : _btb_36_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_23 = _btb_36_bht_T_10 ? 2'h0 : _btb_36_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_24 = _btb_36_bht_T_7 ? 2'h3 : _btb_36_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_25 = _btb_36_bht_T_5 ? 2'h3 : _btb_36_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_26 = _btb_36_bht_T_3 ? 2'h3 : _btb_36_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_36_bht_T_27 = _btb_36_bht_T_1 ? 2'h1 : _btb_36_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8850 = btb_36_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6692; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8852 = btb_36_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_36_bht_T_27 : _GEN_8228; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_37_bht_T = btb_37_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_37_bht_T_1 = io_i_branch_resolve_pack_taken & btb_37_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_37_bht_T_2 = btb_37_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_37_bht_T_3 = io_i_branch_resolve_pack_taken & btb_37_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_37_bht_T_4 = btb_37_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_37_bht_T_5 = io_i_branch_resolve_pack_taken & btb_37_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_37_bht_T_6 = btb_37_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_37_bht_T_7 = io_i_branch_resolve_pack_taken & btb_37_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_37_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_37_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_37_bht_T_13 = _btb_0_bht_T_8 & _btb_37_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_37_bht_T_16 = _btb_0_bht_T_8 & _btb_37_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_37_bht_T_19 = _btb_0_bht_T_8 & _btb_37_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_37_bht_T_20 = _btb_37_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_21 = _btb_37_bht_T_16 ? 2'h0 : _btb_37_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_22 = _btb_37_bht_T_13 ? 2'h0 : _btb_37_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_23 = _btb_37_bht_T_10 ? 2'h0 : _btb_37_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_24 = _btb_37_bht_T_7 ? 2'h3 : _btb_37_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_25 = _btb_37_bht_T_5 ? 2'h3 : _btb_37_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_26 = _btb_37_bht_T_3 ? 2'h3 : _btb_37_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_37_bht_T_27 = _btb_37_bht_T_1 ? 2'h1 : _btb_37_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8854 = btb_37_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6693; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8856 = btb_37_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_37_bht_T_27 : _GEN_8229; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_38_bht_T = btb_38_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_38_bht_T_1 = io_i_branch_resolve_pack_taken & btb_38_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_38_bht_T_2 = btb_38_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_38_bht_T_3 = io_i_branch_resolve_pack_taken & btb_38_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_38_bht_T_4 = btb_38_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_38_bht_T_5 = io_i_branch_resolve_pack_taken & btb_38_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_38_bht_T_6 = btb_38_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_38_bht_T_7 = io_i_branch_resolve_pack_taken & btb_38_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_38_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_38_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_38_bht_T_13 = _btb_0_bht_T_8 & _btb_38_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_38_bht_T_16 = _btb_0_bht_T_8 & _btb_38_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_38_bht_T_19 = _btb_0_bht_T_8 & _btb_38_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_38_bht_T_20 = _btb_38_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_21 = _btb_38_bht_T_16 ? 2'h0 : _btb_38_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_22 = _btb_38_bht_T_13 ? 2'h0 : _btb_38_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_23 = _btb_38_bht_T_10 ? 2'h0 : _btb_38_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_24 = _btb_38_bht_T_7 ? 2'h3 : _btb_38_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_25 = _btb_38_bht_T_5 ? 2'h3 : _btb_38_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_26 = _btb_38_bht_T_3 ? 2'h3 : _btb_38_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_38_bht_T_27 = _btb_38_bht_T_1 ? 2'h1 : _btb_38_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8858 = btb_38_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6694; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8860 = btb_38_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_38_bht_T_27 : _GEN_8230; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_39_bht_T = btb_39_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_39_bht_T_1 = io_i_branch_resolve_pack_taken & btb_39_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_39_bht_T_2 = btb_39_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_39_bht_T_3 = io_i_branch_resolve_pack_taken & btb_39_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_39_bht_T_4 = btb_39_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_39_bht_T_5 = io_i_branch_resolve_pack_taken & btb_39_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_39_bht_T_6 = btb_39_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_39_bht_T_7 = io_i_branch_resolve_pack_taken & btb_39_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_39_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_39_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_39_bht_T_13 = _btb_0_bht_T_8 & _btb_39_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_39_bht_T_16 = _btb_0_bht_T_8 & _btb_39_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_39_bht_T_19 = _btb_0_bht_T_8 & _btb_39_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_39_bht_T_20 = _btb_39_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_21 = _btb_39_bht_T_16 ? 2'h0 : _btb_39_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_22 = _btb_39_bht_T_13 ? 2'h0 : _btb_39_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_23 = _btb_39_bht_T_10 ? 2'h0 : _btb_39_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_24 = _btb_39_bht_T_7 ? 2'h3 : _btb_39_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_25 = _btb_39_bht_T_5 ? 2'h3 : _btb_39_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_26 = _btb_39_bht_T_3 ? 2'h3 : _btb_39_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_39_bht_T_27 = _btb_39_bht_T_1 ? 2'h1 : _btb_39_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8862 = btb_39_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6695; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8864 = btb_39_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_39_bht_T_27 : _GEN_8231; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_40_bht_T = btb_40_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_40_bht_T_1 = io_i_branch_resolve_pack_taken & btb_40_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_40_bht_T_2 = btb_40_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_40_bht_T_3 = io_i_branch_resolve_pack_taken & btb_40_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_40_bht_T_4 = btb_40_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_40_bht_T_5 = io_i_branch_resolve_pack_taken & btb_40_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_40_bht_T_6 = btb_40_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_40_bht_T_7 = io_i_branch_resolve_pack_taken & btb_40_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_40_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_40_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_40_bht_T_13 = _btb_0_bht_T_8 & _btb_40_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_40_bht_T_16 = _btb_0_bht_T_8 & _btb_40_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_40_bht_T_19 = _btb_0_bht_T_8 & _btb_40_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_40_bht_T_20 = _btb_40_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_21 = _btb_40_bht_T_16 ? 2'h0 : _btb_40_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_22 = _btb_40_bht_T_13 ? 2'h0 : _btb_40_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_23 = _btb_40_bht_T_10 ? 2'h0 : _btb_40_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_24 = _btb_40_bht_T_7 ? 2'h3 : _btb_40_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_25 = _btb_40_bht_T_5 ? 2'h3 : _btb_40_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_26 = _btb_40_bht_T_3 ? 2'h3 : _btb_40_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_40_bht_T_27 = _btb_40_bht_T_1 ? 2'h1 : _btb_40_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8866 = btb_40_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6696; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8868 = btb_40_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_40_bht_T_27 : _GEN_8232; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_41_bht_T = btb_41_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_41_bht_T_1 = io_i_branch_resolve_pack_taken & btb_41_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_41_bht_T_2 = btb_41_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_41_bht_T_3 = io_i_branch_resolve_pack_taken & btb_41_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_41_bht_T_4 = btb_41_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_41_bht_T_5 = io_i_branch_resolve_pack_taken & btb_41_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_41_bht_T_6 = btb_41_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_41_bht_T_7 = io_i_branch_resolve_pack_taken & btb_41_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_41_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_41_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_41_bht_T_13 = _btb_0_bht_T_8 & _btb_41_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_41_bht_T_16 = _btb_0_bht_T_8 & _btb_41_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_41_bht_T_19 = _btb_0_bht_T_8 & _btb_41_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_41_bht_T_20 = _btb_41_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_21 = _btb_41_bht_T_16 ? 2'h0 : _btb_41_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_22 = _btb_41_bht_T_13 ? 2'h0 : _btb_41_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_23 = _btb_41_bht_T_10 ? 2'h0 : _btb_41_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_24 = _btb_41_bht_T_7 ? 2'h3 : _btb_41_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_25 = _btb_41_bht_T_5 ? 2'h3 : _btb_41_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_26 = _btb_41_bht_T_3 ? 2'h3 : _btb_41_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_41_bht_T_27 = _btb_41_bht_T_1 ? 2'h1 : _btb_41_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8870 = btb_41_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6697; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8872 = btb_41_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_41_bht_T_27 : _GEN_8233; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_42_bht_T = btb_42_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_42_bht_T_1 = io_i_branch_resolve_pack_taken & btb_42_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_42_bht_T_2 = btb_42_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_42_bht_T_3 = io_i_branch_resolve_pack_taken & btb_42_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_42_bht_T_4 = btb_42_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_42_bht_T_5 = io_i_branch_resolve_pack_taken & btb_42_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_42_bht_T_6 = btb_42_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_42_bht_T_7 = io_i_branch_resolve_pack_taken & btb_42_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_42_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_42_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_42_bht_T_13 = _btb_0_bht_T_8 & _btb_42_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_42_bht_T_16 = _btb_0_bht_T_8 & _btb_42_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_42_bht_T_19 = _btb_0_bht_T_8 & _btb_42_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_42_bht_T_20 = _btb_42_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_21 = _btb_42_bht_T_16 ? 2'h0 : _btb_42_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_22 = _btb_42_bht_T_13 ? 2'h0 : _btb_42_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_23 = _btb_42_bht_T_10 ? 2'h0 : _btb_42_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_24 = _btb_42_bht_T_7 ? 2'h3 : _btb_42_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_25 = _btb_42_bht_T_5 ? 2'h3 : _btb_42_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_26 = _btb_42_bht_T_3 ? 2'h3 : _btb_42_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_42_bht_T_27 = _btb_42_bht_T_1 ? 2'h1 : _btb_42_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8874 = btb_42_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6698; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8876 = btb_42_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_42_bht_T_27 : _GEN_8234; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_43_bht_T = btb_43_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_43_bht_T_1 = io_i_branch_resolve_pack_taken & btb_43_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_43_bht_T_2 = btb_43_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_43_bht_T_3 = io_i_branch_resolve_pack_taken & btb_43_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_43_bht_T_4 = btb_43_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_43_bht_T_5 = io_i_branch_resolve_pack_taken & btb_43_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_43_bht_T_6 = btb_43_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_43_bht_T_7 = io_i_branch_resolve_pack_taken & btb_43_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_43_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_43_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_43_bht_T_13 = _btb_0_bht_T_8 & _btb_43_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_43_bht_T_16 = _btb_0_bht_T_8 & _btb_43_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_43_bht_T_19 = _btb_0_bht_T_8 & _btb_43_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_43_bht_T_20 = _btb_43_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_21 = _btb_43_bht_T_16 ? 2'h0 : _btb_43_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_22 = _btb_43_bht_T_13 ? 2'h0 : _btb_43_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_23 = _btb_43_bht_T_10 ? 2'h0 : _btb_43_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_24 = _btb_43_bht_T_7 ? 2'h3 : _btb_43_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_25 = _btb_43_bht_T_5 ? 2'h3 : _btb_43_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_26 = _btb_43_bht_T_3 ? 2'h3 : _btb_43_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_43_bht_T_27 = _btb_43_bht_T_1 ? 2'h1 : _btb_43_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8878 = btb_43_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6699; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8880 = btb_43_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_43_bht_T_27 : _GEN_8235; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_44_bht_T = btb_44_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_44_bht_T_1 = io_i_branch_resolve_pack_taken & btb_44_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_44_bht_T_2 = btb_44_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_44_bht_T_3 = io_i_branch_resolve_pack_taken & btb_44_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_44_bht_T_4 = btb_44_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_44_bht_T_5 = io_i_branch_resolve_pack_taken & btb_44_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_44_bht_T_6 = btb_44_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_44_bht_T_7 = io_i_branch_resolve_pack_taken & btb_44_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_44_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_44_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_44_bht_T_13 = _btb_0_bht_T_8 & _btb_44_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_44_bht_T_16 = _btb_0_bht_T_8 & _btb_44_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_44_bht_T_19 = _btb_0_bht_T_8 & _btb_44_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_44_bht_T_20 = _btb_44_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_21 = _btb_44_bht_T_16 ? 2'h0 : _btb_44_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_22 = _btb_44_bht_T_13 ? 2'h0 : _btb_44_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_23 = _btb_44_bht_T_10 ? 2'h0 : _btb_44_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_24 = _btb_44_bht_T_7 ? 2'h3 : _btb_44_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_25 = _btb_44_bht_T_5 ? 2'h3 : _btb_44_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_26 = _btb_44_bht_T_3 ? 2'h3 : _btb_44_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_44_bht_T_27 = _btb_44_bht_T_1 ? 2'h1 : _btb_44_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_8881 = btb_44_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_43_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_42_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_41_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_40_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_39_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_38_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_37_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_36_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_35_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_34_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_33_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_32_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_31_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_30_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_8821)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_8882 = btb_44_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6700; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8884 = btb_44_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_44_bht_T_27 : _GEN_8236; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_45_bht_T = btb_45_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_45_bht_T_1 = io_i_branch_resolve_pack_taken & btb_45_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_45_bht_T_2 = btb_45_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_45_bht_T_3 = io_i_branch_resolve_pack_taken & btb_45_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_45_bht_T_4 = btb_45_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_45_bht_T_5 = io_i_branch_resolve_pack_taken & btb_45_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_45_bht_T_6 = btb_45_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_45_bht_T_7 = io_i_branch_resolve_pack_taken & btb_45_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_45_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_45_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_45_bht_T_13 = _btb_0_bht_T_8 & _btb_45_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_45_bht_T_16 = _btb_0_bht_T_8 & _btb_45_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_45_bht_T_19 = _btb_0_bht_T_8 & _btb_45_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_45_bht_T_20 = _btb_45_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_21 = _btb_45_bht_T_16 ? 2'h0 : _btb_45_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_22 = _btb_45_bht_T_13 ? 2'h0 : _btb_45_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_23 = _btb_45_bht_T_10 ? 2'h0 : _btb_45_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_24 = _btb_45_bht_T_7 ? 2'h3 : _btb_45_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_25 = _btb_45_bht_T_5 ? 2'h3 : _btb_45_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_26 = _btb_45_bht_T_3 ? 2'h3 : _btb_45_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_45_bht_T_27 = _btb_45_bht_T_1 ? 2'h1 : _btb_45_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8886 = btb_45_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6701; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8888 = btb_45_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_45_bht_T_27 : _GEN_8237; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_46_bht_T = btb_46_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_46_bht_T_1 = io_i_branch_resolve_pack_taken & btb_46_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_46_bht_T_2 = btb_46_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_46_bht_T_3 = io_i_branch_resolve_pack_taken & btb_46_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_46_bht_T_4 = btb_46_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_46_bht_T_5 = io_i_branch_resolve_pack_taken & btb_46_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_46_bht_T_6 = btb_46_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_46_bht_T_7 = io_i_branch_resolve_pack_taken & btb_46_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_46_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_46_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_46_bht_T_13 = _btb_0_bht_T_8 & _btb_46_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_46_bht_T_16 = _btb_0_bht_T_8 & _btb_46_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_46_bht_T_19 = _btb_0_bht_T_8 & _btb_46_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_46_bht_T_20 = _btb_46_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_21 = _btb_46_bht_T_16 ? 2'h0 : _btb_46_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_22 = _btb_46_bht_T_13 ? 2'h0 : _btb_46_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_23 = _btb_46_bht_T_10 ? 2'h0 : _btb_46_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_24 = _btb_46_bht_T_7 ? 2'h3 : _btb_46_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_25 = _btb_46_bht_T_5 ? 2'h3 : _btb_46_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_26 = _btb_46_bht_T_3 ? 2'h3 : _btb_46_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_46_bht_T_27 = _btb_46_bht_T_1 ? 2'h1 : _btb_46_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8890 = btb_46_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6702; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8892 = btb_46_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_46_bht_T_27 : _GEN_8238; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_47_bht_T = btb_47_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_47_bht_T_1 = io_i_branch_resolve_pack_taken & btb_47_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_47_bht_T_2 = btb_47_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_47_bht_T_3 = io_i_branch_resolve_pack_taken & btb_47_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_47_bht_T_4 = btb_47_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_47_bht_T_5 = io_i_branch_resolve_pack_taken & btb_47_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_47_bht_T_6 = btb_47_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_47_bht_T_7 = io_i_branch_resolve_pack_taken & btb_47_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_47_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_47_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_47_bht_T_13 = _btb_0_bht_T_8 & _btb_47_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_47_bht_T_16 = _btb_0_bht_T_8 & _btb_47_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_47_bht_T_19 = _btb_0_bht_T_8 & _btb_47_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_47_bht_T_20 = _btb_47_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_21 = _btb_47_bht_T_16 ? 2'h0 : _btb_47_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_22 = _btb_47_bht_T_13 ? 2'h0 : _btb_47_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_23 = _btb_47_bht_T_10 ? 2'h0 : _btb_47_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_24 = _btb_47_bht_T_7 ? 2'h3 : _btb_47_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_25 = _btb_47_bht_T_5 ? 2'h3 : _btb_47_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_26 = _btb_47_bht_T_3 ? 2'h3 : _btb_47_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_47_bht_T_27 = _btb_47_bht_T_1 ? 2'h1 : _btb_47_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8894 = btb_47_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6703; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8896 = btb_47_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_47_bht_T_27 : _GEN_8239; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_48_bht_T = btb_48_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_48_bht_T_1 = io_i_branch_resolve_pack_taken & btb_48_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_48_bht_T_2 = btb_48_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_48_bht_T_3 = io_i_branch_resolve_pack_taken & btb_48_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_48_bht_T_4 = btb_48_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_48_bht_T_5 = io_i_branch_resolve_pack_taken & btb_48_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_48_bht_T_6 = btb_48_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_48_bht_T_7 = io_i_branch_resolve_pack_taken & btb_48_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_48_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_48_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_48_bht_T_13 = _btb_0_bht_T_8 & _btb_48_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_48_bht_T_16 = _btb_0_bht_T_8 & _btb_48_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_48_bht_T_19 = _btb_0_bht_T_8 & _btb_48_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_48_bht_T_20 = _btb_48_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_21 = _btb_48_bht_T_16 ? 2'h0 : _btb_48_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_22 = _btb_48_bht_T_13 ? 2'h0 : _btb_48_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_23 = _btb_48_bht_T_10 ? 2'h0 : _btb_48_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_24 = _btb_48_bht_T_7 ? 2'h3 : _btb_48_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_25 = _btb_48_bht_T_5 ? 2'h3 : _btb_48_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_26 = _btb_48_bht_T_3 ? 2'h3 : _btb_48_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_48_bht_T_27 = _btb_48_bht_T_1 ? 2'h1 : _btb_48_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8898 = btb_48_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6704; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8900 = btb_48_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_48_bht_T_27 : _GEN_8240; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_49_bht_T = btb_49_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_49_bht_T_1 = io_i_branch_resolve_pack_taken & btb_49_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_49_bht_T_2 = btb_49_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_49_bht_T_3 = io_i_branch_resolve_pack_taken & btb_49_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_49_bht_T_4 = btb_49_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_49_bht_T_5 = io_i_branch_resolve_pack_taken & btb_49_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_49_bht_T_6 = btb_49_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_49_bht_T_7 = io_i_branch_resolve_pack_taken & btb_49_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_49_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_49_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_49_bht_T_13 = _btb_0_bht_T_8 & _btb_49_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_49_bht_T_16 = _btb_0_bht_T_8 & _btb_49_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_49_bht_T_19 = _btb_0_bht_T_8 & _btb_49_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_49_bht_T_20 = _btb_49_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_21 = _btb_49_bht_T_16 ? 2'h0 : _btb_49_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_22 = _btb_49_bht_T_13 ? 2'h0 : _btb_49_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_23 = _btb_49_bht_T_10 ? 2'h0 : _btb_49_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_24 = _btb_49_bht_T_7 ? 2'h3 : _btb_49_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_25 = _btb_49_bht_T_5 ? 2'h3 : _btb_49_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_26 = _btb_49_bht_T_3 ? 2'h3 : _btb_49_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_49_bht_T_27 = _btb_49_bht_T_1 ? 2'h1 : _btb_49_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8902 = btb_49_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6705; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8904 = btb_49_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_49_bht_T_27 : _GEN_8241; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_50_bht_T = btb_50_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_50_bht_T_1 = io_i_branch_resolve_pack_taken & btb_50_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_50_bht_T_2 = btb_50_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_50_bht_T_3 = io_i_branch_resolve_pack_taken & btb_50_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_50_bht_T_4 = btb_50_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_50_bht_T_5 = io_i_branch_resolve_pack_taken & btb_50_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_50_bht_T_6 = btb_50_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_50_bht_T_7 = io_i_branch_resolve_pack_taken & btb_50_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_50_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_50_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_50_bht_T_13 = _btb_0_bht_T_8 & _btb_50_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_50_bht_T_16 = _btb_0_bht_T_8 & _btb_50_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_50_bht_T_19 = _btb_0_bht_T_8 & _btb_50_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_50_bht_T_20 = _btb_50_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_21 = _btb_50_bht_T_16 ? 2'h0 : _btb_50_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_22 = _btb_50_bht_T_13 ? 2'h0 : _btb_50_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_23 = _btb_50_bht_T_10 ? 2'h0 : _btb_50_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_24 = _btb_50_bht_T_7 ? 2'h3 : _btb_50_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_25 = _btb_50_bht_T_5 ? 2'h3 : _btb_50_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_26 = _btb_50_bht_T_3 ? 2'h3 : _btb_50_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_50_bht_T_27 = _btb_50_bht_T_1 ? 2'h1 : _btb_50_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8906 = btb_50_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6706; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8908 = btb_50_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_50_bht_T_27 : _GEN_8242; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_51_bht_T = btb_51_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_51_bht_T_1 = io_i_branch_resolve_pack_taken & btb_51_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_51_bht_T_2 = btb_51_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_51_bht_T_3 = io_i_branch_resolve_pack_taken & btb_51_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_51_bht_T_4 = btb_51_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_51_bht_T_5 = io_i_branch_resolve_pack_taken & btb_51_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_51_bht_T_6 = btb_51_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_51_bht_T_7 = io_i_branch_resolve_pack_taken & btb_51_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_51_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_51_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_51_bht_T_13 = _btb_0_bht_T_8 & _btb_51_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_51_bht_T_16 = _btb_0_bht_T_8 & _btb_51_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_51_bht_T_19 = _btb_0_bht_T_8 & _btb_51_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_51_bht_T_20 = _btb_51_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_21 = _btb_51_bht_T_16 ? 2'h0 : _btb_51_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_22 = _btb_51_bht_T_13 ? 2'h0 : _btb_51_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_23 = _btb_51_bht_T_10 ? 2'h0 : _btb_51_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_24 = _btb_51_bht_T_7 ? 2'h3 : _btb_51_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_25 = _btb_51_bht_T_5 ? 2'h3 : _btb_51_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_26 = _btb_51_bht_T_3 ? 2'h3 : _btb_51_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_51_bht_T_27 = _btb_51_bht_T_1 ? 2'h1 : _btb_51_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8910 = btb_51_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6707; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8912 = btb_51_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_51_bht_T_27 : _GEN_8243; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_52_bht_T = btb_52_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_52_bht_T_1 = io_i_branch_resolve_pack_taken & btb_52_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_52_bht_T_2 = btb_52_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_52_bht_T_3 = io_i_branch_resolve_pack_taken & btb_52_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_52_bht_T_4 = btb_52_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_52_bht_T_5 = io_i_branch_resolve_pack_taken & btb_52_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_52_bht_T_6 = btb_52_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_52_bht_T_7 = io_i_branch_resolve_pack_taken & btb_52_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_52_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_52_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_52_bht_T_13 = _btb_0_bht_T_8 & _btb_52_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_52_bht_T_16 = _btb_0_bht_T_8 & _btb_52_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_52_bht_T_19 = _btb_0_bht_T_8 & _btb_52_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_52_bht_T_20 = _btb_52_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_21 = _btb_52_bht_T_16 ? 2'h0 : _btb_52_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_22 = _btb_52_bht_T_13 ? 2'h0 : _btb_52_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_23 = _btb_52_bht_T_10 ? 2'h0 : _btb_52_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_24 = _btb_52_bht_T_7 ? 2'h3 : _btb_52_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_25 = _btb_52_bht_T_5 ? 2'h3 : _btb_52_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_26 = _btb_52_bht_T_3 ? 2'h3 : _btb_52_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_52_bht_T_27 = _btb_52_bht_T_1 ? 2'h1 : _btb_52_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8914 = btb_52_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6708; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8916 = btb_52_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_52_bht_T_27 : _GEN_8244; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_53_bht_T = btb_53_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_53_bht_T_1 = io_i_branch_resolve_pack_taken & btb_53_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_53_bht_T_2 = btb_53_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_53_bht_T_3 = io_i_branch_resolve_pack_taken & btb_53_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_53_bht_T_4 = btb_53_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_53_bht_T_5 = io_i_branch_resolve_pack_taken & btb_53_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_53_bht_T_6 = btb_53_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_53_bht_T_7 = io_i_branch_resolve_pack_taken & btb_53_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_53_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_53_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_53_bht_T_13 = _btb_0_bht_T_8 & _btb_53_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_53_bht_T_16 = _btb_0_bht_T_8 & _btb_53_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_53_bht_T_19 = _btb_0_bht_T_8 & _btb_53_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_53_bht_T_20 = _btb_53_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_21 = _btb_53_bht_T_16 ? 2'h0 : _btb_53_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_22 = _btb_53_bht_T_13 ? 2'h0 : _btb_53_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_23 = _btb_53_bht_T_10 ? 2'h0 : _btb_53_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_24 = _btb_53_bht_T_7 ? 2'h3 : _btb_53_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_25 = _btb_53_bht_T_5 ? 2'h3 : _btb_53_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_26 = _btb_53_bht_T_3 ? 2'h3 : _btb_53_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_53_bht_T_27 = _btb_53_bht_T_1 ? 2'h1 : _btb_53_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8918 = btb_53_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6709; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8920 = btb_53_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_53_bht_T_27 : _GEN_8245; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_54_bht_T = btb_54_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_54_bht_T_1 = io_i_branch_resolve_pack_taken & btb_54_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_54_bht_T_2 = btb_54_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_54_bht_T_3 = io_i_branch_resolve_pack_taken & btb_54_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_54_bht_T_4 = btb_54_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_54_bht_T_5 = io_i_branch_resolve_pack_taken & btb_54_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_54_bht_T_6 = btb_54_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_54_bht_T_7 = io_i_branch_resolve_pack_taken & btb_54_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_54_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_54_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_54_bht_T_13 = _btb_0_bht_T_8 & _btb_54_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_54_bht_T_16 = _btb_0_bht_T_8 & _btb_54_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_54_bht_T_19 = _btb_0_bht_T_8 & _btb_54_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_54_bht_T_20 = _btb_54_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_21 = _btb_54_bht_T_16 ? 2'h0 : _btb_54_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_22 = _btb_54_bht_T_13 ? 2'h0 : _btb_54_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_23 = _btb_54_bht_T_10 ? 2'h0 : _btb_54_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_24 = _btb_54_bht_T_7 ? 2'h3 : _btb_54_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_25 = _btb_54_bht_T_5 ? 2'h3 : _btb_54_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_26 = _btb_54_bht_T_3 ? 2'h3 : _btb_54_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_54_bht_T_27 = _btb_54_bht_T_1 ? 2'h1 : _btb_54_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8922 = btb_54_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6710; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8924 = btb_54_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_54_bht_T_27 : _GEN_8246; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_55_bht_T = btb_55_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_55_bht_T_1 = io_i_branch_resolve_pack_taken & btb_55_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_55_bht_T_2 = btb_55_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_55_bht_T_3 = io_i_branch_resolve_pack_taken & btb_55_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_55_bht_T_4 = btb_55_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_55_bht_T_5 = io_i_branch_resolve_pack_taken & btb_55_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_55_bht_T_6 = btb_55_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_55_bht_T_7 = io_i_branch_resolve_pack_taken & btb_55_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_55_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_55_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_55_bht_T_13 = _btb_0_bht_T_8 & _btb_55_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_55_bht_T_16 = _btb_0_bht_T_8 & _btb_55_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_55_bht_T_19 = _btb_0_bht_T_8 & _btb_55_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_55_bht_T_20 = _btb_55_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_21 = _btb_55_bht_T_16 ? 2'h0 : _btb_55_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_22 = _btb_55_bht_T_13 ? 2'h0 : _btb_55_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_23 = _btb_55_bht_T_10 ? 2'h0 : _btb_55_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_24 = _btb_55_bht_T_7 ? 2'h3 : _btb_55_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_25 = _btb_55_bht_T_5 ? 2'h3 : _btb_55_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_26 = _btb_55_bht_T_3 ? 2'h3 : _btb_55_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_55_bht_T_27 = _btb_55_bht_T_1 ? 2'h1 : _btb_55_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8926 = btb_55_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6711; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8928 = btb_55_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_55_bht_T_27 : _GEN_8247; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_56_bht_T = btb_56_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_56_bht_T_1 = io_i_branch_resolve_pack_taken & btb_56_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_56_bht_T_2 = btb_56_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_56_bht_T_3 = io_i_branch_resolve_pack_taken & btb_56_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_56_bht_T_4 = btb_56_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_56_bht_T_5 = io_i_branch_resolve_pack_taken & btb_56_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_56_bht_T_6 = btb_56_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_56_bht_T_7 = io_i_branch_resolve_pack_taken & btb_56_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_56_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_56_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_56_bht_T_13 = _btb_0_bht_T_8 & _btb_56_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_56_bht_T_16 = _btb_0_bht_T_8 & _btb_56_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_56_bht_T_19 = _btb_0_bht_T_8 & _btb_56_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_56_bht_T_20 = _btb_56_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_21 = _btb_56_bht_T_16 ? 2'h0 : _btb_56_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_22 = _btb_56_bht_T_13 ? 2'h0 : _btb_56_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_23 = _btb_56_bht_T_10 ? 2'h0 : _btb_56_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_24 = _btb_56_bht_T_7 ? 2'h3 : _btb_56_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_25 = _btb_56_bht_T_5 ? 2'h3 : _btb_56_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_26 = _btb_56_bht_T_3 ? 2'h3 : _btb_56_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_56_bht_T_27 = _btb_56_bht_T_1 ? 2'h1 : _btb_56_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8930 = btb_56_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6712; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8932 = btb_56_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_56_bht_T_27 : _GEN_8248; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_57_bht_T = btb_57_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_57_bht_T_1 = io_i_branch_resolve_pack_taken & btb_57_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_57_bht_T_2 = btb_57_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_57_bht_T_3 = io_i_branch_resolve_pack_taken & btb_57_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_57_bht_T_4 = btb_57_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_57_bht_T_5 = io_i_branch_resolve_pack_taken & btb_57_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_57_bht_T_6 = btb_57_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_57_bht_T_7 = io_i_branch_resolve_pack_taken & btb_57_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_57_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_57_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_57_bht_T_13 = _btb_0_bht_T_8 & _btb_57_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_57_bht_T_16 = _btb_0_bht_T_8 & _btb_57_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_57_bht_T_19 = _btb_0_bht_T_8 & _btb_57_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_57_bht_T_20 = _btb_57_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_21 = _btb_57_bht_T_16 ? 2'h0 : _btb_57_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_22 = _btb_57_bht_T_13 ? 2'h0 : _btb_57_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_23 = _btb_57_bht_T_10 ? 2'h0 : _btb_57_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_24 = _btb_57_bht_T_7 ? 2'h3 : _btb_57_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_25 = _btb_57_bht_T_5 ? 2'h3 : _btb_57_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_26 = _btb_57_bht_T_3 ? 2'h3 : _btb_57_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_57_bht_T_27 = _btb_57_bht_T_1 ? 2'h1 : _btb_57_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8934 = btb_57_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6713; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8936 = btb_57_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_57_bht_T_27 : _GEN_8249; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_58_bht_T = btb_58_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_58_bht_T_1 = io_i_branch_resolve_pack_taken & btb_58_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_58_bht_T_2 = btb_58_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_58_bht_T_3 = io_i_branch_resolve_pack_taken & btb_58_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_58_bht_T_4 = btb_58_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_58_bht_T_5 = io_i_branch_resolve_pack_taken & btb_58_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_58_bht_T_6 = btb_58_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_58_bht_T_7 = io_i_branch_resolve_pack_taken & btb_58_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_58_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_58_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_58_bht_T_13 = _btb_0_bht_T_8 & _btb_58_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_58_bht_T_16 = _btb_0_bht_T_8 & _btb_58_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_58_bht_T_19 = _btb_0_bht_T_8 & _btb_58_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_58_bht_T_20 = _btb_58_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_21 = _btb_58_bht_T_16 ? 2'h0 : _btb_58_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_22 = _btb_58_bht_T_13 ? 2'h0 : _btb_58_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_23 = _btb_58_bht_T_10 ? 2'h0 : _btb_58_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_24 = _btb_58_bht_T_7 ? 2'h3 : _btb_58_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_25 = _btb_58_bht_T_5 ? 2'h3 : _btb_58_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_26 = _btb_58_bht_T_3 ? 2'h3 : _btb_58_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_58_bht_T_27 = _btb_58_bht_T_1 ? 2'h1 : _btb_58_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8938 = btb_58_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6714; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8940 = btb_58_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_58_bht_T_27 : _GEN_8250; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_59_bht_T = btb_59_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_59_bht_T_1 = io_i_branch_resolve_pack_taken & btb_59_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_59_bht_T_2 = btb_59_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_59_bht_T_3 = io_i_branch_resolve_pack_taken & btb_59_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_59_bht_T_4 = btb_59_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_59_bht_T_5 = io_i_branch_resolve_pack_taken & btb_59_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_59_bht_T_6 = btb_59_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_59_bht_T_7 = io_i_branch_resolve_pack_taken & btb_59_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_59_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_59_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_59_bht_T_13 = _btb_0_bht_T_8 & _btb_59_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_59_bht_T_16 = _btb_0_bht_T_8 & _btb_59_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_59_bht_T_19 = _btb_0_bht_T_8 & _btb_59_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_59_bht_T_20 = _btb_59_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_21 = _btb_59_bht_T_16 ? 2'h0 : _btb_59_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_22 = _btb_59_bht_T_13 ? 2'h0 : _btb_59_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_23 = _btb_59_bht_T_10 ? 2'h0 : _btb_59_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_24 = _btb_59_bht_T_7 ? 2'h3 : _btb_59_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_25 = _btb_59_bht_T_5 ? 2'h3 : _btb_59_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_26 = _btb_59_bht_T_3 ? 2'h3 : _btb_59_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_59_bht_T_27 = _btb_59_bht_T_1 ? 2'h1 : _btb_59_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_8941 = btb_59_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_58_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_57_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_56_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_55_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_54_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_53_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_52_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_51_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_50_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_49_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_48_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_47_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_46_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_45_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_8881)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_8942 = btb_59_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6715; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8944 = btb_59_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_59_bht_T_27 : _GEN_8251; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_60_bht_T = btb_60_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_60_bht_T_1 = io_i_branch_resolve_pack_taken & btb_60_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_60_bht_T_2 = btb_60_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_60_bht_T_3 = io_i_branch_resolve_pack_taken & btb_60_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_60_bht_T_4 = btb_60_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_60_bht_T_5 = io_i_branch_resolve_pack_taken & btb_60_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_60_bht_T_6 = btb_60_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_60_bht_T_7 = io_i_branch_resolve_pack_taken & btb_60_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_60_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_60_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_60_bht_T_13 = _btb_0_bht_T_8 & _btb_60_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_60_bht_T_16 = _btb_0_bht_T_8 & _btb_60_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_60_bht_T_19 = _btb_0_bht_T_8 & _btb_60_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_60_bht_T_20 = _btb_60_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_21 = _btb_60_bht_T_16 ? 2'h0 : _btb_60_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_22 = _btb_60_bht_T_13 ? 2'h0 : _btb_60_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_23 = _btb_60_bht_T_10 ? 2'h0 : _btb_60_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_24 = _btb_60_bht_T_7 ? 2'h3 : _btb_60_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_25 = _btb_60_bht_T_5 ? 2'h3 : _btb_60_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_26 = _btb_60_bht_T_3 ? 2'h3 : _btb_60_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_60_bht_T_27 = _btb_60_bht_T_1 ? 2'h1 : _btb_60_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8946 = btb_60_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6716; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8948 = btb_60_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_60_bht_T_27 : _GEN_8252; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_61_bht_T = btb_61_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_61_bht_T_1 = io_i_branch_resolve_pack_taken & btb_61_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_61_bht_T_2 = btb_61_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_61_bht_T_3 = io_i_branch_resolve_pack_taken & btb_61_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_61_bht_T_4 = btb_61_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_61_bht_T_5 = io_i_branch_resolve_pack_taken & btb_61_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_61_bht_T_6 = btb_61_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_61_bht_T_7 = io_i_branch_resolve_pack_taken & btb_61_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_61_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_61_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_61_bht_T_13 = _btb_0_bht_T_8 & _btb_61_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_61_bht_T_16 = _btb_0_bht_T_8 & _btb_61_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_61_bht_T_19 = _btb_0_bht_T_8 & _btb_61_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_61_bht_T_20 = _btb_61_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_21 = _btb_61_bht_T_16 ? 2'h0 : _btb_61_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_22 = _btb_61_bht_T_13 ? 2'h0 : _btb_61_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_23 = _btb_61_bht_T_10 ? 2'h0 : _btb_61_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_24 = _btb_61_bht_T_7 ? 2'h3 : _btb_61_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_25 = _btb_61_bht_T_5 ? 2'h3 : _btb_61_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_26 = _btb_61_bht_T_3 ? 2'h3 : _btb_61_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_61_bht_T_27 = _btb_61_bht_T_1 ? 2'h1 : _btb_61_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8950 = btb_61_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6717; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8952 = btb_61_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_61_bht_T_27 : _GEN_8253; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_62_bht_T = btb_62_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_62_bht_T_1 = io_i_branch_resolve_pack_taken & btb_62_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_62_bht_T_2 = btb_62_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_62_bht_T_3 = io_i_branch_resolve_pack_taken & btb_62_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_62_bht_T_4 = btb_62_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_62_bht_T_5 = io_i_branch_resolve_pack_taken & btb_62_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_62_bht_T_6 = btb_62_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_62_bht_T_7 = io_i_branch_resolve_pack_taken & btb_62_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_62_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_62_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_62_bht_T_13 = _btb_0_bht_T_8 & _btb_62_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_62_bht_T_16 = _btb_0_bht_T_8 & _btb_62_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_62_bht_T_19 = _btb_0_bht_T_8 & _btb_62_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_62_bht_T_20 = _btb_62_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_21 = _btb_62_bht_T_16 ? 2'h0 : _btb_62_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_22 = _btb_62_bht_T_13 ? 2'h0 : _btb_62_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_23 = _btb_62_bht_T_10 ? 2'h0 : _btb_62_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_24 = _btb_62_bht_T_7 ? 2'h3 : _btb_62_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_25 = _btb_62_bht_T_5 ? 2'h3 : _btb_62_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_26 = _btb_62_bht_T_3 ? 2'h3 : _btb_62_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_62_bht_T_27 = _btb_62_bht_T_1 ? 2'h1 : _btb_62_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8954 = btb_62_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6718; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8956 = btb_62_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_62_bht_T_27 : _GEN_8254; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_63_bht_T = btb_63_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_63_bht_T_1 = io_i_branch_resolve_pack_taken & btb_63_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_63_bht_T_2 = btb_63_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_63_bht_T_3 = io_i_branch_resolve_pack_taken & btb_63_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_63_bht_T_4 = btb_63_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_63_bht_T_5 = io_i_branch_resolve_pack_taken & btb_63_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_63_bht_T_6 = btb_63_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_63_bht_T_7 = io_i_branch_resolve_pack_taken & btb_63_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_63_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_63_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_63_bht_T_13 = _btb_0_bht_T_8 & _btb_63_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_63_bht_T_16 = _btb_0_bht_T_8 & _btb_63_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_63_bht_T_19 = _btb_0_bht_T_8 & _btb_63_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_63_bht_T_20 = _btb_63_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_21 = _btb_63_bht_T_16 ? 2'h0 : _btb_63_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_22 = _btb_63_bht_T_13 ? 2'h0 : _btb_63_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_23 = _btb_63_bht_T_10 ? 2'h0 : _btb_63_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_24 = _btb_63_bht_T_7 ? 2'h3 : _btb_63_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_25 = _btb_63_bht_T_5 ? 2'h3 : _btb_63_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_26 = _btb_63_bht_T_3 ? 2'h3 : _btb_63_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_63_bht_T_27 = _btb_63_bht_T_1 ? 2'h1 : _btb_63_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8958 = btb_63_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6719; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8960 = btb_63_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_63_bht_T_27 : _GEN_8255; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_64_bht_T = btb_64_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_64_bht_T_1 = io_i_branch_resolve_pack_taken & btb_64_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_64_bht_T_2 = btb_64_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_64_bht_T_3 = io_i_branch_resolve_pack_taken & btb_64_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_64_bht_T_4 = btb_64_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_64_bht_T_5 = io_i_branch_resolve_pack_taken & btb_64_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_64_bht_T_6 = btb_64_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_64_bht_T_7 = io_i_branch_resolve_pack_taken & btb_64_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_64_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_64_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_64_bht_T_13 = _btb_0_bht_T_8 & _btb_64_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_64_bht_T_16 = _btb_0_bht_T_8 & _btb_64_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_64_bht_T_19 = _btb_0_bht_T_8 & _btb_64_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_64_bht_T_20 = _btb_64_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_21 = _btb_64_bht_T_16 ? 2'h0 : _btb_64_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_22 = _btb_64_bht_T_13 ? 2'h0 : _btb_64_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_23 = _btb_64_bht_T_10 ? 2'h0 : _btb_64_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_24 = _btb_64_bht_T_7 ? 2'h3 : _btb_64_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_25 = _btb_64_bht_T_5 ? 2'h3 : _btb_64_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_26 = _btb_64_bht_T_3 ? 2'h3 : _btb_64_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_64_bht_T_27 = _btb_64_bht_T_1 ? 2'h1 : _btb_64_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8962 = btb_64_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6720; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8964 = btb_64_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_64_bht_T_27 : _GEN_8256; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_65_bht_T = btb_65_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_65_bht_T_1 = io_i_branch_resolve_pack_taken & btb_65_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_65_bht_T_2 = btb_65_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_65_bht_T_3 = io_i_branch_resolve_pack_taken & btb_65_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_65_bht_T_4 = btb_65_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_65_bht_T_5 = io_i_branch_resolve_pack_taken & btb_65_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_65_bht_T_6 = btb_65_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_65_bht_T_7 = io_i_branch_resolve_pack_taken & btb_65_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_65_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_65_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_65_bht_T_13 = _btb_0_bht_T_8 & _btb_65_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_65_bht_T_16 = _btb_0_bht_T_8 & _btb_65_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_65_bht_T_19 = _btb_0_bht_T_8 & _btb_65_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_65_bht_T_20 = _btb_65_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_21 = _btb_65_bht_T_16 ? 2'h0 : _btb_65_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_22 = _btb_65_bht_T_13 ? 2'h0 : _btb_65_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_23 = _btb_65_bht_T_10 ? 2'h0 : _btb_65_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_24 = _btb_65_bht_T_7 ? 2'h3 : _btb_65_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_25 = _btb_65_bht_T_5 ? 2'h3 : _btb_65_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_26 = _btb_65_bht_T_3 ? 2'h3 : _btb_65_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_65_bht_T_27 = _btb_65_bht_T_1 ? 2'h1 : _btb_65_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8966 = btb_65_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6721; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8968 = btb_65_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_65_bht_T_27 : _GEN_8257; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_66_bht_T = btb_66_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_66_bht_T_1 = io_i_branch_resolve_pack_taken & btb_66_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_66_bht_T_2 = btb_66_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_66_bht_T_3 = io_i_branch_resolve_pack_taken & btb_66_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_66_bht_T_4 = btb_66_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_66_bht_T_5 = io_i_branch_resolve_pack_taken & btb_66_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_66_bht_T_6 = btb_66_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_66_bht_T_7 = io_i_branch_resolve_pack_taken & btb_66_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_66_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_66_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_66_bht_T_13 = _btb_0_bht_T_8 & _btb_66_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_66_bht_T_16 = _btb_0_bht_T_8 & _btb_66_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_66_bht_T_19 = _btb_0_bht_T_8 & _btb_66_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_66_bht_T_20 = _btb_66_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_21 = _btb_66_bht_T_16 ? 2'h0 : _btb_66_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_22 = _btb_66_bht_T_13 ? 2'h0 : _btb_66_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_23 = _btb_66_bht_T_10 ? 2'h0 : _btb_66_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_24 = _btb_66_bht_T_7 ? 2'h3 : _btb_66_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_25 = _btb_66_bht_T_5 ? 2'h3 : _btb_66_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_26 = _btb_66_bht_T_3 ? 2'h3 : _btb_66_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_66_bht_T_27 = _btb_66_bht_T_1 ? 2'h1 : _btb_66_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8970 = btb_66_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6722; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8972 = btb_66_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_66_bht_T_27 : _GEN_8258; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_67_bht_T = btb_67_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_67_bht_T_1 = io_i_branch_resolve_pack_taken & btb_67_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_67_bht_T_2 = btb_67_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_67_bht_T_3 = io_i_branch_resolve_pack_taken & btb_67_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_67_bht_T_4 = btb_67_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_67_bht_T_5 = io_i_branch_resolve_pack_taken & btb_67_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_67_bht_T_6 = btb_67_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_67_bht_T_7 = io_i_branch_resolve_pack_taken & btb_67_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_67_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_67_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_67_bht_T_13 = _btb_0_bht_T_8 & _btb_67_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_67_bht_T_16 = _btb_0_bht_T_8 & _btb_67_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_67_bht_T_19 = _btb_0_bht_T_8 & _btb_67_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_67_bht_T_20 = _btb_67_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_21 = _btb_67_bht_T_16 ? 2'h0 : _btb_67_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_22 = _btb_67_bht_T_13 ? 2'h0 : _btb_67_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_23 = _btb_67_bht_T_10 ? 2'h0 : _btb_67_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_24 = _btb_67_bht_T_7 ? 2'h3 : _btb_67_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_25 = _btb_67_bht_T_5 ? 2'h3 : _btb_67_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_26 = _btb_67_bht_T_3 ? 2'h3 : _btb_67_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_67_bht_T_27 = _btb_67_bht_T_1 ? 2'h1 : _btb_67_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8974 = btb_67_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6723; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8976 = btb_67_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_67_bht_T_27 : _GEN_8259; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_68_bht_T = btb_68_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_68_bht_T_1 = io_i_branch_resolve_pack_taken & btb_68_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_68_bht_T_2 = btb_68_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_68_bht_T_3 = io_i_branch_resolve_pack_taken & btb_68_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_68_bht_T_4 = btb_68_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_68_bht_T_5 = io_i_branch_resolve_pack_taken & btb_68_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_68_bht_T_6 = btb_68_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_68_bht_T_7 = io_i_branch_resolve_pack_taken & btb_68_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_68_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_68_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_68_bht_T_13 = _btb_0_bht_T_8 & _btb_68_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_68_bht_T_16 = _btb_0_bht_T_8 & _btb_68_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_68_bht_T_19 = _btb_0_bht_T_8 & _btb_68_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_68_bht_T_20 = _btb_68_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_21 = _btb_68_bht_T_16 ? 2'h0 : _btb_68_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_22 = _btb_68_bht_T_13 ? 2'h0 : _btb_68_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_23 = _btb_68_bht_T_10 ? 2'h0 : _btb_68_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_24 = _btb_68_bht_T_7 ? 2'h3 : _btb_68_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_25 = _btb_68_bht_T_5 ? 2'h3 : _btb_68_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_26 = _btb_68_bht_T_3 ? 2'h3 : _btb_68_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_68_bht_T_27 = _btb_68_bht_T_1 ? 2'h1 : _btb_68_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8978 = btb_68_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6724; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8980 = btb_68_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_68_bht_T_27 : _GEN_8260; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_69_bht_T = btb_69_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_69_bht_T_1 = io_i_branch_resolve_pack_taken & btb_69_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_69_bht_T_2 = btb_69_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_69_bht_T_3 = io_i_branch_resolve_pack_taken & btb_69_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_69_bht_T_4 = btb_69_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_69_bht_T_5 = io_i_branch_resolve_pack_taken & btb_69_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_69_bht_T_6 = btb_69_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_69_bht_T_7 = io_i_branch_resolve_pack_taken & btb_69_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_69_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_69_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_69_bht_T_13 = _btb_0_bht_T_8 & _btb_69_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_69_bht_T_16 = _btb_0_bht_T_8 & _btb_69_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_69_bht_T_19 = _btb_0_bht_T_8 & _btb_69_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_69_bht_T_20 = _btb_69_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_21 = _btb_69_bht_T_16 ? 2'h0 : _btb_69_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_22 = _btb_69_bht_T_13 ? 2'h0 : _btb_69_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_23 = _btb_69_bht_T_10 ? 2'h0 : _btb_69_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_24 = _btb_69_bht_T_7 ? 2'h3 : _btb_69_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_25 = _btb_69_bht_T_5 ? 2'h3 : _btb_69_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_26 = _btb_69_bht_T_3 ? 2'h3 : _btb_69_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_69_bht_T_27 = _btb_69_bht_T_1 ? 2'h1 : _btb_69_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8982 = btb_69_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6725; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8984 = btb_69_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_69_bht_T_27 : _GEN_8261; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_70_bht_T = btb_70_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_70_bht_T_1 = io_i_branch_resolve_pack_taken & btb_70_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_70_bht_T_2 = btb_70_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_70_bht_T_3 = io_i_branch_resolve_pack_taken & btb_70_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_70_bht_T_4 = btb_70_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_70_bht_T_5 = io_i_branch_resolve_pack_taken & btb_70_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_70_bht_T_6 = btb_70_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_70_bht_T_7 = io_i_branch_resolve_pack_taken & btb_70_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_70_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_70_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_70_bht_T_13 = _btb_0_bht_T_8 & _btb_70_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_70_bht_T_16 = _btb_0_bht_T_8 & _btb_70_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_70_bht_T_19 = _btb_0_bht_T_8 & _btb_70_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_70_bht_T_20 = _btb_70_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_21 = _btb_70_bht_T_16 ? 2'h0 : _btb_70_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_22 = _btb_70_bht_T_13 ? 2'h0 : _btb_70_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_23 = _btb_70_bht_T_10 ? 2'h0 : _btb_70_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_24 = _btb_70_bht_T_7 ? 2'h3 : _btb_70_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_25 = _btb_70_bht_T_5 ? 2'h3 : _btb_70_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_26 = _btb_70_bht_T_3 ? 2'h3 : _btb_70_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_70_bht_T_27 = _btb_70_bht_T_1 ? 2'h1 : _btb_70_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8986 = btb_70_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6726; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8988 = btb_70_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_70_bht_T_27 : _GEN_8262; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_71_bht_T = btb_71_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_71_bht_T_1 = io_i_branch_resolve_pack_taken & btb_71_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_71_bht_T_2 = btb_71_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_71_bht_T_3 = io_i_branch_resolve_pack_taken & btb_71_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_71_bht_T_4 = btb_71_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_71_bht_T_5 = io_i_branch_resolve_pack_taken & btb_71_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_71_bht_T_6 = btb_71_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_71_bht_T_7 = io_i_branch_resolve_pack_taken & btb_71_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_71_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_71_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_71_bht_T_13 = _btb_0_bht_T_8 & _btb_71_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_71_bht_T_16 = _btb_0_bht_T_8 & _btb_71_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_71_bht_T_19 = _btb_0_bht_T_8 & _btb_71_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_71_bht_T_20 = _btb_71_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_21 = _btb_71_bht_T_16 ? 2'h0 : _btb_71_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_22 = _btb_71_bht_T_13 ? 2'h0 : _btb_71_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_23 = _btb_71_bht_T_10 ? 2'h0 : _btb_71_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_24 = _btb_71_bht_T_7 ? 2'h3 : _btb_71_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_25 = _btb_71_bht_T_5 ? 2'h3 : _btb_71_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_26 = _btb_71_bht_T_3 ? 2'h3 : _btb_71_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_71_bht_T_27 = _btb_71_bht_T_1 ? 2'h1 : _btb_71_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8990 = btb_71_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6727; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8992 = btb_71_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_71_bht_T_27 : _GEN_8263; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_72_bht_T = btb_72_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_72_bht_T_1 = io_i_branch_resolve_pack_taken & btb_72_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_72_bht_T_2 = btb_72_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_72_bht_T_3 = io_i_branch_resolve_pack_taken & btb_72_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_72_bht_T_4 = btb_72_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_72_bht_T_5 = io_i_branch_resolve_pack_taken & btb_72_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_72_bht_T_6 = btb_72_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_72_bht_T_7 = io_i_branch_resolve_pack_taken & btb_72_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_72_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_72_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_72_bht_T_13 = _btb_0_bht_T_8 & _btb_72_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_72_bht_T_16 = _btb_0_bht_T_8 & _btb_72_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_72_bht_T_19 = _btb_0_bht_T_8 & _btb_72_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_72_bht_T_20 = _btb_72_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_21 = _btb_72_bht_T_16 ? 2'h0 : _btb_72_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_22 = _btb_72_bht_T_13 ? 2'h0 : _btb_72_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_23 = _btb_72_bht_T_10 ? 2'h0 : _btb_72_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_24 = _btb_72_bht_T_7 ? 2'h3 : _btb_72_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_25 = _btb_72_bht_T_5 ? 2'h3 : _btb_72_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_26 = _btb_72_bht_T_3 ? 2'h3 : _btb_72_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_72_bht_T_27 = _btb_72_bht_T_1 ? 2'h1 : _btb_72_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8994 = btb_72_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6728; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_8996 = btb_72_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_72_bht_T_27 : _GEN_8264; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_73_bht_T = btb_73_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_73_bht_T_1 = io_i_branch_resolve_pack_taken & btb_73_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_73_bht_T_2 = btb_73_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_73_bht_T_3 = io_i_branch_resolve_pack_taken & btb_73_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_73_bht_T_4 = btb_73_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_73_bht_T_5 = io_i_branch_resolve_pack_taken & btb_73_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_73_bht_T_6 = btb_73_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_73_bht_T_7 = io_i_branch_resolve_pack_taken & btb_73_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_73_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_73_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_73_bht_T_13 = _btb_0_bht_T_8 & _btb_73_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_73_bht_T_16 = _btb_0_bht_T_8 & _btb_73_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_73_bht_T_19 = _btb_0_bht_T_8 & _btb_73_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_73_bht_T_20 = _btb_73_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_21 = _btb_73_bht_T_16 ? 2'h0 : _btb_73_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_22 = _btb_73_bht_T_13 ? 2'h0 : _btb_73_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_23 = _btb_73_bht_T_10 ? 2'h0 : _btb_73_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_24 = _btb_73_bht_T_7 ? 2'h3 : _btb_73_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_25 = _btb_73_bht_T_5 ? 2'h3 : _btb_73_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_26 = _btb_73_bht_T_3 ? 2'h3 : _btb_73_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_73_bht_T_27 = _btb_73_bht_T_1 ? 2'h1 : _btb_73_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_8998 = btb_73_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6729; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9000 = btb_73_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_73_bht_T_27 : _GEN_8265; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_74_bht_T = btb_74_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_74_bht_T_1 = io_i_branch_resolve_pack_taken & btb_74_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_74_bht_T_2 = btb_74_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_74_bht_T_3 = io_i_branch_resolve_pack_taken & btb_74_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_74_bht_T_4 = btb_74_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_74_bht_T_5 = io_i_branch_resolve_pack_taken & btb_74_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_74_bht_T_6 = btb_74_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_74_bht_T_7 = io_i_branch_resolve_pack_taken & btb_74_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_74_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_74_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_74_bht_T_13 = _btb_0_bht_T_8 & _btb_74_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_74_bht_T_16 = _btb_0_bht_T_8 & _btb_74_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_74_bht_T_19 = _btb_0_bht_T_8 & _btb_74_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_74_bht_T_20 = _btb_74_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_21 = _btb_74_bht_T_16 ? 2'h0 : _btb_74_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_22 = _btb_74_bht_T_13 ? 2'h0 : _btb_74_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_23 = _btb_74_bht_T_10 ? 2'h0 : _btb_74_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_24 = _btb_74_bht_T_7 ? 2'h3 : _btb_74_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_25 = _btb_74_bht_T_5 ? 2'h3 : _btb_74_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_26 = _btb_74_bht_T_3 ? 2'h3 : _btb_74_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_74_bht_T_27 = _btb_74_bht_T_1 ? 2'h1 : _btb_74_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9001 = btb_74_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_73_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_72_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_71_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_70_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_69_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_68_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_67_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_66_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_65_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_64_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_63_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_62_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_61_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_60_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_8941)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9002 = btb_74_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6730; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9004 = btb_74_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_74_bht_T_27 : _GEN_8266; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_75_bht_T = btb_75_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_75_bht_T_1 = io_i_branch_resolve_pack_taken & btb_75_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_75_bht_T_2 = btb_75_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_75_bht_T_3 = io_i_branch_resolve_pack_taken & btb_75_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_75_bht_T_4 = btb_75_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_75_bht_T_5 = io_i_branch_resolve_pack_taken & btb_75_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_75_bht_T_6 = btb_75_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_75_bht_T_7 = io_i_branch_resolve_pack_taken & btb_75_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_75_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_75_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_75_bht_T_13 = _btb_0_bht_T_8 & _btb_75_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_75_bht_T_16 = _btb_0_bht_T_8 & _btb_75_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_75_bht_T_19 = _btb_0_bht_T_8 & _btb_75_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_75_bht_T_20 = _btb_75_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_21 = _btb_75_bht_T_16 ? 2'h0 : _btb_75_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_22 = _btb_75_bht_T_13 ? 2'h0 : _btb_75_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_23 = _btb_75_bht_T_10 ? 2'h0 : _btb_75_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_24 = _btb_75_bht_T_7 ? 2'h3 : _btb_75_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_25 = _btb_75_bht_T_5 ? 2'h3 : _btb_75_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_26 = _btb_75_bht_T_3 ? 2'h3 : _btb_75_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_75_bht_T_27 = _btb_75_bht_T_1 ? 2'h1 : _btb_75_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9006 = btb_75_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6731; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9008 = btb_75_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_75_bht_T_27 : _GEN_8267; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_76_bht_T = btb_76_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_76_bht_T_1 = io_i_branch_resolve_pack_taken & btb_76_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_76_bht_T_2 = btb_76_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_76_bht_T_3 = io_i_branch_resolve_pack_taken & btb_76_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_76_bht_T_4 = btb_76_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_76_bht_T_5 = io_i_branch_resolve_pack_taken & btb_76_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_76_bht_T_6 = btb_76_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_76_bht_T_7 = io_i_branch_resolve_pack_taken & btb_76_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_76_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_76_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_76_bht_T_13 = _btb_0_bht_T_8 & _btb_76_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_76_bht_T_16 = _btb_0_bht_T_8 & _btb_76_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_76_bht_T_19 = _btb_0_bht_T_8 & _btb_76_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_76_bht_T_20 = _btb_76_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_21 = _btb_76_bht_T_16 ? 2'h0 : _btb_76_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_22 = _btb_76_bht_T_13 ? 2'h0 : _btb_76_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_23 = _btb_76_bht_T_10 ? 2'h0 : _btb_76_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_24 = _btb_76_bht_T_7 ? 2'h3 : _btb_76_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_25 = _btb_76_bht_T_5 ? 2'h3 : _btb_76_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_26 = _btb_76_bht_T_3 ? 2'h3 : _btb_76_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_76_bht_T_27 = _btb_76_bht_T_1 ? 2'h1 : _btb_76_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9010 = btb_76_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6732; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9012 = btb_76_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_76_bht_T_27 : _GEN_8268; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_77_bht_T = btb_77_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_77_bht_T_1 = io_i_branch_resolve_pack_taken & btb_77_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_77_bht_T_2 = btb_77_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_77_bht_T_3 = io_i_branch_resolve_pack_taken & btb_77_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_77_bht_T_4 = btb_77_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_77_bht_T_5 = io_i_branch_resolve_pack_taken & btb_77_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_77_bht_T_6 = btb_77_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_77_bht_T_7 = io_i_branch_resolve_pack_taken & btb_77_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_77_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_77_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_77_bht_T_13 = _btb_0_bht_T_8 & _btb_77_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_77_bht_T_16 = _btb_0_bht_T_8 & _btb_77_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_77_bht_T_19 = _btb_0_bht_T_8 & _btb_77_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_77_bht_T_20 = _btb_77_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_21 = _btb_77_bht_T_16 ? 2'h0 : _btb_77_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_22 = _btb_77_bht_T_13 ? 2'h0 : _btb_77_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_23 = _btb_77_bht_T_10 ? 2'h0 : _btb_77_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_24 = _btb_77_bht_T_7 ? 2'h3 : _btb_77_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_25 = _btb_77_bht_T_5 ? 2'h3 : _btb_77_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_26 = _btb_77_bht_T_3 ? 2'h3 : _btb_77_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_77_bht_T_27 = _btb_77_bht_T_1 ? 2'h1 : _btb_77_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9014 = btb_77_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6733; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9016 = btb_77_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_77_bht_T_27 : _GEN_8269; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_78_bht_T = btb_78_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_78_bht_T_1 = io_i_branch_resolve_pack_taken & btb_78_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_78_bht_T_2 = btb_78_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_78_bht_T_3 = io_i_branch_resolve_pack_taken & btb_78_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_78_bht_T_4 = btb_78_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_78_bht_T_5 = io_i_branch_resolve_pack_taken & btb_78_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_78_bht_T_6 = btb_78_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_78_bht_T_7 = io_i_branch_resolve_pack_taken & btb_78_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_78_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_78_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_78_bht_T_13 = _btb_0_bht_T_8 & _btb_78_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_78_bht_T_16 = _btb_0_bht_T_8 & _btb_78_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_78_bht_T_19 = _btb_0_bht_T_8 & _btb_78_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_78_bht_T_20 = _btb_78_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_21 = _btb_78_bht_T_16 ? 2'h0 : _btb_78_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_22 = _btb_78_bht_T_13 ? 2'h0 : _btb_78_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_23 = _btb_78_bht_T_10 ? 2'h0 : _btb_78_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_24 = _btb_78_bht_T_7 ? 2'h3 : _btb_78_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_25 = _btb_78_bht_T_5 ? 2'h3 : _btb_78_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_26 = _btb_78_bht_T_3 ? 2'h3 : _btb_78_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_78_bht_T_27 = _btb_78_bht_T_1 ? 2'h1 : _btb_78_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9018 = btb_78_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6734; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9020 = btb_78_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_78_bht_T_27 : _GEN_8270; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_79_bht_T = btb_79_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_79_bht_T_1 = io_i_branch_resolve_pack_taken & btb_79_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_79_bht_T_2 = btb_79_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_79_bht_T_3 = io_i_branch_resolve_pack_taken & btb_79_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_79_bht_T_4 = btb_79_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_79_bht_T_5 = io_i_branch_resolve_pack_taken & btb_79_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_79_bht_T_6 = btb_79_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_79_bht_T_7 = io_i_branch_resolve_pack_taken & btb_79_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_79_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_79_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_79_bht_T_13 = _btb_0_bht_T_8 & _btb_79_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_79_bht_T_16 = _btb_0_bht_T_8 & _btb_79_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_79_bht_T_19 = _btb_0_bht_T_8 & _btb_79_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_79_bht_T_20 = _btb_79_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_21 = _btb_79_bht_T_16 ? 2'h0 : _btb_79_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_22 = _btb_79_bht_T_13 ? 2'h0 : _btb_79_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_23 = _btb_79_bht_T_10 ? 2'h0 : _btb_79_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_24 = _btb_79_bht_T_7 ? 2'h3 : _btb_79_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_25 = _btb_79_bht_T_5 ? 2'h3 : _btb_79_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_26 = _btb_79_bht_T_3 ? 2'h3 : _btb_79_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_79_bht_T_27 = _btb_79_bht_T_1 ? 2'h1 : _btb_79_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9022 = btb_79_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6735; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9024 = btb_79_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_79_bht_T_27 : _GEN_8271; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_80_bht_T = btb_80_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_80_bht_T_1 = io_i_branch_resolve_pack_taken & btb_80_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_80_bht_T_2 = btb_80_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_80_bht_T_3 = io_i_branch_resolve_pack_taken & btb_80_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_80_bht_T_4 = btb_80_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_80_bht_T_5 = io_i_branch_resolve_pack_taken & btb_80_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_80_bht_T_6 = btb_80_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_80_bht_T_7 = io_i_branch_resolve_pack_taken & btb_80_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_80_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_80_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_80_bht_T_13 = _btb_0_bht_T_8 & _btb_80_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_80_bht_T_16 = _btb_0_bht_T_8 & _btb_80_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_80_bht_T_19 = _btb_0_bht_T_8 & _btb_80_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_80_bht_T_20 = _btb_80_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_21 = _btb_80_bht_T_16 ? 2'h0 : _btb_80_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_22 = _btb_80_bht_T_13 ? 2'h0 : _btb_80_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_23 = _btb_80_bht_T_10 ? 2'h0 : _btb_80_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_24 = _btb_80_bht_T_7 ? 2'h3 : _btb_80_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_25 = _btb_80_bht_T_5 ? 2'h3 : _btb_80_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_26 = _btb_80_bht_T_3 ? 2'h3 : _btb_80_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_80_bht_T_27 = _btb_80_bht_T_1 ? 2'h1 : _btb_80_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9026 = btb_80_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6736; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9028 = btb_80_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_80_bht_T_27 : _GEN_8272; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_81_bht_T = btb_81_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_81_bht_T_1 = io_i_branch_resolve_pack_taken & btb_81_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_81_bht_T_2 = btb_81_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_81_bht_T_3 = io_i_branch_resolve_pack_taken & btb_81_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_81_bht_T_4 = btb_81_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_81_bht_T_5 = io_i_branch_resolve_pack_taken & btb_81_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_81_bht_T_6 = btb_81_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_81_bht_T_7 = io_i_branch_resolve_pack_taken & btb_81_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_81_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_81_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_81_bht_T_13 = _btb_0_bht_T_8 & _btb_81_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_81_bht_T_16 = _btb_0_bht_T_8 & _btb_81_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_81_bht_T_19 = _btb_0_bht_T_8 & _btb_81_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_81_bht_T_20 = _btb_81_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_21 = _btb_81_bht_T_16 ? 2'h0 : _btb_81_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_22 = _btb_81_bht_T_13 ? 2'h0 : _btb_81_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_23 = _btb_81_bht_T_10 ? 2'h0 : _btb_81_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_24 = _btb_81_bht_T_7 ? 2'h3 : _btb_81_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_25 = _btb_81_bht_T_5 ? 2'h3 : _btb_81_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_26 = _btb_81_bht_T_3 ? 2'h3 : _btb_81_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_81_bht_T_27 = _btb_81_bht_T_1 ? 2'h1 : _btb_81_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9030 = btb_81_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6737; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9032 = btb_81_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_81_bht_T_27 : _GEN_8273; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_82_bht_T = btb_82_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_82_bht_T_1 = io_i_branch_resolve_pack_taken & btb_82_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_82_bht_T_2 = btb_82_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_82_bht_T_3 = io_i_branch_resolve_pack_taken & btb_82_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_82_bht_T_4 = btb_82_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_82_bht_T_5 = io_i_branch_resolve_pack_taken & btb_82_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_82_bht_T_6 = btb_82_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_82_bht_T_7 = io_i_branch_resolve_pack_taken & btb_82_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_82_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_82_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_82_bht_T_13 = _btb_0_bht_T_8 & _btb_82_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_82_bht_T_16 = _btb_0_bht_T_8 & _btb_82_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_82_bht_T_19 = _btb_0_bht_T_8 & _btb_82_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_82_bht_T_20 = _btb_82_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_21 = _btb_82_bht_T_16 ? 2'h0 : _btb_82_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_22 = _btb_82_bht_T_13 ? 2'h0 : _btb_82_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_23 = _btb_82_bht_T_10 ? 2'h0 : _btb_82_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_24 = _btb_82_bht_T_7 ? 2'h3 : _btb_82_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_25 = _btb_82_bht_T_5 ? 2'h3 : _btb_82_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_26 = _btb_82_bht_T_3 ? 2'h3 : _btb_82_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_82_bht_T_27 = _btb_82_bht_T_1 ? 2'h1 : _btb_82_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9034 = btb_82_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6738; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9036 = btb_82_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_82_bht_T_27 : _GEN_8274; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_83_bht_T = btb_83_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_83_bht_T_1 = io_i_branch_resolve_pack_taken & btb_83_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_83_bht_T_2 = btb_83_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_83_bht_T_3 = io_i_branch_resolve_pack_taken & btb_83_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_83_bht_T_4 = btb_83_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_83_bht_T_5 = io_i_branch_resolve_pack_taken & btb_83_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_83_bht_T_6 = btb_83_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_83_bht_T_7 = io_i_branch_resolve_pack_taken & btb_83_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_83_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_83_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_83_bht_T_13 = _btb_0_bht_T_8 & _btb_83_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_83_bht_T_16 = _btb_0_bht_T_8 & _btb_83_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_83_bht_T_19 = _btb_0_bht_T_8 & _btb_83_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_83_bht_T_20 = _btb_83_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_21 = _btb_83_bht_T_16 ? 2'h0 : _btb_83_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_22 = _btb_83_bht_T_13 ? 2'h0 : _btb_83_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_23 = _btb_83_bht_T_10 ? 2'h0 : _btb_83_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_24 = _btb_83_bht_T_7 ? 2'h3 : _btb_83_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_25 = _btb_83_bht_T_5 ? 2'h3 : _btb_83_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_26 = _btb_83_bht_T_3 ? 2'h3 : _btb_83_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_83_bht_T_27 = _btb_83_bht_T_1 ? 2'h1 : _btb_83_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9038 = btb_83_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6739; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9040 = btb_83_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_83_bht_T_27 : _GEN_8275; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_84_bht_T = btb_84_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_84_bht_T_1 = io_i_branch_resolve_pack_taken & btb_84_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_84_bht_T_2 = btb_84_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_84_bht_T_3 = io_i_branch_resolve_pack_taken & btb_84_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_84_bht_T_4 = btb_84_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_84_bht_T_5 = io_i_branch_resolve_pack_taken & btb_84_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_84_bht_T_6 = btb_84_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_84_bht_T_7 = io_i_branch_resolve_pack_taken & btb_84_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_84_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_84_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_84_bht_T_13 = _btb_0_bht_T_8 & _btb_84_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_84_bht_T_16 = _btb_0_bht_T_8 & _btb_84_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_84_bht_T_19 = _btb_0_bht_T_8 & _btb_84_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_84_bht_T_20 = _btb_84_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_21 = _btb_84_bht_T_16 ? 2'h0 : _btb_84_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_22 = _btb_84_bht_T_13 ? 2'h0 : _btb_84_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_23 = _btb_84_bht_T_10 ? 2'h0 : _btb_84_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_24 = _btb_84_bht_T_7 ? 2'h3 : _btb_84_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_25 = _btb_84_bht_T_5 ? 2'h3 : _btb_84_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_26 = _btb_84_bht_T_3 ? 2'h3 : _btb_84_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_84_bht_T_27 = _btb_84_bht_T_1 ? 2'h1 : _btb_84_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9042 = btb_84_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6740; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9044 = btb_84_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_84_bht_T_27 : _GEN_8276; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_85_bht_T = btb_85_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_85_bht_T_1 = io_i_branch_resolve_pack_taken & btb_85_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_85_bht_T_2 = btb_85_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_85_bht_T_3 = io_i_branch_resolve_pack_taken & btb_85_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_85_bht_T_4 = btb_85_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_85_bht_T_5 = io_i_branch_resolve_pack_taken & btb_85_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_85_bht_T_6 = btb_85_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_85_bht_T_7 = io_i_branch_resolve_pack_taken & btb_85_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_85_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_85_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_85_bht_T_13 = _btb_0_bht_T_8 & _btb_85_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_85_bht_T_16 = _btb_0_bht_T_8 & _btb_85_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_85_bht_T_19 = _btb_0_bht_T_8 & _btb_85_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_85_bht_T_20 = _btb_85_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_21 = _btb_85_bht_T_16 ? 2'h0 : _btb_85_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_22 = _btb_85_bht_T_13 ? 2'h0 : _btb_85_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_23 = _btb_85_bht_T_10 ? 2'h0 : _btb_85_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_24 = _btb_85_bht_T_7 ? 2'h3 : _btb_85_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_25 = _btb_85_bht_T_5 ? 2'h3 : _btb_85_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_26 = _btb_85_bht_T_3 ? 2'h3 : _btb_85_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_85_bht_T_27 = _btb_85_bht_T_1 ? 2'h1 : _btb_85_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9046 = btb_85_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6741; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9048 = btb_85_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_85_bht_T_27 : _GEN_8277; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_86_bht_T = btb_86_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_86_bht_T_1 = io_i_branch_resolve_pack_taken & btb_86_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_86_bht_T_2 = btb_86_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_86_bht_T_3 = io_i_branch_resolve_pack_taken & btb_86_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_86_bht_T_4 = btb_86_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_86_bht_T_5 = io_i_branch_resolve_pack_taken & btb_86_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_86_bht_T_6 = btb_86_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_86_bht_T_7 = io_i_branch_resolve_pack_taken & btb_86_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_86_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_86_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_86_bht_T_13 = _btb_0_bht_T_8 & _btb_86_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_86_bht_T_16 = _btb_0_bht_T_8 & _btb_86_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_86_bht_T_19 = _btb_0_bht_T_8 & _btb_86_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_86_bht_T_20 = _btb_86_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_21 = _btb_86_bht_T_16 ? 2'h0 : _btb_86_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_22 = _btb_86_bht_T_13 ? 2'h0 : _btb_86_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_23 = _btb_86_bht_T_10 ? 2'h0 : _btb_86_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_24 = _btb_86_bht_T_7 ? 2'h3 : _btb_86_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_25 = _btb_86_bht_T_5 ? 2'h3 : _btb_86_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_26 = _btb_86_bht_T_3 ? 2'h3 : _btb_86_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_86_bht_T_27 = _btb_86_bht_T_1 ? 2'h1 : _btb_86_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9050 = btb_86_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6742; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9052 = btb_86_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_86_bht_T_27 : _GEN_8278; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_87_bht_T = btb_87_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_87_bht_T_1 = io_i_branch_resolve_pack_taken & btb_87_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_87_bht_T_2 = btb_87_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_87_bht_T_3 = io_i_branch_resolve_pack_taken & btb_87_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_87_bht_T_4 = btb_87_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_87_bht_T_5 = io_i_branch_resolve_pack_taken & btb_87_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_87_bht_T_6 = btb_87_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_87_bht_T_7 = io_i_branch_resolve_pack_taken & btb_87_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_87_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_87_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_87_bht_T_13 = _btb_0_bht_T_8 & _btb_87_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_87_bht_T_16 = _btb_0_bht_T_8 & _btb_87_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_87_bht_T_19 = _btb_0_bht_T_8 & _btb_87_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_87_bht_T_20 = _btb_87_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_21 = _btb_87_bht_T_16 ? 2'h0 : _btb_87_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_22 = _btb_87_bht_T_13 ? 2'h0 : _btb_87_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_23 = _btb_87_bht_T_10 ? 2'h0 : _btb_87_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_24 = _btb_87_bht_T_7 ? 2'h3 : _btb_87_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_25 = _btb_87_bht_T_5 ? 2'h3 : _btb_87_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_26 = _btb_87_bht_T_3 ? 2'h3 : _btb_87_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_87_bht_T_27 = _btb_87_bht_T_1 ? 2'h1 : _btb_87_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9054 = btb_87_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6743; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9056 = btb_87_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_87_bht_T_27 : _GEN_8279; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_88_bht_T = btb_88_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_88_bht_T_1 = io_i_branch_resolve_pack_taken & btb_88_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_88_bht_T_2 = btb_88_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_88_bht_T_3 = io_i_branch_resolve_pack_taken & btb_88_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_88_bht_T_4 = btb_88_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_88_bht_T_5 = io_i_branch_resolve_pack_taken & btb_88_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_88_bht_T_6 = btb_88_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_88_bht_T_7 = io_i_branch_resolve_pack_taken & btb_88_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_88_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_88_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_88_bht_T_13 = _btb_0_bht_T_8 & _btb_88_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_88_bht_T_16 = _btb_0_bht_T_8 & _btb_88_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_88_bht_T_19 = _btb_0_bht_T_8 & _btb_88_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_88_bht_T_20 = _btb_88_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_21 = _btb_88_bht_T_16 ? 2'h0 : _btb_88_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_22 = _btb_88_bht_T_13 ? 2'h0 : _btb_88_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_23 = _btb_88_bht_T_10 ? 2'h0 : _btb_88_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_24 = _btb_88_bht_T_7 ? 2'h3 : _btb_88_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_25 = _btb_88_bht_T_5 ? 2'h3 : _btb_88_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_26 = _btb_88_bht_T_3 ? 2'h3 : _btb_88_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_88_bht_T_27 = _btb_88_bht_T_1 ? 2'h1 : _btb_88_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9058 = btb_88_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6744; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9060 = btb_88_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_88_bht_T_27 : _GEN_8280; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_89_bht_T = btb_89_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_89_bht_T_1 = io_i_branch_resolve_pack_taken & btb_89_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_89_bht_T_2 = btb_89_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_89_bht_T_3 = io_i_branch_resolve_pack_taken & btb_89_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_89_bht_T_4 = btb_89_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_89_bht_T_5 = io_i_branch_resolve_pack_taken & btb_89_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_89_bht_T_6 = btb_89_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_89_bht_T_7 = io_i_branch_resolve_pack_taken & btb_89_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_89_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_89_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_89_bht_T_13 = _btb_0_bht_T_8 & _btb_89_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_89_bht_T_16 = _btb_0_bht_T_8 & _btb_89_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_89_bht_T_19 = _btb_0_bht_T_8 & _btb_89_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_89_bht_T_20 = _btb_89_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_21 = _btb_89_bht_T_16 ? 2'h0 : _btb_89_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_22 = _btb_89_bht_T_13 ? 2'h0 : _btb_89_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_23 = _btb_89_bht_T_10 ? 2'h0 : _btb_89_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_24 = _btb_89_bht_T_7 ? 2'h3 : _btb_89_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_25 = _btb_89_bht_T_5 ? 2'h3 : _btb_89_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_26 = _btb_89_bht_T_3 ? 2'h3 : _btb_89_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_89_bht_T_27 = _btb_89_bht_T_1 ? 2'h1 : _btb_89_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9061 = btb_89_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_88_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_87_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_86_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_85_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_84_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_83_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_82_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_81_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_80_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_79_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_78_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_77_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_76_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_75_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9001)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9062 = btb_89_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6745; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9064 = btb_89_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_89_bht_T_27 : _GEN_8281; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_90_bht_T = btb_90_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_90_bht_T_1 = io_i_branch_resolve_pack_taken & btb_90_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_90_bht_T_2 = btb_90_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_90_bht_T_3 = io_i_branch_resolve_pack_taken & btb_90_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_90_bht_T_4 = btb_90_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_90_bht_T_5 = io_i_branch_resolve_pack_taken & btb_90_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_90_bht_T_6 = btb_90_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_90_bht_T_7 = io_i_branch_resolve_pack_taken & btb_90_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_90_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_90_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_90_bht_T_13 = _btb_0_bht_T_8 & _btb_90_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_90_bht_T_16 = _btb_0_bht_T_8 & _btb_90_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_90_bht_T_19 = _btb_0_bht_T_8 & _btb_90_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_90_bht_T_20 = _btb_90_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_21 = _btb_90_bht_T_16 ? 2'h0 : _btb_90_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_22 = _btb_90_bht_T_13 ? 2'h0 : _btb_90_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_23 = _btb_90_bht_T_10 ? 2'h0 : _btb_90_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_24 = _btb_90_bht_T_7 ? 2'h3 : _btb_90_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_25 = _btb_90_bht_T_5 ? 2'h3 : _btb_90_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_26 = _btb_90_bht_T_3 ? 2'h3 : _btb_90_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_90_bht_T_27 = _btb_90_bht_T_1 ? 2'h1 : _btb_90_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9066 = btb_90_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6746; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9068 = btb_90_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_90_bht_T_27 : _GEN_8282; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_91_bht_T = btb_91_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_91_bht_T_1 = io_i_branch_resolve_pack_taken & btb_91_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_91_bht_T_2 = btb_91_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_91_bht_T_3 = io_i_branch_resolve_pack_taken & btb_91_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_91_bht_T_4 = btb_91_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_91_bht_T_5 = io_i_branch_resolve_pack_taken & btb_91_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_91_bht_T_6 = btb_91_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_91_bht_T_7 = io_i_branch_resolve_pack_taken & btb_91_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_91_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_91_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_91_bht_T_13 = _btb_0_bht_T_8 & _btb_91_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_91_bht_T_16 = _btb_0_bht_T_8 & _btb_91_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_91_bht_T_19 = _btb_0_bht_T_8 & _btb_91_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_91_bht_T_20 = _btb_91_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_21 = _btb_91_bht_T_16 ? 2'h0 : _btb_91_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_22 = _btb_91_bht_T_13 ? 2'h0 : _btb_91_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_23 = _btb_91_bht_T_10 ? 2'h0 : _btb_91_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_24 = _btb_91_bht_T_7 ? 2'h3 : _btb_91_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_25 = _btb_91_bht_T_5 ? 2'h3 : _btb_91_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_26 = _btb_91_bht_T_3 ? 2'h3 : _btb_91_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_91_bht_T_27 = _btb_91_bht_T_1 ? 2'h1 : _btb_91_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9070 = btb_91_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6747; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9072 = btb_91_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_91_bht_T_27 : _GEN_8283; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_92_bht_T = btb_92_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_92_bht_T_1 = io_i_branch_resolve_pack_taken & btb_92_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_92_bht_T_2 = btb_92_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_92_bht_T_3 = io_i_branch_resolve_pack_taken & btb_92_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_92_bht_T_4 = btb_92_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_92_bht_T_5 = io_i_branch_resolve_pack_taken & btb_92_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_92_bht_T_6 = btb_92_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_92_bht_T_7 = io_i_branch_resolve_pack_taken & btb_92_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_92_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_92_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_92_bht_T_13 = _btb_0_bht_T_8 & _btb_92_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_92_bht_T_16 = _btb_0_bht_T_8 & _btb_92_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_92_bht_T_19 = _btb_0_bht_T_8 & _btb_92_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_92_bht_T_20 = _btb_92_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_21 = _btb_92_bht_T_16 ? 2'h0 : _btb_92_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_22 = _btb_92_bht_T_13 ? 2'h0 : _btb_92_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_23 = _btb_92_bht_T_10 ? 2'h0 : _btb_92_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_24 = _btb_92_bht_T_7 ? 2'h3 : _btb_92_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_25 = _btb_92_bht_T_5 ? 2'h3 : _btb_92_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_26 = _btb_92_bht_T_3 ? 2'h3 : _btb_92_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_92_bht_T_27 = _btb_92_bht_T_1 ? 2'h1 : _btb_92_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9074 = btb_92_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6748; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9076 = btb_92_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_92_bht_T_27 : _GEN_8284; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_93_bht_T = btb_93_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_93_bht_T_1 = io_i_branch_resolve_pack_taken & btb_93_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_93_bht_T_2 = btb_93_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_93_bht_T_3 = io_i_branch_resolve_pack_taken & btb_93_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_93_bht_T_4 = btb_93_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_93_bht_T_5 = io_i_branch_resolve_pack_taken & btb_93_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_93_bht_T_6 = btb_93_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_93_bht_T_7 = io_i_branch_resolve_pack_taken & btb_93_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_93_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_93_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_93_bht_T_13 = _btb_0_bht_T_8 & _btb_93_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_93_bht_T_16 = _btb_0_bht_T_8 & _btb_93_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_93_bht_T_19 = _btb_0_bht_T_8 & _btb_93_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_93_bht_T_20 = _btb_93_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_21 = _btb_93_bht_T_16 ? 2'h0 : _btb_93_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_22 = _btb_93_bht_T_13 ? 2'h0 : _btb_93_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_23 = _btb_93_bht_T_10 ? 2'h0 : _btb_93_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_24 = _btb_93_bht_T_7 ? 2'h3 : _btb_93_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_25 = _btb_93_bht_T_5 ? 2'h3 : _btb_93_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_26 = _btb_93_bht_T_3 ? 2'h3 : _btb_93_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_93_bht_T_27 = _btb_93_bht_T_1 ? 2'h1 : _btb_93_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9078 = btb_93_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6749; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9080 = btb_93_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_93_bht_T_27 : _GEN_8285; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_94_bht_T = btb_94_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_94_bht_T_1 = io_i_branch_resolve_pack_taken & btb_94_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_94_bht_T_2 = btb_94_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_94_bht_T_3 = io_i_branch_resolve_pack_taken & btb_94_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_94_bht_T_4 = btb_94_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_94_bht_T_5 = io_i_branch_resolve_pack_taken & btb_94_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_94_bht_T_6 = btb_94_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_94_bht_T_7 = io_i_branch_resolve_pack_taken & btb_94_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_94_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_94_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_94_bht_T_13 = _btb_0_bht_T_8 & _btb_94_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_94_bht_T_16 = _btb_0_bht_T_8 & _btb_94_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_94_bht_T_19 = _btb_0_bht_T_8 & _btb_94_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_94_bht_T_20 = _btb_94_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_21 = _btb_94_bht_T_16 ? 2'h0 : _btb_94_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_22 = _btb_94_bht_T_13 ? 2'h0 : _btb_94_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_23 = _btb_94_bht_T_10 ? 2'h0 : _btb_94_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_24 = _btb_94_bht_T_7 ? 2'h3 : _btb_94_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_25 = _btb_94_bht_T_5 ? 2'h3 : _btb_94_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_26 = _btb_94_bht_T_3 ? 2'h3 : _btb_94_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_94_bht_T_27 = _btb_94_bht_T_1 ? 2'h1 : _btb_94_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9082 = btb_94_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6750; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9084 = btb_94_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_94_bht_T_27 : _GEN_8286; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_95_bht_T = btb_95_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_95_bht_T_1 = io_i_branch_resolve_pack_taken & btb_95_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_95_bht_T_2 = btb_95_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_95_bht_T_3 = io_i_branch_resolve_pack_taken & btb_95_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_95_bht_T_4 = btb_95_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_95_bht_T_5 = io_i_branch_resolve_pack_taken & btb_95_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_95_bht_T_6 = btb_95_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_95_bht_T_7 = io_i_branch_resolve_pack_taken & btb_95_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_95_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_95_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_95_bht_T_13 = _btb_0_bht_T_8 & _btb_95_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_95_bht_T_16 = _btb_0_bht_T_8 & _btb_95_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_95_bht_T_19 = _btb_0_bht_T_8 & _btb_95_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_95_bht_T_20 = _btb_95_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_21 = _btb_95_bht_T_16 ? 2'h0 : _btb_95_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_22 = _btb_95_bht_T_13 ? 2'h0 : _btb_95_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_23 = _btb_95_bht_T_10 ? 2'h0 : _btb_95_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_24 = _btb_95_bht_T_7 ? 2'h3 : _btb_95_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_25 = _btb_95_bht_T_5 ? 2'h3 : _btb_95_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_26 = _btb_95_bht_T_3 ? 2'h3 : _btb_95_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_95_bht_T_27 = _btb_95_bht_T_1 ? 2'h1 : _btb_95_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9086 = btb_95_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6751; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9088 = btb_95_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_95_bht_T_27 : _GEN_8287; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_96_bht_T = btb_96_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_96_bht_T_1 = io_i_branch_resolve_pack_taken & btb_96_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_96_bht_T_2 = btb_96_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_96_bht_T_3 = io_i_branch_resolve_pack_taken & btb_96_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_96_bht_T_4 = btb_96_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_96_bht_T_5 = io_i_branch_resolve_pack_taken & btb_96_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_96_bht_T_6 = btb_96_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_96_bht_T_7 = io_i_branch_resolve_pack_taken & btb_96_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_96_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_96_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_96_bht_T_13 = _btb_0_bht_T_8 & _btb_96_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_96_bht_T_16 = _btb_0_bht_T_8 & _btb_96_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_96_bht_T_19 = _btb_0_bht_T_8 & _btb_96_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_96_bht_T_20 = _btb_96_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_21 = _btb_96_bht_T_16 ? 2'h0 : _btb_96_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_22 = _btb_96_bht_T_13 ? 2'h0 : _btb_96_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_23 = _btb_96_bht_T_10 ? 2'h0 : _btb_96_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_24 = _btb_96_bht_T_7 ? 2'h3 : _btb_96_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_25 = _btb_96_bht_T_5 ? 2'h3 : _btb_96_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_26 = _btb_96_bht_T_3 ? 2'h3 : _btb_96_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_96_bht_T_27 = _btb_96_bht_T_1 ? 2'h1 : _btb_96_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9090 = btb_96_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6752; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9092 = btb_96_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_96_bht_T_27 : _GEN_8288; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_97_bht_T = btb_97_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_97_bht_T_1 = io_i_branch_resolve_pack_taken & btb_97_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_97_bht_T_2 = btb_97_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_97_bht_T_3 = io_i_branch_resolve_pack_taken & btb_97_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_97_bht_T_4 = btb_97_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_97_bht_T_5 = io_i_branch_resolve_pack_taken & btb_97_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_97_bht_T_6 = btb_97_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_97_bht_T_7 = io_i_branch_resolve_pack_taken & btb_97_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_97_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_97_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_97_bht_T_13 = _btb_0_bht_T_8 & _btb_97_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_97_bht_T_16 = _btb_0_bht_T_8 & _btb_97_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_97_bht_T_19 = _btb_0_bht_T_8 & _btb_97_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_97_bht_T_20 = _btb_97_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_21 = _btb_97_bht_T_16 ? 2'h0 : _btb_97_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_22 = _btb_97_bht_T_13 ? 2'h0 : _btb_97_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_23 = _btb_97_bht_T_10 ? 2'h0 : _btb_97_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_24 = _btb_97_bht_T_7 ? 2'h3 : _btb_97_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_25 = _btb_97_bht_T_5 ? 2'h3 : _btb_97_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_26 = _btb_97_bht_T_3 ? 2'h3 : _btb_97_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_97_bht_T_27 = _btb_97_bht_T_1 ? 2'h1 : _btb_97_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9094 = btb_97_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6753; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9096 = btb_97_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_97_bht_T_27 : _GEN_8289; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_98_bht_T = btb_98_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_98_bht_T_1 = io_i_branch_resolve_pack_taken & btb_98_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_98_bht_T_2 = btb_98_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_98_bht_T_3 = io_i_branch_resolve_pack_taken & btb_98_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_98_bht_T_4 = btb_98_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_98_bht_T_5 = io_i_branch_resolve_pack_taken & btb_98_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_98_bht_T_6 = btb_98_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_98_bht_T_7 = io_i_branch_resolve_pack_taken & btb_98_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_98_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_98_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_98_bht_T_13 = _btb_0_bht_T_8 & _btb_98_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_98_bht_T_16 = _btb_0_bht_T_8 & _btb_98_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_98_bht_T_19 = _btb_0_bht_T_8 & _btb_98_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_98_bht_T_20 = _btb_98_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_21 = _btb_98_bht_T_16 ? 2'h0 : _btb_98_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_22 = _btb_98_bht_T_13 ? 2'h0 : _btb_98_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_23 = _btb_98_bht_T_10 ? 2'h0 : _btb_98_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_24 = _btb_98_bht_T_7 ? 2'h3 : _btb_98_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_25 = _btb_98_bht_T_5 ? 2'h3 : _btb_98_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_26 = _btb_98_bht_T_3 ? 2'h3 : _btb_98_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_98_bht_T_27 = _btb_98_bht_T_1 ? 2'h1 : _btb_98_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9098 = btb_98_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6754; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9100 = btb_98_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_98_bht_T_27 : _GEN_8290; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_99_bht_T = btb_99_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_99_bht_T_1 = io_i_branch_resolve_pack_taken & btb_99_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_99_bht_T_2 = btb_99_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_99_bht_T_3 = io_i_branch_resolve_pack_taken & btb_99_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_99_bht_T_4 = btb_99_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_99_bht_T_5 = io_i_branch_resolve_pack_taken & btb_99_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_99_bht_T_6 = btb_99_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_99_bht_T_7 = io_i_branch_resolve_pack_taken & btb_99_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_99_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_99_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_99_bht_T_13 = _btb_0_bht_T_8 & _btb_99_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_99_bht_T_16 = _btb_0_bht_T_8 & _btb_99_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_99_bht_T_19 = _btb_0_bht_T_8 & _btb_99_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_99_bht_T_20 = _btb_99_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_21 = _btb_99_bht_T_16 ? 2'h0 : _btb_99_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_22 = _btb_99_bht_T_13 ? 2'h0 : _btb_99_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_23 = _btb_99_bht_T_10 ? 2'h0 : _btb_99_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_24 = _btb_99_bht_T_7 ? 2'h3 : _btb_99_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_25 = _btb_99_bht_T_5 ? 2'h3 : _btb_99_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_26 = _btb_99_bht_T_3 ? 2'h3 : _btb_99_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_99_bht_T_27 = _btb_99_bht_T_1 ? 2'h1 : _btb_99_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9102 = btb_99_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6755; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9104 = btb_99_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_99_bht_T_27 : _GEN_8291; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_100_bht_T = btb_100_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_100_bht_T_1 = io_i_branch_resolve_pack_taken & btb_100_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_100_bht_T_2 = btb_100_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_100_bht_T_3 = io_i_branch_resolve_pack_taken & btb_100_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_100_bht_T_4 = btb_100_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_100_bht_T_5 = io_i_branch_resolve_pack_taken & btb_100_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_100_bht_T_6 = btb_100_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_100_bht_T_7 = io_i_branch_resolve_pack_taken & btb_100_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_100_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_100_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_100_bht_T_13 = _btb_0_bht_T_8 & _btb_100_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_100_bht_T_16 = _btb_0_bht_T_8 & _btb_100_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_100_bht_T_19 = _btb_0_bht_T_8 & _btb_100_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_100_bht_T_20 = _btb_100_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_21 = _btb_100_bht_T_16 ? 2'h0 : _btb_100_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_22 = _btb_100_bht_T_13 ? 2'h0 : _btb_100_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_23 = _btb_100_bht_T_10 ? 2'h0 : _btb_100_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_24 = _btb_100_bht_T_7 ? 2'h3 : _btb_100_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_25 = _btb_100_bht_T_5 ? 2'h3 : _btb_100_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_26 = _btb_100_bht_T_3 ? 2'h3 : _btb_100_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_100_bht_T_27 = _btb_100_bht_T_1 ? 2'h1 : _btb_100_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9106 = btb_100_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6756
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9108 = btb_100_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_100_bht_T_27 : _GEN_8292; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_101_bht_T = btb_101_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_101_bht_T_1 = io_i_branch_resolve_pack_taken & btb_101_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_101_bht_T_2 = btb_101_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_101_bht_T_3 = io_i_branch_resolve_pack_taken & btb_101_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_101_bht_T_4 = btb_101_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_101_bht_T_5 = io_i_branch_resolve_pack_taken & btb_101_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_101_bht_T_6 = btb_101_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_101_bht_T_7 = io_i_branch_resolve_pack_taken & btb_101_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_101_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_101_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_101_bht_T_13 = _btb_0_bht_T_8 & _btb_101_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_101_bht_T_16 = _btb_0_bht_T_8 & _btb_101_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_101_bht_T_19 = _btb_0_bht_T_8 & _btb_101_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_101_bht_T_20 = _btb_101_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_21 = _btb_101_bht_T_16 ? 2'h0 : _btb_101_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_22 = _btb_101_bht_T_13 ? 2'h0 : _btb_101_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_23 = _btb_101_bht_T_10 ? 2'h0 : _btb_101_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_24 = _btb_101_bht_T_7 ? 2'h3 : _btb_101_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_25 = _btb_101_bht_T_5 ? 2'h3 : _btb_101_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_26 = _btb_101_bht_T_3 ? 2'h3 : _btb_101_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_101_bht_T_27 = _btb_101_bht_T_1 ? 2'h1 : _btb_101_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9110 = btb_101_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6757
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9112 = btb_101_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_101_bht_T_27 : _GEN_8293; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_102_bht_T = btb_102_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_102_bht_T_1 = io_i_branch_resolve_pack_taken & btb_102_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_102_bht_T_2 = btb_102_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_102_bht_T_3 = io_i_branch_resolve_pack_taken & btb_102_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_102_bht_T_4 = btb_102_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_102_bht_T_5 = io_i_branch_resolve_pack_taken & btb_102_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_102_bht_T_6 = btb_102_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_102_bht_T_7 = io_i_branch_resolve_pack_taken & btb_102_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_102_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_102_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_102_bht_T_13 = _btb_0_bht_T_8 & _btb_102_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_102_bht_T_16 = _btb_0_bht_T_8 & _btb_102_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_102_bht_T_19 = _btb_0_bht_T_8 & _btb_102_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_102_bht_T_20 = _btb_102_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_21 = _btb_102_bht_T_16 ? 2'h0 : _btb_102_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_22 = _btb_102_bht_T_13 ? 2'h0 : _btb_102_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_23 = _btb_102_bht_T_10 ? 2'h0 : _btb_102_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_24 = _btb_102_bht_T_7 ? 2'h3 : _btb_102_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_25 = _btb_102_bht_T_5 ? 2'h3 : _btb_102_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_26 = _btb_102_bht_T_3 ? 2'h3 : _btb_102_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_102_bht_T_27 = _btb_102_bht_T_1 ? 2'h1 : _btb_102_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9114 = btb_102_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6758
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9116 = btb_102_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_102_bht_T_27 : _GEN_8294; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_103_bht_T = btb_103_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_103_bht_T_1 = io_i_branch_resolve_pack_taken & btb_103_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_103_bht_T_2 = btb_103_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_103_bht_T_3 = io_i_branch_resolve_pack_taken & btb_103_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_103_bht_T_4 = btb_103_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_103_bht_T_5 = io_i_branch_resolve_pack_taken & btb_103_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_103_bht_T_6 = btb_103_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_103_bht_T_7 = io_i_branch_resolve_pack_taken & btb_103_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_103_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_103_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_103_bht_T_13 = _btb_0_bht_T_8 & _btb_103_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_103_bht_T_16 = _btb_0_bht_T_8 & _btb_103_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_103_bht_T_19 = _btb_0_bht_T_8 & _btb_103_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_103_bht_T_20 = _btb_103_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_21 = _btb_103_bht_T_16 ? 2'h0 : _btb_103_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_22 = _btb_103_bht_T_13 ? 2'h0 : _btb_103_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_23 = _btb_103_bht_T_10 ? 2'h0 : _btb_103_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_24 = _btb_103_bht_T_7 ? 2'h3 : _btb_103_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_25 = _btb_103_bht_T_5 ? 2'h3 : _btb_103_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_26 = _btb_103_bht_T_3 ? 2'h3 : _btb_103_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_103_bht_T_27 = _btb_103_bht_T_1 ? 2'h1 : _btb_103_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9118 = btb_103_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6759
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9120 = btb_103_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_103_bht_T_27 : _GEN_8295; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_104_bht_T = btb_104_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_104_bht_T_1 = io_i_branch_resolve_pack_taken & btb_104_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_104_bht_T_2 = btb_104_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_104_bht_T_3 = io_i_branch_resolve_pack_taken & btb_104_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_104_bht_T_4 = btb_104_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_104_bht_T_5 = io_i_branch_resolve_pack_taken & btb_104_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_104_bht_T_6 = btb_104_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_104_bht_T_7 = io_i_branch_resolve_pack_taken & btb_104_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_104_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_104_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_104_bht_T_13 = _btb_0_bht_T_8 & _btb_104_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_104_bht_T_16 = _btb_0_bht_T_8 & _btb_104_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_104_bht_T_19 = _btb_0_bht_T_8 & _btb_104_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_104_bht_T_20 = _btb_104_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_21 = _btb_104_bht_T_16 ? 2'h0 : _btb_104_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_22 = _btb_104_bht_T_13 ? 2'h0 : _btb_104_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_23 = _btb_104_bht_T_10 ? 2'h0 : _btb_104_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_24 = _btb_104_bht_T_7 ? 2'h3 : _btb_104_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_25 = _btb_104_bht_T_5 ? 2'h3 : _btb_104_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_26 = _btb_104_bht_T_3 ? 2'h3 : _btb_104_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_104_bht_T_27 = _btb_104_bht_T_1 ? 2'h1 : _btb_104_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9121 = btb_104_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_103_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_102_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_101_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_100_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_99_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_98_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_97_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_96_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_95_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_94_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_93_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_92_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_91_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_90_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9061)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9122 = btb_104_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6760
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9124 = btb_104_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_104_bht_T_27 : _GEN_8296; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_105_bht_T = btb_105_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_105_bht_T_1 = io_i_branch_resolve_pack_taken & btb_105_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_105_bht_T_2 = btb_105_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_105_bht_T_3 = io_i_branch_resolve_pack_taken & btb_105_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_105_bht_T_4 = btb_105_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_105_bht_T_5 = io_i_branch_resolve_pack_taken & btb_105_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_105_bht_T_6 = btb_105_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_105_bht_T_7 = io_i_branch_resolve_pack_taken & btb_105_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_105_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_105_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_105_bht_T_13 = _btb_0_bht_T_8 & _btb_105_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_105_bht_T_16 = _btb_0_bht_T_8 & _btb_105_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_105_bht_T_19 = _btb_0_bht_T_8 & _btb_105_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_105_bht_T_20 = _btb_105_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_21 = _btb_105_bht_T_16 ? 2'h0 : _btb_105_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_22 = _btb_105_bht_T_13 ? 2'h0 : _btb_105_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_23 = _btb_105_bht_T_10 ? 2'h0 : _btb_105_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_24 = _btb_105_bht_T_7 ? 2'h3 : _btb_105_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_25 = _btb_105_bht_T_5 ? 2'h3 : _btb_105_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_26 = _btb_105_bht_T_3 ? 2'h3 : _btb_105_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_105_bht_T_27 = _btb_105_bht_T_1 ? 2'h1 : _btb_105_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9126 = btb_105_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6761
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9128 = btb_105_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_105_bht_T_27 : _GEN_8297; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_106_bht_T = btb_106_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_106_bht_T_1 = io_i_branch_resolve_pack_taken & btb_106_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_106_bht_T_2 = btb_106_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_106_bht_T_3 = io_i_branch_resolve_pack_taken & btb_106_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_106_bht_T_4 = btb_106_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_106_bht_T_5 = io_i_branch_resolve_pack_taken & btb_106_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_106_bht_T_6 = btb_106_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_106_bht_T_7 = io_i_branch_resolve_pack_taken & btb_106_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_106_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_106_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_106_bht_T_13 = _btb_0_bht_T_8 & _btb_106_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_106_bht_T_16 = _btb_0_bht_T_8 & _btb_106_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_106_bht_T_19 = _btb_0_bht_T_8 & _btb_106_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_106_bht_T_20 = _btb_106_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_21 = _btb_106_bht_T_16 ? 2'h0 : _btb_106_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_22 = _btb_106_bht_T_13 ? 2'h0 : _btb_106_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_23 = _btb_106_bht_T_10 ? 2'h0 : _btb_106_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_24 = _btb_106_bht_T_7 ? 2'h3 : _btb_106_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_25 = _btb_106_bht_T_5 ? 2'h3 : _btb_106_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_26 = _btb_106_bht_T_3 ? 2'h3 : _btb_106_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_106_bht_T_27 = _btb_106_bht_T_1 ? 2'h1 : _btb_106_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9130 = btb_106_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6762
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9132 = btb_106_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_106_bht_T_27 : _GEN_8298; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_107_bht_T = btb_107_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_107_bht_T_1 = io_i_branch_resolve_pack_taken & btb_107_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_107_bht_T_2 = btb_107_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_107_bht_T_3 = io_i_branch_resolve_pack_taken & btb_107_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_107_bht_T_4 = btb_107_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_107_bht_T_5 = io_i_branch_resolve_pack_taken & btb_107_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_107_bht_T_6 = btb_107_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_107_bht_T_7 = io_i_branch_resolve_pack_taken & btb_107_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_107_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_107_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_107_bht_T_13 = _btb_0_bht_T_8 & _btb_107_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_107_bht_T_16 = _btb_0_bht_T_8 & _btb_107_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_107_bht_T_19 = _btb_0_bht_T_8 & _btb_107_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_107_bht_T_20 = _btb_107_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_21 = _btb_107_bht_T_16 ? 2'h0 : _btb_107_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_22 = _btb_107_bht_T_13 ? 2'h0 : _btb_107_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_23 = _btb_107_bht_T_10 ? 2'h0 : _btb_107_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_24 = _btb_107_bht_T_7 ? 2'h3 : _btb_107_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_25 = _btb_107_bht_T_5 ? 2'h3 : _btb_107_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_26 = _btb_107_bht_T_3 ? 2'h3 : _btb_107_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_107_bht_T_27 = _btb_107_bht_T_1 ? 2'h1 : _btb_107_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9134 = btb_107_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6763
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9136 = btb_107_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_107_bht_T_27 : _GEN_8299; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_108_bht_T = btb_108_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_108_bht_T_1 = io_i_branch_resolve_pack_taken & btb_108_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_108_bht_T_2 = btb_108_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_108_bht_T_3 = io_i_branch_resolve_pack_taken & btb_108_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_108_bht_T_4 = btb_108_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_108_bht_T_5 = io_i_branch_resolve_pack_taken & btb_108_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_108_bht_T_6 = btb_108_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_108_bht_T_7 = io_i_branch_resolve_pack_taken & btb_108_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_108_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_108_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_108_bht_T_13 = _btb_0_bht_T_8 & _btb_108_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_108_bht_T_16 = _btb_0_bht_T_8 & _btb_108_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_108_bht_T_19 = _btb_0_bht_T_8 & _btb_108_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_108_bht_T_20 = _btb_108_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_21 = _btb_108_bht_T_16 ? 2'h0 : _btb_108_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_22 = _btb_108_bht_T_13 ? 2'h0 : _btb_108_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_23 = _btb_108_bht_T_10 ? 2'h0 : _btb_108_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_24 = _btb_108_bht_T_7 ? 2'h3 : _btb_108_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_25 = _btb_108_bht_T_5 ? 2'h3 : _btb_108_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_26 = _btb_108_bht_T_3 ? 2'h3 : _btb_108_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_108_bht_T_27 = _btb_108_bht_T_1 ? 2'h1 : _btb_108_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9138 = btb_108_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6764
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9140 = btb_108_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_108_bht_T_27 : _GEN_8300; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_109_bht_T = btb_109_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_109_bht_T_1 = io_i_branch_resolve_pack_taken & btb_109_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_109_bht_T_2 = btb_109_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_109_bht_T_3 = io_i_branch_resolve_pack_taken & btb_109_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_109_bht_T_4 = btb_109_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_109_bht_T_5 = io_i_branch_resolve_pack_taken & btb_109_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_109_bht_T_6 = btb_109_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_109_bht_T_7 = io_i_branch_resolve_pack_taken & btb_109_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_109_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_109_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_109_bht_T_13 = _btb_0_bht_T_8 & _btb_109_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_109_bht_T_16 = _btb_0_bht_T_8 & _btb_109_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_109_bht_T_19 = _btb_0_bht_T_8 & _btb_109_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_109_bht_T_20 = _btb_109_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_21 = _btb_109_bht_T_16 ? 2'h0 : _btb_109_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_22 = _btb_109_bht_T_13 ? 2'h0 : _btb_109_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_23 = _btb_109_bht_T_10 ? 2'h0 : _btb_109_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_24 = _btb_109_bht_T_7 ? 2'h3 : _btb_109_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_25 = _btb_109_bht_T_5 ? 2'h3 : _btb_109_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_26 = _btb_109_bht_T_3 ? 2'h3 : _btb_109_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_109_bht_T_27 = _btb_109_bht_T_1 ? 2'h1 : _btb_109_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9142 = btb_109_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6765
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9144 = btb_109_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_109_bht_T_27 : _GEN_8301; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_110_bht_T = btb_110_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_110_bht_T_1 = io_i_branch_resolve_pack_taken & btb_110_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_110_bht_T_2 = btb_110_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_110_bht_T_3 = io_i_branch_resolve_pack_taken & btb_110_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_110_bht_T_4 = btb_110_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_110_bht_T_5 = io_i_branch_resolve_pack_taken & btb_110_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_110_bht_T_6 = btb_110_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_110_bht_T_7 = io_i_branch_resolve_pack_taken & btb_110_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_110_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_110_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_110_bht_T_13 = _btb_0_bht_T_8 & _btb_110_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_110_bht_T_16 = _btb_0_bht_T_8 & _btb_110_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_110_bht_T_19 = _btb_0_bht_T_8 & _btb_110_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_110_bht_T_20 = _btb_110_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_21 = _btb_110_bht_T_16 ? 2'h0 : _btb_110_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_22 = _btb_110_bht_T_13 ? 2'h0 : _btb_110_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_23 = _btb_110_bht_T_10 ? 2'h0 : _btb_110_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_24 = _btb_110_bht_T_7 ? 2'h3 : _btb_110_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_25 = _btb_110_bht_T_5 ? 2'h3 : _btb_110_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_26 = _btb_110_bht_T_3 ? 2'h3 : _btb_110_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_110_bht_T_27 = _btb_110_bht_T_1 ? 2'h1 : _btb_110_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9146 = btb_110_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6766
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9148 = btb_110_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_110_bht_T_27 : _GEN_8302; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_111_bht_T = btb_111_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_111_bht_T_1 = io_i_branch_resolve_pack_taken & btb_111_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_111_bht_T_2 = btb_111_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_111_bht_T_3 = io_i_branch_resolve_pack_taken & btb_111_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_111_bht_T_4 = btb_111_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_111_bht_T_5 = io_i_branch_resolve_pack_taken & btb_111_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_111_bht_T_6 = btb_111_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_111_bht_T_7 = io_i_branch_resolve_pack_taken & btb_111_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_111_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_111_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_111_bht_T_13 = _btb_0_bht_T_8 & _btb_111_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_111_bht_T_16 = _btb_0_bht_T_8 & _btb_111_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_111_bht_T_19 = _btb_0_bht_T_8 & _btb_111_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_111_bht_T_20 = _btb_111_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_21 = _btb_111_bht_T_16 ? 2'h0 : _btb_111_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_22 = _btb_111_bht_T_13 ? 2'h0 : _btb_111_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_23 = _btb_111_bht_T_10 ? 2'h0 : _btb_111_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_24 = _btb_111_bht_T_7 ? 2'h3 : _btb_111_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_25 = _btb_111_bht_T_5 ? 2'h3 : _btb_111_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_26 = _btb_111_bht_T_3 ? 2'h3 : _btb_111_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_111_bht_T_27 = _btb_111_bht_T_1 ? 2'h1 : _btb_111_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9150 = btb_111_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6767
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9152 = btb_111_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_111_bht_T_27 : _GEN_8303; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_112_bht_T = btb_112_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_112_bht_T_1 = io_i_branch_resolve_pack_taken & btb_112_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_112_bht_T_2 = btb_112_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_112_bht_T_3 = io_i_branch_resolve_pack_taken & btb_112_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_112_bht_T_4 = btb_112_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_112_bht_T_5 = io_i_branch_resolve_pack_taken & btb_112_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_112_bht_T_6 = btb_112_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_112_bht_T_7 = io_i_branch_resolve_pack_taken & btb_112_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_112_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_112_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_112_bht_T_13 = _btb_0_bht_T_8 & _btb_112_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_112_bht_T_16 = _btb_0_bht_T_8 & _btb_112_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_112_bht_T_19 = _btb_0_bht_T_8 & _btb_112_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_112_bht_T_20 = _btb_112_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_21 = _btb_112_bht_T_16 ? 2'h0 : _btb_112_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_22 = _btb_112_bht_T_13 ? 2'h0 : _btb_112_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_23 = _btb_112_bht_T_10 ? 2'h0 : _btb_112_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_24 = _btb_112_bht_T_7 ? 2'h3 : _btb_112_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_25 = _btb_112_bht_T_5 ? 2'h3 : _btb_112_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_26 = _btb_112_bht_T_3 ? 2'h3 : _btb_112_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_112_bht_T_27 = _btb_112_bht_T_1 ? 2'h1 : _btb_112_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9154 = btb_112_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6768
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9156 = btb_112_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_112_bht_T_27 : _GEN_8304; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_113_bht_T = btb_113_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_113_bht_T_1 = io_i_branch_resolve_pack_taken & btb_113_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_113_bht_T_2 = btb_113_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_113_bht_T_3 = io_i_branch_resolve_pack_taken & btb_113_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_113_bht_T_4 = btb_113_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_113_bht_T_5 = io_i_branch_resolve_pack_taken & btb_113_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_113_bht_T_6 = btb_113_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_113_bht_T_7 = io_i_branch_resolve_pack_taken & btb_113_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_113_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_113_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_113_bht_T_13 = _btb_0_bht_T_8 & _btb_113_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_113_bht_T_16 = _btb_0_bht_T_8 & _btb_113_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_113_bht_T_19 = _btb_0_bht_T_8 & _btb_113_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_113_bht_T_20 = _btb_113_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_21 = _btb_113_bht_T_16 ? 2'h0 : _btb_113_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_22 = _btb_113_bht_T_13 ? 2'h0 : _btb_113_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_23 = _btb_113_bht_T_10 ? 2'h0 : _btb_113_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_24 = _btb_113_bht_T_7 ? 2'h3 : _btb_113_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_25 = _btb_113_bht_T_5 ? 2'h3 : _btb_113_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_26 = _btb_113_bht_T_3 ? 2'h3 : _btb_113_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_113_bht_T_27 = _btb_113_bht_T_1 ? 2'h1 : _btb_113_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9158 = btb_113_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6769
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9160 = btb_113_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_113_bht_T_27 : _GEN_8305; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_114_bht_T = btb_114_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_114_bht_T_1 = io_i_branch_resolve_pack_taken & btb_114_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_114_bht_T_2 = btb_114_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_114_bht_T_3 = io_i_branch_resolve_pack_taken & btb_114_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_114_bht_T_4 = btb_114_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_114_bht_T_5 = io_i_branch_resolve_pack_taken & btb_114_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_114_bht_T_6 = btb_114_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_114_bht_T_7 = io_i_branch_resolve_pack_taken & btb_114_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_114_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_114_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_114_bht_T_13 = _btb_0_bht_T_8 & _btb_114_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_114_bht_T_16 = _btb_0_bht_T_8 & _btb_114_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_114_bht_T_19 = _btb_0_bht_T_8 & _btb_114_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_114_bht_T_20 = _btb_114_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_21 = _btb_114_bht_T_16 ? 2'h0 : _btb_114_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_22 = _btb_114_bht_T_13 ? 2'h0 : _btb_114_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_23 = _btb_114_bht_T_10 ? 2'h0 : _btb_114_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_24 = _btb_114_bht_T_7 ? 2'h3 : _btb_114_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_25 = _btb_114_bht_T_5 ? 2'h3 : _btb_114_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_26 = _btb_114_bht_T_3 ? 2'h3 : _btb_114_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_114_bht_T_27 = _btb_114_bht_T_1 ? 2'h1 : _btb_114_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9162 = btb_114_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6770
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9164 = btb_114_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_114_bht_T_27 : _GEN_8306; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_115_bht_T = btb_115_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_115_bht_T_1 = io_i_branch_resolve_pack_taken & btb_115_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_115_bht_T_2 = btb_115_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_115_bht_T_3 = io_i_branch_resolve_pack_taken & btb_115_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_115_bht_T_4 = btb_115_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_115_bht_T_5 = io_i_branch_resolve_pack_taken & btb_115_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_115_bht_T_6 = btb_115_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_115_bht_T_7 = io_i_branch_resolve_pack_taken & btb_115_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_115_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_115_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_115_bht_T_13 = _btb_0_bht_T_8 & _btb_115_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_115_bht_T_16 = _btb_0_bht_T_8 & _btb_115_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_115_bht_T_19 = _btb_0_bht_T_8 & _btb_115_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_115_bht_T_20 = _btb_115_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_21 = _btb_115_bht_T_16 ? 2'h0 : _btb_115_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_22 = _btb_115_bht_T_13 ? 2'h0 : _btb_115_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_23 = _btb_115_bht_T_10 ? 2'h0 : _btb_115_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_24 = _btb_115_bht_T_7 ? 2'h3 : _btb_115_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_25 = _btb_115_bht_T_5 ? 2'h3 : _btb_115_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_26 = _btb_115_bht_T_3 ? 2'h3 : _btb_115_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_115_bht_T_27 = _btb_115_bht_T_1 ? 2'h1 : _btb_115_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9166 = btb_115_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6771
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9168 = btb_115_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_115_bht_T_27 : _GEN_8307; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_116_bht_T = btb_116_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_116_bht_T_1 = io_i_branch_resolve_pack_taken & btb_116_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_116_bht_T_2 = btb_116_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_116_bht_T_3 = io_i_branch_resolve_pack_taken & btb_116_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_116_bht_T_4 = btb_116_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_116_bht_T_5 = io_i_branch_resolve_pack_taken & btb_116_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_116_bht_T_6 = btb_116_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_116_bht_T_7 = io_i_branch_resolve_pack_taken & btb_116_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_116_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_116_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_116_bht_T_13 = _btb_0_bht_T_8 & _btb_116_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_116_bht_T_16 = _btb_0_bht_T_8 & _btb_116_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_116_bht_T_19 = _btb_0_bht_T_8 & _btb_116_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_116_bht_T_20 = _btb_116_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_21 = _btb_116_bht_T_16 ? 2'h0 : _btb_116_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_22 = _btb_116_bht_T_13 ? 2'h0 : _btb_116_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_23 = _btb_116_bht_T_10 ? 2'h0 : _btb_116_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_24 = _btb_116_bht_T_7 ? 2'h3 : _btb_116_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_25 = _btb_116_bht_T_5 ? 2'h3 : _btb_116_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_26 = _btb_116_bht_T_3 ? 2'h3 : _btb_116_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_116_bht_T_27 = _btb_116_bht_T_1 ? 2'h1 : _btb_116_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9170 = btb_116_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6772
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9172 = btb_116_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_116_bht_T_27 : _GEN_8308; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_117_bht_T = btb_117_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_117_bht_T_1 = io_i_branch_resolve_pack_taken & btb_117_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_117_bht_T_2 = btb_117_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_117_bht_T_3 = io_i_branch_resolve_pack_taken & btb_117_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_117_bht_T_4 = btb_117_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_117_bht_T_5 = io_i_branch_resolve_pack_taken & btb_117_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_117_bht_T_6 = btb_117_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_117_bht_T_7 = io_i_branch_resolve_pack_taken & btb_117_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_117_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_117_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_117_bht_T_13 = _btb_0_bht_T_8 & _btb_117_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_117_bht_T_16 = _btb_0_bht_T_8 & _btb_117_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_117_bht_T_19 = _btb_0_bht_T_8 & _btb_117_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_117_bht_T_20 = _btb_117_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_21 = _btb_117_bht_T_16 ? 2'h0 : _btb_117_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_22 = _btb_117_bht_T_13 ? 2'h0 : _btb_117_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_23 = _btb_117_bht_T_10 ? 2'h0 : _btb_117_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_24 = _btb_117_bht_T_7 ? 2'h3 : _btb_117_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_25 = _btb_117_bht_T_5 ? 2'h3 : _btb_117_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_26 = _btb_117_bht_T_3 ? 2'h3 : _btb_117_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_117_bht_T_27 = _btb_117_bht_T_1 ? 2'h1 : _btb_117_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9174 = btb_117_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6773
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9176 = btb_117_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_117_bht_T_27 : _GEN_8309; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_118_bht_T = btb_118_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_118_bht_T_1 = io_i_branch_resolve_pack_taken & btb_118_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_118_bht_T_2 = btb_118_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_118_bht_T_3 = io_i_branch_resolve_pack_taken & btb_118_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_118_bht_T_4 = btb_118_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_118_bht_T_5 = io_i_branch_resolve_pack_taken & btb_118_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_118_bht_T_6 = btb_118_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_118_bht_T_7 = io_i_branch_resolve_pack_taken & btb_118_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_118_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_118_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_118_bht_T_13 = _btb_0_bht_T_8 & _btb_118_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_118_bht_T_16 = _btb_0_bht_T_8 & _btb_118_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_118_bht_T_19 = _btb_0_bht_T_8 & _btb_118_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_118_bht_T_20 = _btb_118_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_21 = _btb_118_bht_T_16 ? 2'h0 : _btb_118_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_22 = _btb_118_bht_T_13 ? 2'h0 : _btb_118_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_23 = _btb_118_bht_T_10 ? 2'h0 : _btb_118_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_24 = _btb_118_bht_T_7 ? 2'h3 : _btb_118_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_25 = _btb_118_bht_T_5 ? 2'h3 : _btb_118_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_26 = _btb_118_bht_T_3 ? 2'h3 : _btb_118_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_118_bht_T_27 = _btb_118_bht_T_1 ? 2'h1 : _btb_118_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9178 = btb_118_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6774
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9180 = btb_118_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_118_bht_T_27 : _GEN_8310; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_119_bht_T = btb_119_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_119_bht_T_1 = io_i_branch_resolve_pack_taken & btb_119_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_119_bht_T_2 = btb_119_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_119_bht_T_3 = io_i_branch_resolve_pack_taken & btb_119_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_119_bht_T_4 = btb_119_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_119_bht_T_5 = io_i_branch_resolve_pack_taken & btb_119_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_119_bht_T_6 = btb_119_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_119_bht_T_7 = io_i_branch_resolve_pack_taken & btb_119_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_119_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_119_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_119_bht_T_13 = _btb_0_bht_T_8 & _btb_119_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_119_bht_T_16 = _btb_0_bht_T_8 & _btb_119_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_119_bht_T_19 = _btb_0_bht_T_8 & _btb_119_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_119_bht_T_20 = _btb_119_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_21 = _btb_119_bht_T_16 ? 2'h0 : _btb_119_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_22 = _btb_119_bht_T_13 ? 2'h0 : _btb_119_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_23 = _btb_119_bht_T_10 ? 2'h0 : _btb_119_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_24 = _btb_119_bht_T_7 ? 2'h3 : _btb_119_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_25 = _btb_119_bht_T_5 ? 2'h3 : _btb_119_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_26 = _btb_119_bht_T_3 ? 2'h3 : _btb_119_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_119_bht_T_27 = _btb_119_bht_T_1 ? 2'h1 : _btb_119_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9181 = btb_119_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_118_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_117_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_116_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_115_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_114_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_113_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_112_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_111_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_110_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_109_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_108_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_107_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_106_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_105_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9121)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9182 = btb_119_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6775
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9184 = btb_119_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_119_bht_T_27 : _GEN_8311; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_120_bht_T = btb_120_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_120_bht_T_1 = io_i_branch_resolve_pack_taken & btb_120_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_120_bht_T_2 = btb_120_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_120_bht_T_3 = io_i_branch_resolve_pack_taken & btb_120_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_120_bht_T_4 = btb_120_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_120_bht_T_5 = io_i_branch_resolve_pack_taken & btb_120_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_120_bht_T_6 = btb_120_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_120_bht_T_7 = io_i_branch_resolve_pack_taken & btb_120_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_120_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_120_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_120_bht_T_13 = _btb_0_bht_T_8 & _btb_120_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_120_bht_T_16 = _btb_0_bht_T_8 & _btb_120_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_120_bht_T_19 = _btb_0_bht_T_8 & _btb_120_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_120_bht_T_20 = _btb_120_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_21 = _btb_120_bht_T_16 ? 2'h0 : _btb_120_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_22 = _btb_120_bht_T_13 ? 2'h0 : _btb_120_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_23 = _btb_120_bht_T_10 ? 2'h0 : _btb_120_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_24 = _btb_120_bht_T_7 ? 2'h3 : _btb_120_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_25 = _btb_120_bht_T_5 ? 2'h3 : _btb_120_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_26 = _btb_120_bht_T_3 ? 2'h3 : _btb_120_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_120_bht_T_27 = _btb_120_bht_T_1 ? 2'h1 : _btb_120_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9186 = btb_120_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6776
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9188 = btb_120_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_120_bht_T_27 : _GEN_8312; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_121_bht_T = btb_121_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_121_bht_T_1 = io_i_branch_resolve_pack_taken & btb_121_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_121_bht_T_2 = btb_121_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_121_bht_T_3 = io_i_branch_resolve_pack_taken & btb_121_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_121_bht_T_4 = btb_121_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_121_bht_T_5 = io_i_branch_resolve_pack_taken & btb_121_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_121_bht_T_6 = btb_121_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_121_bht_T_7 = io_i_branch_resolve_pack_taken & btb_121_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_121_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_121_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_121_bht_T_13 = _btb_0_bht_T_8 & _btb_121_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_121_bht_T_16 = _btb_0_bht_T_8 & _btb_121_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_121_bht_T_19 = _btb_0_bht_T_8 & _btb_121_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_121_bht_T_20 = _btb_121_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_21 = _btb_121_bht_T_16 ? 2'h0 : _btb_121_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_22 = _btb_121_bht_T_13 ? 2'h0 : _btb_121_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_23 = _btb_121_bht_T_10 ? 2'h0 : _btb_121_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_24 = _btb_121_bht_T_7 ? 2'h3 : _btb_121_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_25 = _btb_121_bht_T_5 ? 2'h3 : _btb_121_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_26 = _btb_121_bht_T_3 ? 2'h3 : _btb_121_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_121_bht_T_27 = _btb_121_bht_T_1 ? 2'h1 : _btb_121_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9190 = btb_121_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6777
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9192 = btb_121_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_121_bht_T_27 : _GEN_8313; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_122_bht_T = btb_122_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_122_bht_T_1 = io_i_branch_resolve_pack_taken & btb_122_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_122_bht_T_2 = btb_122_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_122_bht_T_3 = io_i_branch_resolve_pack_taken & btb_122_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_122_bht_T_4 = btb_122_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_122_bht_T_5 = io_i_branch_resolve_pack_taken & btb_122_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_122_bht_T_6 = btb_122_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_122_bht_T_7 = io_i_branch_resolve_pack_taken & btb_122_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_122_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_122_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_122_bht_T_13 = _btb_0_bht_T_8 & _btb_122_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_122_bht_T_16 = _btb_0_bht_T_8 & _btb_122_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_122_bht_T_19 = _btb_0_bht_T_8 & _btb_122_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_122_bht_T_20 = _btb_122_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_21 = _btb_122_bht_T_16 ? 2'h0 : _btb_122_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_22 = _btb_122_bht_T_13 ? 2'h0 : _btb_122_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_23 = _btb_122_bht_T_10 ? 2'h0 : _btb_122_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_24 = _btb_122_bht_T_7 ? 2'h3 : _btb_122_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_25 = _btb_122_bht_T_5 ? 2'h3 : _btb_122_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_26 = _btb_122_bht_T_3 ? 2'h3 : _btb_122_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_122_bht_T_27 = _btb_122_bht_T_1 ? 2'h1 : _btb_122_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9194 = btb_122_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6778
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9196 = btb_122_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_122_bht_T_27 : _GEN_8314; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_123_bht_T = btb_123_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_123_bht_T_1 = io_i_branch_resolve_pack_taken & btb_123_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_123_bht_T_2 = btb_123_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_123_bht_T_3 = io_i_branch_resolve_pack_taken & btb_123_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_123_bht_T_4 = btb_123_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_123_bht_T_5 = io_i_branch_resolve_pack_taken & btb_123_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_123_bht_T_6 = btb_123_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_123_bht_T_7 = io_i_branch_resolve_pack_taken & btb_123_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_123_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_123_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_123_bht_T_13 = _btb_0_bht_T_8 & _btb_123_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_123_bht_T_16 = _btb_0_bht_T_8 & _btb_123_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_123_bht_T_19 = _btb_0_bht_T_8 & _btb_123_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_123_bht_T_20 = _btb_123_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_21 = _btb_123_bht_T_16 ? 2'h0 : _btb_123_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_22 = _btb_123_bht_T_13 ? 2'h0 : _btb_123_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_23 = _btb_123_bht_T_10 ? 2'h0 : _btb_123_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_24 = _btb_123_bht_T_7 ? 2'h3 : _btb_123_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_25 = _btb_123_bht_T_5 ? 2'h3 : _btb_123_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_26 = _btb_123_bht_T_3 ? 2'h3 : _btb_123_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_123_bht_T_27 = _btb_123_bht_T_1 ? 2'h1 : _btb_123_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9198 = btb_123_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6779
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9200 = btb_123_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_123_bht_T_27 : _GEN_8315; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_124_bht_T = btb_124_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_124_bht_T_1 = io_i_branch_resolve_pack_taken & btb_124_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_124_bht_T_2 = btb_124_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_124_bht_T_3 = io_i_branch_resolve_pack_taken & btb_124_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_124_bht_T_4 = btb_124_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_124_bht_T_5 = io_i_branch_resolve_pack_taken & btb_124_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_124_bht_T_6 = btb_124_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_124_bht_T_7 = io_i_branch_resolve_pack_taken & btb_124_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_124_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_124_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_124_bht_T_13 = _btb_0_bht_T_8 & _btb_124_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_124_bht_T_16 = _btb_0_bht_T_8 & _btb_124_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_124_bht_T_19 = _btb_0_bht_T_8 & _btb_124_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_124_bht_T_20 = _btb_124_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_21 = _btb_124_bht_T_16 ? 2'h0 : _btb_124_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_22 = _btb_124_bht_T_13 ? 2'h0 : _btb_124_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_23 = _btb_124_bht_T_10 ? 2'h0 : _btb_124_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_24 = _btb_124_bht_T_7 ? 2'h3 : _btb_124_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_25 = _btb_124_bht_T_5 ? 2'h3 : _btb_124_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_26 = _btb_124_bht_T_3 ? 2'h3 : _btb_124_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_124_bht_T_27 = _btb_124_bht_T_1 ? 2'h1 : _btb_124_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9202 = btb_124_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6780
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9204 = btb_124_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_124_bht_T_27 : _GEN_8316; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_125_bht_T = btb_125_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_125_bht_T_1 = io_i_branch_resolve_pack_taken & btb_125_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_125_bht_T_2 = btb_125_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_125_bht_T_3 = io_i_branch_resolve_pack_taken & btb_125_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_125_bht_T_4 = btb_125_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_125_bht_T_5 = io_i_branch_resolve_pack_taken & btb_125_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_125_bht_T_6 = btb_125_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_125_bht_T_7 = io_i_branch_resolve_pack_taken & btb_125_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_125_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_125_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_125_bht_T_13 = _btb_0_bht_T_8 & _btb_125_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_125_bht_T_16 = _btb_0_bht_T_8 & _btb_125_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_125_bht_T_19 = _btb_0_bht_T_8 & _btb_125_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_125_bht_T_20 = _btb_125_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_21 = _btb_125_bht_T_16 ? 2'h0 : _btb_125_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_22 = _btb_125_bht_T_13 ? 2'h0 : _btb_125_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_23 = _btb_125_bht_T_10 ? 2'h0 : _btb_125_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_24 = _btb_125_bht_T_7 ? 2'h3 : _btb_125_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_25 = _btb_125_bht_T_5 ? 2'h3 : _btb_125_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_26 = _btb_125_bht_T_3 ? 2'h3 : _btb_125_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_125_bht_T_27 = _btb_125_bht_T_1 ? 2'h1 : _btb_125_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9206 = btb_125_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6781
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9208 = btb_125_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_125_bht_T_27 : _GEN_8317; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_126_bht_T = btb_126_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_126_bht_T_1 = io_i_branch_resolve_pack_taken & btb_126_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_126_bht_T_2 = btb_126_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_126_bht_T_3 = io_i_branch_resolve_pack_taken & btb_126_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_126_bht_T_4 = btb_126_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_126_bht_T_5 = io_i_branch_resolve_pack_taken & btb_126_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_126_bht_T_6 = btb_126_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_126_bht_T_7 = io_i_branch_resolve_pack_taken & btb_126_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_126_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_126_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_126_bht_T_13 = _btb_0_bht_T_8 & _btb_126_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_126_bht_T_16 = _btb_0_bht_T_8 & _btb_126_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_126_bht_T_19 = _btb_0_bht_T_8 & _btb_126_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_126_bht_T_20 = _btb_126_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_21 = _btb_126_bht_T_16 ? 2'h0 : _btb_126_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_22 = _btb_126_bht_T_13 ? 2'h0 : _btb_126_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_23 = _btb_126_bht_T_10 ? 2'h0 : _btb_126_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_24 = _btb_126_bht_T_7 ? 2'h3 : _btb_126_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_25 = _btb_126_bht_T_5 ? 2'h3 : _btb_126_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_26 = _btb_126_bht_T_3 ? 2'h3 : _btb_126_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_126_bht_T_27 = _btb_126_bht_T_1 ? 2'h1 : _btb_126_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9210 = btb_126_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6782
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9212 = btb_126_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_126_bht_T_27 : _GEN_8318; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_127_bht_T = btb_127_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_127_bht_T_1 = io_i_branch_resolve_pack_taken & btb_127_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_127_bht_T_2 = btb_127_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_127_bht_T_3 = io_i_branch_resolve_pack_taken & btb_127_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_127_bht_T_4 = btb_127_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_127_bht_T_5 = io_i_branch_resolve_pack_taken & btb_127_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_127_bht_T_6 = btb_127_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_127_bht_T_7 = io_i_branch_resolve_pack_taken & btb_127_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_127_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_127_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_127_bht_T_13 = _btb_0_bht_T_8 & _btb_127_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_127_bht_T_16 = _btb_0_bht_T_8 & _btb_127_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_127_bht_T_19 = _btb_0_bht_T_8 & _btb_127_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_127_bht_T_20 = _btb_127_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_21 = _btb_127_bht_T_16 ? 2'h0 : _btb_127_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_22 = _btb_127_bht_T_13 ? 2'h0 : _btb_127_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_23 = _btb_127_bht_T_10 ? 2'h0 : _btb_127_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_24 = _btb_127_bht_T_7 ? 2'h3 : _btb_127_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_25 = _btb_127_bht_T_5 ? 2'h3 : _btb_127_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_26 = _btb_127_bht_T_3 ? 2'h3 : _btb_127_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_127_bht_T_27 = _btb_127_bht_T_1 ? 2'h1 : _btb_127_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9214 = btb_127_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6783
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9216 = btb_127_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_127_bht_T_27 : _GEN_8319; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_128_bht_T = btb_128_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_128_bht_T_1 = io_i_branch_resolve_pack_taken & btb_128_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_128_bht_T_2 = btb_128_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_128_bht_T_3 = io_i_branch_resolve_pack_taken & btb_128_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_128_bht_T_4 = btb_128_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_128_bht_T_5 = io_i_branch_resolve_pack_taken & btb_128_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_128_bht_T_6 = btb_128_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_128_bht_T_7 = io_i_branch_resolve_pack_taken & btb_128_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_128_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_128_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_128_bht_T_13 = _btb_0_bht_T_8 & _btb_128_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_128_bht_T_16 = _btb_0_bht_T_8 & _btb_128_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_128_bht_T_19 = _btb_0_bht_T_8 & _btb_128_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_128_bht_T_20 = _btb_128_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_21 = _btb_128_bht_T_16 ? 2'h0 : _btb_128_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_22 = _btb_128_bht_T_13 ? 2'h0 : _btb_128_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_23 = _btb_128_bht_T_10 ? 2'h0 : _btb_128_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_24 = _btb_128_bht_T_7 ? 2'h3 : _btb_128_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_25 = _btb_128_bht_T_5 ? 2'h3 : _btb_128_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_26 = _btb_128_bht_T_3 ? 2'h3 : _btb_128_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_128_bht_T_27 = _btb_128_bht_T_1 ? 2'h1 : _btb_128_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9218 = btb_128_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6784
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9220 = btb_128_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_128_bht_T_27 : _GEN_8320; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_129_bht_T = btb_129_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_129_bht_T_1 = io_i_branch_resolve_pack_taken & btb_129_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_129_bht_T_2 = btb_129_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_129_bht_T_3 = io_i_branch_resolve_pack_taken & btb_129_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_129_bht_T_4 = btb_129_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_129_bht_T_5 = io_i_branch_resolve_pack_taken & btb_129_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_129_bht_T_6 = btb_129_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_129_bht_T_7 = io_i_branch_resolve_pack_taken & btb_129_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_129_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_129_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_129_bht_T_13 = _btb_0_bht_T_8 & _btb_129_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_129_bht_T_16 = _btb_0_bht_T_8 & _btb_129_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_129_bht_T_19 = _btb_0_bht_T_8 & _btb_129_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_129_bht_T_20 = _btb_129_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_21 = _btb_129_bht_T_16 ? 2'h0 : _btb_129_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_22 = _btb_129_bht_T_13 ? 2'h0 : _btb_129_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_23 = _btb_129_bht_T_10 ? 2'h0 : _btb_129_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_24 = _btb_129_bht_T_7 ? 2'h3 : _btb_129_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_25 = _btb_129_bht_T_5 ? 2'h3 : _btb_129_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_26 = _btb_129_bht_T_3 ? 2'h3 : _btb_129_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_129_bht_T_27 = _btb_129_bht_T_1 ? 2'h1 : _btb_129_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9222 = btb_129_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6785
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9224 = btb_129_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_129_bht_T_27 : _GEN_8321; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_130_bht_T = btb_130_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_130_bht_T_1 = io_i_branch_resolve_pack_taken & btb_130_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_130_bht_T_2 = btb_130_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_130_bht_T_3 = io_i_branch_resolve_pack_taken & btb_130_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_130_bht_T_4 = btb_130_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_130_bht_T_5 = io_i_branch_resolve_pack_taken & btb_130_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_130_bht_T_6 = btb_130_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_130_bht_T_7 = io_i_branch_resolve_pack_taken & btb_130_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_130_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_130_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_130_bht_T_13 = _btb_0_bht_T_8 & _btb_130_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_130_bht_T_16 = _btb_0_bht_T_8 & _btb_130_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_130_bht_T_19 = _btb_0_bht_T_8 & _btb_130_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_130_bht_T_20 = _btb_130_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_21 = _btb_130_bht_T_16 ? 2'h0 : _btb_130_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_22 = _btb_130_bht_T_13 ? 2'h0 : _btb_130_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_23 = _btb_130_bht_T_10 ? 2'h0 : _btb_130_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_24 = _btb_130_bht_T_7 ? 2'h3 : _btb_130_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_25 = _btb_130_bht_T_5 ? 2'h3 : _btb_130_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_26 = _btb_130_bht_T_3 ? 2'h3 : _btb_130_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_130_bht_T_27 = _btb_130_bht_T_1 ? 2'h1 : _btb_130_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9226 = btb_130_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6786
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9228 = btb_130_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_130_bht_T_27 : _GEN_8322; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_131_bht_T = btb_131_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_131_bht_T_1 = io_i_branch_resolve_pack_taken & btb_131_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_131_bht_T_2 = btb_131_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_131_bht_T_3 = io_i_branch_resolve_pack_taken & btb_131_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_131_bht_T_4 = btb_131_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_131_bht_T_5 = io_i_branch_resolve_pack_taken & btb_131_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_131_bht_T_6 = btb_131_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_131_bht_T_7 = io_i_branch_resolve_pack_taken & btb_131_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_131_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_131_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_131_bht_T_13 = _btb_0_bht_T_8 & _btb_131_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_131_bht_T_16 = _btb_0_bht_T_8 & _btb_131_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_131_bht_T_19 = _btb_0_bht_T_8 & _btb_131_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_131_bht_T_20 = _btb_131_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_21 = _btb_131_bht_T_16 ? 2'h0 : _btb_131_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_22 = _btb_131_bht_T_13 ? 2'h0 : _btb_131_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_23 = _btb_131_bht_T_10 ? 2'h0 : _btb_131_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_24 = _btb_131_bht_T_7 ? 2'h3 : _btb_131_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_25 = _btb_131_bht_T_5 ? 2'h3 : _btb_131_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_26 = _btb_131_bht_T_3 ? 2'h3 : _btb_131_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_131_bht_T_27 = _btb_131_bht_T_1 ? 2'h1 : _btb_131_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9230 = btb_131_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6787
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9232 = btb_131_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_131_bht_T_27 : _GEN_8323; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_132_bht_T = btb_132_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_132_bht_T_1 = io_i_branch_resolve_pack_taken & btb_132_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_132_bht_T_2 = btb_132_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_132_bht_T_3 = io_i_branch_resolve_pack_taken & btb_132_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_132_bht_T_4 = btb_132_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_132_bht_T_5 = io_i_branch_resolve_pack_taken & btb_132_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_132_bht_T_6 = btb_132_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_132_bht_T_7 = io_i_branch_resolve_pack_taken & btb_132_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_132_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_132_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_132_bht_T_13 = _btb_0_bht_T_8 & _btb_132_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_132_bht_T_16 = _btb_0_bht_T_8 & _btb_132_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_132_bht_T_19 = _btb_0_bht_T_8 & _btb_132_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_132_bht_T_20 = _btb_132_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_21 = _btb_132_bht_T_16 ? 2'h0 : _btb_132_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_22 = _btb_132_bht_T_13 ? 2'h0 : _btb_132_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_23 = _btb_132_bht_T_10 ? 2'h0 : _btb_132_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_24 = _btb_132_bht_T_7 ? 2'h3 : _btb_132_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_25 = _btb_132_bht_T_5 ? 2'h3 : _btb_132_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_26 = _btb_132_bht_T_3 ? 2'h3 : _btb_132_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_132_bht_T_27 = _btb_132_bht_T_1 ? 2'h1 : _btb_132_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9234 = btb_132_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6788
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9236 = btb_132_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_132_bht_T_27 : _GEN_8324; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_133_bht_T = btb_133_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_133_bht_T_1 = io_i_branch_resolve_pack_taken & btb_133_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_133_bht_T_2 = btb_133_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_133_bht_T_3 = io_i_branch_resolve_pack_taken & btb_133_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_133_bht_T_4 = btb_133_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_133_bht_T_5 = io_i_branch_resolve_pack_taken & btb_133_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_133_bht_T_6 = btb_133_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_133_bht_T_7 = io_i_branch_resolve_pack_taken & btb_133_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_133_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_133_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_133_bht_T_13 = _btb_0_bht_T_8 & _btb_133_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_133_bht_T_16 = _btb_0_bht_T_8 & _btb_133_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_133_bht_T_19 = _btb_0_bht_T_8 & _btb_133_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_133_bht_T_20 = _btb_133_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_21 = _btb_133_bht_T_16 ? 2'h0 : _btb_133_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_22 = _btb_133_bht_T_13 ? 2'h0 : _btb_133_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_23 = _btb_133_bht_T_10 ? 2'h0 : _btb_133_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_24 = _btb_133_bht_T_7 ? 2'h3 : _btb_133_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_25 = _btb_133_bht_T_5 ? 2'h3 : _btb_133_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_26 = _btb_133_bht_T_3 ? 2'h3 : _btb_133_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_133_bht_T_27 = _btb_133_bht_T_1 ? 2'h1 : _btb_133_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9238 = btb_133_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6789
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9240 = btb_133_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_133_bht_T_27 : _GEN_8325; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_134_bht_T = btb_134_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_134_bht_T_1 = io_i_branch_resolve_pack_taken & btb_134_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_134_bht_T_2 = btb_134_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_134_bht_T_3 = io_i_branch_resolve_pack_taken & btb_134_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_134_bht_T_4 = btb_134_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_134_bht_T_5 = io_i_branch_resolve_pack_taken & btb_134_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_134_bht_T_6 = btb_134_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_134_bht_T_7 = io_i_branch_resolve_pack_taken & btb_134_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_134_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_134_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_134_bht_T_13 = _btb_0_bht_T_8 & _btb_134_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_134_bht_T_16 = _btb_0_bht_T_8 & _btb_134_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_134_bht_T_19 = _btb_0_bht_T_8 & _btb_134_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_134_bht_T_20 = _btb_134_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_21 = _btb_134_bht_T_16 ? 2'h0 : _btb_134_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_22 = _btb_134_bht_T_13 ? 2'h0 : _btb_134_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_23 = _btb_134_bht_T_10 ? 2'h0 : _btb_134_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_24 = _btb_134_bht_T_7 ? 2'h3 : _btb_134_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_25 = _btb_134_bht_T_5 ? 2'h3 : _btb_134_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_26 = _btb_134_bht_T_3 ? 2'h3 : _btb_134_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_134_bht_T_27 = _btb_134_bht_T_1 ? 2'h1 : _btb_134_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9241 = btb_134_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_133_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_132_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_131_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_130_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_129_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_128_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_127_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_126_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_125_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_124_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_123_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_122_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_121_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_120_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9181)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9242 = btb_134_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6790
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9244 = btb_134_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_134_bht_T_27 : _GEN_8326; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_135_bht_T = btb_135_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_135_bht_T_1 = io_i_branch_resolve_pack_taken & btb_135_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_135_bht_T_2 = btb_135_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_135_bht_T_3 = io_i_branch_resolve_pack_taken & btb_135_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_135_bht_T_4 = btb_135_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_135_bht_T_5 = io_i_branch_resolve_pack_taken & btb_135_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_135_bht_T_6 = btb_135_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_135_bht_T_7 = io_i_branch_resolve_pack_taken & btb_135_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_135_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_135_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_135_bht_T_13 = _btb_0_bht_T_8 & _btb_135_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_135_bht_T_16 = _btb_0_bht_T_8 & _btb_135_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_135_bht_T_19 = _btb_0_bht_T_8 & _btb_135_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_135_bht_T_20 = _btb_135_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_21 = _btb_135_bht_T_16 ? 2'h0 : _btb_135_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_22 = _btb_135_bht_T_13 ? 2'h0 : _btb_135_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_23 = _btb_135_bht_T_10 ? 2'h0 : _btb_135_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_24 = _btb_135_bht_T_7 ? 2'h3 : _btb_135_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_25 = _btb_135_bht_T_5 ? 2'h3 : _btb_135_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_26 = _btb_135_bht_T_3 ? 2'h3 : _btb_135_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_135_bht_T_27 = _btb_135_bht_T_1 ? 2'h1 : _btb_135_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9246 = btb_135_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6791
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9248 = btb_135_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_135_bht_T_27 : _GEN_8327; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_136_bht_T = btb_136_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_136_bht_T_1 = io_i_branch_resolve_pack_taken & btb_136_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_136_bht_T_2 = btb_136_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_136_bht_T_3 = io_i_branch_resolve_pack_taken & btb_136_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_136_bht_T_4 = btb_136_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_136_bht_T_5 = io_i_branch_resolve_pack_taken & btb_136_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_136_bht_T_6 = btb_136_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_136_bht_T_7 = io_i_branch_resolve_pack_taken & btb_136_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_136_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_136_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_136_bht_T_13 = _btb_0_bht_T_8 & _btb_136_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_136_bht_T_16 = _btb_0_bht_T_8 & _btb_136_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_136_bht_T_19 = _btb_0_bht_T_8 & _btb_136_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_136_bht_T_20 = _btb_136_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_21 = _btb_136_bht_T_16 ? 2'h0 : _btb_136_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_22 = _btb_136_bht_T_13 ? 2'h0 : _btb_136_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_23 = _btb_136_bht_T_10 ? 2'h0 : _btb_136_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_24 = _btb_136_bht_T_7 ? 2'h3 : _btb_136_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_25 = _btb_136_bht_T_5 ? 2'h3 : _btb_136_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_26 = _btb_136_bht_T_3 ? 2'h3 : _btb_136_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_136_bht_T_27 = _btb_136_bht_T_1 ? 2'h1 : _btb_136_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9250 = btb_136_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6792
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9252 = btb_136_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_136_bht_T_27 : _GEN_8328; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_137_bht_T = btb_137_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_137_bht_T_1 = io_i_branch_resolve_pack_taken & btb_137_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_137_bht_T_2 = btb_137_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_137_bht_T_3 = io_i_branch_resolve_pack_taken & btb_137_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_137_bht_T_4 = btb_137_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_137_bht_T_5 = io_i_branch_resolve_pack_taken & btb_137_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_137_bht_T_6 = btb_137_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_137_bht_T_7 = io_i_branch_resolve_pack_taken & btb_137_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_137_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_137_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_137_bht_T_13 = _btb_0_bht_T_8 & _btb_137_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_137_bht_T_16 = _btb_0_bht_T_8 & _btb_137_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_137_bht_T_19 = _btb_0_bht_T_8 & _btb_137_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_137_bht_T_20 = _btb_137_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_21 = _btb_137_bht_T_16 ? 2'h0 : _btb_137_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_22 = _btb_137_bht_T_13 ? 2'h0 : _btb_137_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_23 = _btb_137_bht_T_10 ? 2'h0 : _btb_137_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_24 = _btb_137_bht_T_7 ? 2'h3 : _btb_137_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_25 = _btb_137_bht_T_5 ? 2'h3 : _btb_137_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_26 = _btb_137_bht_T_3 ? 2'h3 : _btb_137_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_137_bht_T_27 = _btb_137_bht_T_1 ? 2'h1 : _btb_137_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9254 = btb_137_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6793
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9256 = btb_137_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_137_bht_T_27 : _GEN_8329; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_138_bht_T = btb_138_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_138_bht_T_1 = io_i_branch_resolve_pack_taken & btb_138_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_138_bht_T_2 = btb_138_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_138_bht_T_3 = io_i_branch_resolve_pack_taken & btb_138_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_138_bht_T_4 = btb_138_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_138_bht_T_5 = io_i_branch_resolve_pack_taken & btb_138_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_138_bht_T_6 = btb_138_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_138_bht_T_7 = io_i_branch_resolve_pack_taken & btb_138_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_138_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_138_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_138_bht_T_13 = _btb_0_bht_T_8 & _btb_138_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_138_bht_T_16 = _btb_0_bht_T_8 & _btb_138_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_138_bht_T_19 = _btb_0_bht_T_8 & _btb_138_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_138_bht_T_20 = _btb_138_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_21 = _btb_138_bht_T_16 ? 2'h0 : _btb_138_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_22 = _btb_138_bht_T_13 ? 2'h0 : _btb_138_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_23 = _btb_138_bht_T_10 ? 2'h0 : _btb_138_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_24 = _btb_138_bht_T_7 ? 2'h3 : _btb_138_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_25 = _btb_138_bht_T_5 ? 2'h3 : _btb_138_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_26 = _btb_138_bht_T_3 ? 2'h3 : _btb_138_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_138_bht_T_27 = _btb_138_bht_T_1 ? 2'h1 : _btb_138_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9258 = btb_138_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6794
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9260 = btb_138_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_138_bht_T_27 : _GEN_8330; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_139_bht_T = btb_139_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_139_bht_T_1 = io_i_branch_resolve_pack_taken & btb_139_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_139_bht_T_2 = btb_139_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_139_bht_T_3 = io_i_branch_resolve_pack_taken & btb_139_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_139_bht_T_4 = btb_139_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_139_bht_T_5 = io_i_branch_resolve_pack_taken & btb_139_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_139_bht_T_6 = btb_139_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_139_bht_T_7 = io_i_branch_resolve_pack_taken & btb_139_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_139_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_139_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_139_bht_T_13 = _btb_0_bht_T_8 & _btb_139_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_139_bht_T_16 = _btb_0_bht_T_8 & _btb_139_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_139_bht_T_19 = _btb_0_bht_T_8 & _btb_139_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_139_bht_T_20 = _btb_139_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_21 = _btb_139_bht_T_16 ? 2'h0 : _btb_139_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_22 = _btb_139_bht_T_13 ? 2'h0 : _btb_139_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_23 = _btb_139_bht_T_10 ? 2'h0 : _btb_139_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_24 = _btb_139_bht_T_7 ? 2'h3 : _btb_139_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_25 = _btb_139_bht_T_5 ? 2'h3 : _btb_139_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_26 = _btb_139_bht_T_3 ? 2'h3 : _btb_139_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_139_bht_T_27 = _btb_139_bht_T_1 ? 2'h1 : _btb_139_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9262 = btb_139_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6795
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9264 = btb_139_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_139_bht_T_27 : _GEN_8331; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_140_bht_T = btb_140_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_140_bht_T_1 = io_i_branch_resolve_pack_taken & btb_140_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_140_bht_T_2 = btb_140_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_140_bht_T_3 = io_i_branch_resolve_pack_taken & btb_140_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_140_bht_T_4 = btb_140_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_140_bht_T_5 = io_i_branch_resolve_pack_taken & btb_140_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_140_bht_T_6 = btb_140_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_140_bht_T_7 = io_i_branch_resolve_pack_taken & btb_140_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_140_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_140_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_140_bht_T_13 = _btb_0_bht_T_8 & _btb_140_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_140_bht_T_16 = _btb_0_bht_T_8 & _btb_140_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_140_bht_T_19 = _btb_0_bht_T_8 & _btb_140_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_140_bht_T_20 = _btb_140_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_21 = _btb_140_bht_T_16 ? 2'h0 : _btb_140_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_22 = _btb_140_bht_T_13 ? 2'h0 : _btb_140_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_23 = _btb_140_bht_T_10 ? 2'h0 : _btb_140_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_24 = _btb_140_bht_T_7 ? 2'h3 : _btb_140_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_25 = _btb_140_bht_T_5 ? 2'h3 : _btb_140_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_26 = _btb_140_bht_T_3 ? 2'h3 : _btb_140_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_140_bht_T_27 = _btb_140_bht_T_1 ? 2'h1 : _btb_140_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9266 = btb_140_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6796
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9268 = btb_140_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_140_bht_T_27 : _GEN_8332; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_141_bht_T = btb_141_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_141_bht_T_1 = io_i_branch_resolve_pack_taken & btb_141_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_141_bht_T_2 = btb_141_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_141_bht_T_3 = io_i_branch_resolve_pack_taken & btb_141_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_141_bht_T_4 = btb_141_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_141_bht_T_5 = io_i_branch_resolve_pack_taken & btb_141_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_141_bht_T_6 = btb_141_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_141_bht_T_7 = io_i_branch_resolve_pack_taken & btb_141_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_141_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_141_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_141_bht_T_13 = _btb_0_bht_T_8 & _btb_141_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_141_bht_T_16 = _btb_0_bht_T_8 & _btb_141_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_141_bht_T_19 = _btb_0_bht_T_8 & _btb_141_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_141_bht_T_20 = _btb_141_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_21 = _btb_141_bht_T_16 ? 2'h0 : _btb_141_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_22 = _btb_141_bht_T_13 ? 2'h0 : _btb_141_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_23 = _btb_141_bht_T_10 ? 2'h0 : _btb_141_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_24 = _btb_141_bht_T_7 ? 2'h3 : _btb_141_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_25 = _btb_141_bht_T_5 ? 2'h3 : _btb_141_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_26 = _btb_141_bht_T_3 ? 2'h3 : _btb_141_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_141_bht_T_27 = _btb_141_bht_T_1 ? 2'h1 : _btb_141_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9270 = btb_141_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6797
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9272 = btb_141_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_141_bht_T_27 : _GEN_8333; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_142_bht_T = btb_142_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_142_bht_T_1 = io_i_branch_resolve_pack_taken & btb_142_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_142_bht_T_2 = btb_142_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_142_bht_T_3 = io_i_branch_resolve_pack_taken & btb_142_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_142_bht_T_4 = btb_142_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_142_bht_T_5 = io_i_branch_resolve_pack_taken & btb_142_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_142_bht_T_6 = btb_142_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_142_bht_T_7 = io_i_branch_resolve_pack_taken & btb_142_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_142_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_142_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_142_bht_T_13 = _btb_0_bht_T_8 & _btb_142_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_142_bht_T_16 = _btb_0_bht_T_8 & _btb_142_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_142_bht_T_19 = _btb_0_bht_T_8 & _btb_142_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_142_bht_T_20 = _btb_142_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_21 = _btb_142_bht_T_16 ? 2'h0 : _btb_142_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_22 = _btb_142_bht_T_13 ? 2'h0 : _btb_142_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_23 = _btb_142_bht_T_10 ? 2'h0 : _btb_142_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_24 = _btb_142_bht_T_7 ? 2'h3 : _btb_142_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_25 = _btb_142_bht_T_5 ? 2'h3 : _btb_142_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_26 = _btb_142_bht_T_3 ? 2'h3 : _btb_142_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_142_bht_T_27 = _btb_142_bht_T_1 ? 2'h1 : _btb_142_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9274 = btb_142_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6798
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9276 = btb_142_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_142_bht_T_27 : _GEN_8334; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_143_bht_T = btb_143_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_143_bht_T_1 = io_i_branch_resolve_pack_taken & btb_143_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_143_bht_T_2 = btb_143_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_143_bht_T_3 = io_i_branch_resolve_pack_taken & btb_143_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_143_bht_T_4 = btb_143_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_143_bht_T_5 = io_i_branch_resolve_pack_taken & btb_143_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_143_bht_T_6 = btb_143_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_143_bht_T_7 = io_i_branch_resolve_pack_taken & btb_143_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_143_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_143_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_143_bht_T_13 = _btb_0_bht_T_8 & _btb_143_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_143_bht_T_16 = _btb_0_bht_T_8 & _btb_143_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_143_bht_T_19 = _btb_0_bht_T_8 & _btb_143_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_143_bht_T_20 = _btb_143_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_21 = _btb_143_bht_T_16 ? 2'h0 : _btb_143_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_22 = _btb_143_bht_T_13 ? 2'h0 : _btb_143_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_23 = _btb_143_bht_T_10 ? 2'h0 : _btb_143_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_24 = _btb_143_bht_T_7 ? 2'h3 : _btb_143_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_25 = _btb_143_bht_T_5 ? 2'h3 : _btb_143_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_26 = _btb_143_bht_T_3 ? 2'h3 : _btb_143_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_143_bht_T_27 = _btb_143_bht_T_1 ? 2'h1 : _btb_143_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9278 = btb_143_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6799
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9280 = btb_143_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_143_bht_T_27 : _GEN_8335; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_144_bht_T = btb_144_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_144_bht_T_1 = io_i_branch_resolve_pack_taken & btb_144_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_144_bht_T_2 = btb_144_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_144_bht_T_3 = io_i_branch_resolve_pack_taken & btb_144_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_144_bht_T_4 = btb_144_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_144_bht_T_5 = io_i_branch_resolve_pack_taken & btb_144_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_144_bht_T_6 = btb_144_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_144_bht_T_7 = io_i_branch_resolve_pack_taken & btb_144_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_144_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_144_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_144_bht_T_13 = _btb_0_bht_T_8 & _btb_144_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_144_bht_T_16 = _btb_0_bht_T_8 & _btb_144_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_144_bht_T_19 = _btb_0_bht_T_8 & _btb_144_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_144_bht_T_20 = _btb_144_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_21 = _btb_144_bht_T_16 ? 2'h0 : _btb_144_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_22 = _btb_144_bht_T_13 ? 2'h0 : _btb_144_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_23 = _btb_144_bht_T_10 ? 2'h0 : _btb_144_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_24 = _btb_144_bht_T_7 ? 2'h3 : _btb_144_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_25 = _btb_144_bht_T_5 ? 2'h3 : _btb_144_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_26 = _btb_144_bht_T_3 ? 2'h3 : _btb_144_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_144_bht_T_27 = _btb_144_bht_T_1 ? 2'h1 : _btb_144_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9282 = btb_144_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6800
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9284 = btb_144_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_144_bht_T_27 : _GEN_8336; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_145_bht_T = btb_145_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_145_bht_T_1 = io_i_branch_resolve_pack_taken & btb_145_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_145_bht_T_2 = btb_145_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_145_bht_T_3 = io_i_branch_resolve_pack_taken & btb_145_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_145_bht_T_4 = btb_145_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_145_bht_T_5 = io_i_branch_resolve_pack_taken & btb_145_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_145_bht_T_6 = btb_145_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_145_bht_T_7 = io_i_branch_resolve_pack_taken & btb_145_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_145_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_145_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_145_bht_T_13 = _btb_0_bht_T_8 & _btb_145_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_145_bht_T_16 = _btb_0_bht_T_8 & _btb_145_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_145_bht_T_19 = _btb_0_bht_T_8 & _btb_145_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_145_bht_T_20 = _btb_145_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_21 = _btb_145_bht_T_16 ? 2'h0 : _btb_145_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_22 = _btb_145_bht_T_13 ? 2'h0 : _btb_145_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_23 = _btb_145_bht_T_10 ? 2'h0 : _btb_145_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_24 = _btb_145_bht_T_7 ? 2'h3 : _btb_145_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_25 = _btb_145_bht_T_5 ? 2'h3 : _btb_145_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_26 = _btb_145_bht_T_3 ? 2'h3 : _btb_145_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_145_bht_T_27 = _btb_145_bht_T_1 ? 2'h1 : _btb_145_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9286 = btb_145_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6801
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9288 = btb_145_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_145_bht_T_27 : _GEN_8337; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_146_bht_T = btb_146_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_146_bht_T_1 = io_i_branch_resolve_pack_taken & btb_146_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_146_bht_T_2 = btb_146_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_146_bht_T_3 = io_i_branch_resolve_pack_taken & btb_146_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_146_bht_T_4 = btb_146_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_146_bht_T_5 = io_i_branch_resolve_pack_taken & btb_146_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_146_bht_T_6 = btb_146_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_146_bht_T_7 = io_i_branch_resolve_pack_taken & btb_146_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_146_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_146_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_146_bht_T_13 = _btb_0_bht_T_8 & _btb_146_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_146_bht_T_16 = _btb_0_bht_T_8 & _btb_146_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_146_bht_T_19 = _btb_0_bht_T_8 & _btb_146_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_146_bht_T_20 = _btb_146_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_21 = _btb_146_bht_T_16 ? 2'h0 : _btb_146_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_22 = _btb_146_bht_T_13 ? 2'h0 : _btb_146_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_23 = _btb_146_bht_T_10 ? 2'h0 : _btb_146_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_24 = _btb_146_bht_T_7 ? 2'h3 : _btb_146_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_25 = _btb_146_bht_T_5 ? 2'h3 : _btb_146_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_26 = _btb_146_bht_T_3 ? 2'h3 : _btb_146_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_146_bht_T_27 = _btb_146_bht_T_1 ? 2'h1 : _btb_146_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9290 = btb_146_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6802
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9292 = btb_146_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_146_bht_T_27 : _GEN_8338; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_147_bht_T = btb_147_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_147_bht_T_1 = io_i_branch_resolve_pack_taken & btb_147_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_147_bht_T_2 = btb_147_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_147_bht_T_3 = io_i_branch_resolve_pack_taken & btb_147_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_147_bht_T_4 = btb_147_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_147_bht_T_5 = io_i_branch_resolve_pack_taken & btb_147_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_147_bht_T_6 = btb_147_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_147_bht_T_7 = io_i_branch_resolve_pack_taken & btb_147_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_147_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_147_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_147_bht_T_13 = _btb_0_bht_T_8 & _btb_147_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_147_bht_T_16 = _btb_0_bht_T_8 & _btb_147_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_147_bht_T_19 = _btb_0_bht_T_8 & _btb_147_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_147_bht_T_20 = _btb_147_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_21 = _btb_147_bht_T_16 ? 2'h0 : _btb_147_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_22 = _btb_147_bht_T_13 ? 2'h0 : _btb_147_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_23 = _btb_147_bht_T_10 ? 2'h0 : _btb_147_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_24 = _btb_147_bht_T_7 ? 2'h3 : _btb_147_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_25 = _btb_147_bht_T_5 ? 2'h3 : _btb_147_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_26 = _btb_147_bht_T_3 ? 2'h3 : _btb_147_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_147_bht_T_27 = _btb_147_bht_T_1 ? 2'h1 : _btb_147_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9294 = btb_147_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6803
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9296 = btb_147_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_147_bht_T_27 : _GEN_8339; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_148_bht_T = btb_148_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_148_bht_T_1 = io_i_branch_resolve_pack_taken & btb_148_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_148_bht_T_2 = btb_148_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_148_bht_T_3 = io_i_branch_resolve_pack_taken & btb_148_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_148_bht_T_4 = btb_148_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_148_bht_T_5 = io_i_branch_resolve_pack_taken & btb_148_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_148_bht_T_6 = btb_148_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_148_bht_T_7 = io_i_branch_resolve_pack_taken & btb_148_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_148_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_148_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_148_bht_T_13 = _btb_0_bht_T_8 & _btb_148_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_148_bht_T_16 = _btb_0_bht_T_8 & _btb_148_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_148_bht_T_19 = _btb_0_bht_T_8 & _btb_148_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_148_bht_T_20 = _btb_148_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_21 = _btb_148_bht_T_16 ? 2'h0 : _btb_148_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_22 = _btb_148_bht_T_13 ? 2'h0 : _btb_148_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_23 = _btb_148_bht_T_10 ? 2'h0 : _btb_148_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_24 = _btb_148_bht_T_7 ? 2'h3 : _btb_148_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_25 = _btb_148_bht_T_5 ? 2'h3 : _btb_148_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_26 = _btb_148_bht_T_3 ? 2'h3 : _btb_148_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_148_bht_T_27 = _btb_148_bht_T_1 ? 2'h1 : _btb_148_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9298 = btb_148_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6804
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9300 = btb_148_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_148_bht_T_27 : _GEN_8340; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_149_bht_T = btb_149_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_149_bht_T_1 = io_i_branch_resolve_pack_taken & btb_149_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_149_bht_T_2 = btb_149_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_149_bht_T_3 = io_i_branch_resolve_pack_taken & btb_149_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_149_bht_T_4 = btb_149_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_149_bht_T_5 = io_i_branch_resolve_pack_taken & btb_149_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_149_bht_T_6 = btb_149_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_149_bht_T_7 = io_i_branch_resolve_pack_taken & btb_149_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_149_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_149_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_149_bht_T_13 = _btb_0_bht_T_8 & _btb_149_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_149_bht_T_16 = _btb_0_bht_T_8 & _btb_149_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_149_bht_T_19 = _btb_0_bht_T_8 & _btb_149_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_149_bht_T_20 = _btb_149_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_21 = _btb_149_bht_T_16 ? 2'h0 : _btb_149_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_22 = _btb_149_bht_T_13 ? 2'h0 : _btb_149_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_23 = _btb_149_bht_T_10 ? 2'h0 : _btb_149_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_24 = _btb_149_bht_T_7 ? 2'h3 : _btb_149_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_25 = _btb_149_bht_T_5 ? 2'h3 : _btb_149_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_26 = _btb_149_bht_T_3 ? 2'h3 : _btb_149_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_149_bht_T_27 = _btb_149_bht_T_1 ? 2'h1 : _btb_149_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9301 = btb_149_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_148_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_147_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_146_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_145_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_144_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_143_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_142_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_141_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_140_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_139_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_138_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_137_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_136_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_135_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9241)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9302 = btb_149_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6805
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9304 = btb_149_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_149_bht_T_27 : _GEN_8341; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_150_bht_T = btb_150_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_150_bht_T_1 = io_i_branch_resolve_pack_taken & btb_150_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_150_bht_T_2 = btb_150_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_150_bht_T_3 = io_i_branch_resolve_pack_taken & btb_150_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_150_bht_T_4 = btb_150_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_150_bht_T_5 = io_i_branch_resolve_pack_taken & btb_150_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_150_bht_T_6 = btb_150_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_150_bht_T_7 = io_i_branch_resolve_pack_taken & btb_150_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_150_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_150_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_150_bht_T_13 = _btb_0_bht_T_8 & _btb_150_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_150_bht_T_16 = _btb_0_bht_T_8 & _btb_150_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_150_bht_T_19 = _btb_0_bht_T_8 & _btb_150_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_150_bht_T_20 = _btb_150_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_21 = _btb_150_bht_T_16 ? 2'h0 : _btb_150_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_22 = _btb_150_bht_T_13 ? 2'h0 : _btb_150_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_23 = _btb_150_bht_T_10 ? 2'h0 : _btb_150_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_24 = _btb_150_bht_T_7 ? 2'h3 : _btb_150_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_25 = _btb_150_bht_T_5 ? 2'h3 : _btb_150_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_26 = _btb_150_bht_T_3 ? 2'h3 : _btb_150_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_150_bht_T_27 = _btb_150_bht_T_1 ? 2'h1 : _btb_150_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9306 = btb_150_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6806
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9308 = btb_150_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_150_bht_T_27 : _GEN_8342; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_151_bht_T = btb_151_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_151_bht_T_1 = io_i_branch_resolve_pack_taken & btb_151_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_151_bht_T_2 = btb_151_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_151_bht_T_3 = io_i_branch_resolve_pack_taken & btb_151_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_151_bht_T_4 = btb_151_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_151_bht_T_5 = io_i_branch_resolve_pack_taken & btb_151_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_151_bht_T_6 = btb_151_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_151_bht_T_7 = io_i_branch_resolve_pack_taken & btb_151_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_151_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_151_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_151_bht_T_13 = _btb_0_bht_T_8 & _btb_151_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_151_bht_T_16 = _btb_0_bht_T_8 & _btb_151_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_151_bht_T_19 = _btb_0_bht_T_8 & _btb_151_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_151_bht_T_20 = _btb_151_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_21 = _btb_151_bht_T_16 ? 2'h0 : _btb_151_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_22 = _btb_151_bht_T_13 ? 2'h0 : _btb_151_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_23 = _btb_151_bht_T_10 ? 2'h0 : _btb_151_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_24 = _btb_151_bht_T_7 ? 2'h3 : _btb_151_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_25 = _btb_151_bht_T_5 ? 2'h3 : _btb_151_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_26 = _btb_151_bht_T_3 ? 2'h3 : _btb_151_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_151_bht_T_27 = _btb_151_bht_T_1 ? 2'h1 : _btb_151_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9310 = btb_151_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6807
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9312 = btb_151_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_151_bht_T_27 : _GEN_8343; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_152_bht_T = btb_152_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_152_bht_T_1 = io_i_branch_resolve_pack_taken & btb_152_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_152_bht_T_2 = btb_152_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_152_bht_T_3 = io_i_branch_resolve_pack_taken & btb_152_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_152_bht_T_4 = btb_152_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_152_bht_T_5 = io_i_branch_resolve_pack_taken & btb_152_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_152_bht_T_6 = btb_152_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_152_bht_T_7 = io_i_branch_resolve_pack_taken & btb_152_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_152_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_152_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_152_bht_T_13 = _btb_0_bht_T_8 & _btb_152_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_152_bht_T_16 = _btb_0_bht_T_8 & _btb_152_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_152_bht_T_19 = _btb_0_bht_T_8 & _btb_152_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_152_bht_T_20 = _btb_152_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_21 = _btb_152_bht_T_16 ? 2'h0 : _btb_152_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_22 = _btb_152_bht_T_13 ? 2'h0 : _btb_152_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_23 = _btb_152_bht_T_10 ? 2'h0 : _btb_152_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_24 = _btb_152_bht_T_7 ? 2'h3 : _btb_152_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_25 = _btb_152_bht_T_5 ? 2'h3 : _btb_152_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_26 = _btb_152_bht_T_3 ? 2'h3 : _btb_152_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_152_bht_T_27 = _btb_152_bht_T_1 ? 2'h1 : _btb_152_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9314 = btb_152_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6808
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9316 = btb_152_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_152_bht_T_27 : _GEN_8344; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_153_bht_T = btb_153_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_153_bht_T_1 = io_i_branch_resolve_pack_taken & btb_153_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_153_bht_T_2 = btb_153_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_153_bht_T_3 = io_i_branch_resolve_pack_taken & btb_153_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_153_bht_T_4 = btb_153_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_153_bht_T_5 = io_i_branch_resolve_pack_taken & btb_153_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_153_bht_T_6 = btb_153_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_153_bht_T_7 = io_i_branch_resolve_pack_taken & btb_153_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_153_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_153_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_153_bht_T_13 = _btb_0_bht_T_8 & _btb_153_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_153_bht_T_16 = _btb_0_bht_T_8 & _btb_153_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_153_bht_T_19 = _btb_0_bht_T_8 & _btb_153_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_153_bht_T_20 = _btb_153_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_21 = _btb_153_bht_T_16 ? 2'h0 : _btb_153_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_22 = _btb_153_bht_T_13 ? 2'h0 : _btb_153_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_23 = _btb_153_bht_T_10 ? 2'h0 : _btb_153_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_24 = _btb_153_bht_T_7 ? 2'h3 : _btb_153_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_25 = _btb_153_bht_T_5 ? 2'h3 : _btb_153_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_26 = _btb_153_bht_T_3 ? 2'h3 : _btb_153_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_153_bht_T_27 = _btb_153_bht_T_1 ? 2'h1 : _btb_153_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9318 = btb_153_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6809
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9320 = btb_153_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_153_bht_T_27 : _GEN_8345; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_154_bht_T = btb_154_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_154_bht_T_1 = io_i_branch_resolve_pack_taken & btb_154_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_154_bht_T_2 = btb_154_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_154_bht_T_3 = io_i_branch_resolve_pack_taken & btb_154_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_154_bht_T_4 = btb_154_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_154_bht_T_5 = io_i_branch_resolve_pack_taken & btb_154_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_154_bht_T_6 = btb_154_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_154_bht_T_7 = io_i_branch_resolve_pack_taken & btb_154_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_154_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_154_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_154_bht_T_13 = _btb_0_bht_T_8 & _btb_154_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_154_bht_T_16 = _btb_0_bht_T_8 & _btb_154_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_154_bht_T_19 = _btb_0_bht_T_8 & _btb_154_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_154_bht_T_20 = _btb_154_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_21 = _btb_154_bht_T_16 ? 2'h0 : _btb_154_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_22 = _btb_154_bht_T_13 ? 2'h0 : _btb_154_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_23 = _btb_154_bht_T_10 ? 2'h0 : _btb_154_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_24 = _btb_154_bht_T_7 ? 2'h3 : _btb_154_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_25 = _btb_154_bht_T_5 ? 2'h3 : _btb_154_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_26 = _btb_154_bht_T_3 ? 2'h3 : _btb_154_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_154_bht_T_27 = _btb_154_bht_T_1 ? 2'h1 : _btb_154_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9322 = btb_154_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6810
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9324 = btb_154_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_154_bht_T_27 : _GEN_8346; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_155_bht_T = btb_155_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_155_bht_T_1 = io_i_branch_resolve_pack_taken & btb_155_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_155_bht_T_2 = btb_155_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_155_bht_T_3 = io_i_branch_resolve_pack_taken & btb_155_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_155_bht_T_4 = btb_155_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_155_bht_T_5 = io_i_branch_resolve_pack_taken & btb_155_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_155_bht_T_6 = btb_155_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_155_bht_T_7 = io_i_branch_resolve_pack_taken & btb_155_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_155_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_155_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_155_bht_T_13 = _btb_0_bht_T_8 & _btb_155_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_155_bht_T_16 = _btb_0_bht_T_8 & _btb_155_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_155_bht_T_19 = _btb_0_bht_T_8 & _btb_155_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_155_bht_T_20 = _btb_155_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_21 = _btb_155_bht_T_16 ? 2'h0 : _btb_155_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_22 = _btb_155_bht_T_13 ? 2'h0 : _btb_155_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_23 = _btb_155_bht_T_10 ? 2'h0 : _btb_155_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_24 = _btb_155_bht_T_7 ? 2'h3 : _btb_155_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_25 = _btb_155_bht_T_5 ? 2'h3 : _btb_155_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_26 = _btb_155_bht_T_3 ? 2'h3 : _btb_155_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_155_bht_T_27 = _btb_155_bht_T_1 ? 2'h1 : _btb_155_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9326 = btb_155_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6811
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9328 = btb_155_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_155_bht_T_27 : _GEN_8347; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_156_bht_T = btb_156_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_156_bht_T_1 = io_i_branch_resolve_pack_taken & btb_156_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_156_bht_T_2 = btb_156_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_156_bht_T_3 = io_i_branch_resolve_pack_taken & btb_156_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_156_bht_T_4 = btb_156_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_156_bht_T_5 = io_i_branch_resolve_pack_taken & btb_156_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_156_bht_T_6 = btb_156_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_156_bht_T_7 = io_i_branch_resolve_pack_taken & btb_156_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_156_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_156_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_156_bht_T_13 = _btb_0_bht_T_8 & _btb_156_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_156_bht_T_16 = _btb_0_bht_T_8 & _btb_156_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_156_bht_T_19 = _btb_0_bht_T_8 & _btb_156_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_156_bht_T_20 = _btb_156_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_21 = _btb_156_bht_T_16 ? 2'h0 : _btb_156_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_22 = _btb_156_bht_T_13 ? 2'h0 : _btb_156_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_23 = _btb_156_bht_T_10 ? 2'h0 : _btb_156_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_24 = _btb_156_bht_T_7 ? 2'h3 : _btb_156_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_25 = _btb_156_bht_T_5 ? 2'h3 : _btb_156_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_26 = _btb_156_bht_T_3 ? 2'h3 : _btb_156_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_156_bht_T_27 = _btb_156_bht_T_1 ? 2'h1 : _btb_156_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9330 = btb_156_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6812
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9332 = btb_156_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_156_bht_T_27 : _GEN_8348; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_157_bht_T = btb_157_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_157_bht_T_1 = io_i_branch_resolve_pack_taken & btb_157_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_157_bht_T_2 = btb_157_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_157_bht_T_3 = io_i_branch_resolve_pack_taken & btb_157_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_157_bht_T_4 = btb_157_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_157_bht_T_5 = io_i_branch_resolve_pack_taken & btb_157_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_157_bht_T_6 = btb_157_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_157_bht_T_7 = io_i_branch_resolve_pack_taken & btb_157_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_157_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_157_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_157_bht_T_13 = _btb_0_bht_T_8 & _btb_157_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_157_bht_T_16 = _btb_0_bht_T_8 & _btb_157_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_157_bht_T_19 = _btb_0_bht_T_8 & _btb_157_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_157_bht_T_20 = _btb_157_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_21 = _btb_157_bht_T_16 ? 2'h0 : _btb_157_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_22 = _btb_157_bht_T_13 ? 2'h0 : _btb_157_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_23 = _btb_157_bht_T_10 ? 2'h0 : _btb_157_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_24 = _btb_157_bht_T_7 ? 2'h3 : _btb_157_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_25 = _btb_157_bht_T_5 ? 2'h3 : _btb_157_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_26 = _btb_157_bht_T_3 ? 2'h3 : _btb_157_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_157_bht_T_27 = _btb_157_bht_T_1 ? 2'h1 : _btb_157_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9334 = btb_157_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6813
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9336 = btb_157_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_157_bht_T_27 : _GEN_8349; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_158_bht_T = btb_158_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_158_bht_T_1 = io_i_branch_resolve_pack_taken & btb_158_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_158_bht_T_2 = btb_158_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_158_bht_T_3 = io_i_branch_resolve_pack_taken & btb_158_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_158_bht_T_4 = btb_158_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_158_bht_T_5 = io_i_branch_resolve_pack_taken & btb_158_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_158_bht_T_6 = btb_158_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_158_bht_T_7 = io_i_branch_resolve_pack_taken & btb_158_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_158_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_158_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_158_bht_T_13 = _btb_0_bht_T_8 & _btb_158_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_158_bht_T_16 = _btb_0_bht_T_8 & _btb_158_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_158_bht_T_19 = _btb_0_bht_T_8 & _btb_158_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_158_bht_T_20 = _btb_158_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_21 = _btb_158_bht_T_16 ? 2'h0 : _btb_158_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_22 = _btb_158_bht_T_13 ? 2'h0 : _btb_158_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_23 = _btb_158_bht_T_10 ? 2'h0 : _btb_158_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_24 = _btb_158_bht_T_7 ? 2'h3 : _btb_158_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_25 = _btb_158_bht_T_5 ? 2'h3 : _btb_158_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_26 = _btb_158_bht_T_3 ? 2'h3 : _btb_158_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_158_bht_T_27 = _btb_158_bht_T_1 ? 2'h1 : _btb_158_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9338 = btb_158_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6814
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9340 = btb_158_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_158_bht_T_27 : _GEN_8350; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_159_bht_T = btb_159_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_159_bht_T_1 = io_i_branch_resolve_pack_taken & btb_159_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_159_bht_T_2 = btb_159_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_159_bht_T_3 = io_i_branch_resolve_pack_taken & btb_159_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_159_bht_T_4 = btb_159_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_159_bht_T_5 = io_i_branch_resolve_pack_taken & btb_159_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_159_bht_T_6 = btb_159_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_159_bht_T_7 = io_i_branch_resolve_pack_taken & btb_159_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_159_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_159_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_159_bht_T_13 = _btb_0_bht_T_8 & _btb_159_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_159_bht_T_16 = _btb_0_bht_T_8 & _btb_159_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_159_bht_T_19 = _btb_0_bht_T_8 & _btb_159_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_159_bht_T_20 = _btb_159_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_21 = _btb_159_bht_T_16 ? 2'h0 : _btb_159_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_22 = _btb_159_bht_T_13 ? 2'h0 : _btb_159_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_23 = _btb_159_bht_T_10 ? 2'h0 : _btb_159_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_24 = _btb_159_bht_T_7 ? 2'h3 : _btb_159_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_25 = _btb_159_bht_T_5 ? 2'h3 : _btb_159_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_26 = _btb_159_bht_T_3 ? 2'h3 : _btb_159_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_159_bht_T_27 = _btb_159_bht_T_1 ? 2'h1 : _btb_159_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9342 = btb_159_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6815
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9344 = btb_159_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_159_bht_T_27 : _GEN_8351; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_160_bht_T = btb_160_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_160_bht_T_1 = io_i_branch_resolve_pack_taken & btb_160_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_160_bht_T_2 = btb_160_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_160_bht_T_3 = io_i_branch_resolve_pack_taken & btb_160_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_160_bht_T_4 = btb_160_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_160_bht_T_5 = io_i_branch_resolve_pack_taken & btb_160_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_160_bht_T_6 = btb_160_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_160_bht_T_7 = io_i_branch_resolve_pack_taken & btb_160_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_160_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_160_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_160_bht_T_13 = _btb_0_bht_T_8 & _btb_160_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_160_bht_T_16 = _btb_0_bht_T_8 & _btb_160_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_160_bht_T_19 = _btb_0_bht_T_8 & _btb_160_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_160_bht_T_20 = _btb_160_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_21 = _btb_160_bht_T_16 ? 2'h0 : _btb_160_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_22 = _btb_160_bht_T_13 ? 2'h0 : _btb_160_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_23 = _btb_160_bht_T_10 ? 2'h0 : _btb_160_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_24 = _btb_160_bht_T_7 ? 2'h3 : _btb_160_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_25 = _btb_160_bht_T_5 ? 2'h3 : _btb_160_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_26 = _btb_160_bht_T_3 ? 2'h3 : _btb_160_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_160_bht_T_27 = _btb_160_bht_T_1 ? 2'h1 : _btb_160_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9346 = btb_160_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6816
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9348 = btb_160_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_160_bht_T_27 : _GEN_8352; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_161_bht_T = btb_161_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_161_bht_T_1 = io_i_branch_resolve_pack_taken & btb_161_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_161_bht_T_2 = btb_161_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_161_bht_T_3 = io_i_branch_resolve_pack_taken & btb_161_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_161_bht_T_4 = btb_161_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_161_bht_T_5 = io_i_branch_resolve_pack_taken & btb_161_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_161_bht_T_6 = btb_161_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_161_bht_T_7 = io_i_branch_resolve_pack_taken & btb_161_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_161_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_161_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_161_bht_T_13 = _btb_0_bht_T_8 & _btb_161_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_161_bht_T_16 = _btb_0_bht_T_8 & _btb_161_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_161_bht_T_19 = _btb_0_bht_T_8 & _btb_161_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_161_bht_T_20 = _btb_161_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_21 = _btb_161_bht_T_16 ? 2'h0 : _btb_161_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_22 = _btb_161_bht_T_13 ? 2'h0 : _btb_161_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_23 = _btb_161_bht_T_10 ? 2'h0 : _btb_161_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_24 = _btb_161_bht_T_7 ? 2'h3 : _btb_161_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_25 = _btb_161_bht_T_5 ? 2'h3 : _btb_161_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_26 = _btb_161_bht_T_3 ? 2'h3 : _btb_161_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_161_bht_T_27 = _btb_161_bht_T_1 ? 2'h1 : _btb_161_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9350 = btb_161_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6817
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9352 = btb_161_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_161_bht_T_27 : _GEN_8353; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_162_bht_T = btb_162_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_162_bht_T_1 = io_i_branch_resolve_pack_taken & btb_162_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_162_bht_T_2 = btb_162_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_162_bht_T_3 = io_i_branch_resolve_pack_taken & btb_162_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_162_bht_T_4 = btb_162_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_162_bht_T_5 = io_i_branch_resolve_pack_taken & btb_162_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_162_bht_T_6 = btb_162_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_162_bht_T_7 = io_i_branch_resolve_pack_taken & btb_162_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_162_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_162_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_162_bht_T_13 = _btb_0_bht_T_8 & _btb_162_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_162_bht_T_16 = _btb_0_bht_T_8 & _btb_162_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_162_bht_T_19 = _btb_0_bht_T_8 & _btb_162_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_162_bht_T_20 = _btb_162_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_21 = _btb_162_bht_T_16 ? 2'h0 : _btb_162_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_22 = _btb_162_bht_T_13 ? 2'h0 : _btb_162_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_23 = _btb_162_bht_T_10 ? 2'h0 : _btb_162_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_24 = _btb_162_bht_T_7 ? 2'h3 : _btb_162_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_25 = _btb_162_bht_T_5 ? 2'h3 : _btb_162_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_26 = _btb_162_bht_T_3 ? 2'h3 : _btb_162_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_162_bht_T_27 = _btb_162_bht_T_1 ? 2'h1 : _btb_162_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9354 = btb_162_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6818
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9356 = btb_162_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_162_bht_T_27 : _GEN_8354; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_163_bht_T = btb_163_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_163_bht_T_1 = io_i_branch_resolve_pack_taken & btb_163_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_163_bht_T_2 = btb_163_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_163_bht_T_3 = io_i_branch_resolve_pack_taken & btb_163_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_163_bht_T_4 = btb_163_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_163_bht_T_5 = io_i_branch_resolve_pack_taken & btb_163_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_163_bht_T_6 = btb_163_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_163_bht_T_7 = io_i_branch_resolve_pack_taken & btb_163_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_163_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_163_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_163_bht_T_13 = _btb_0_bht_T_8 & _btb_163_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_163_bht_T_16 = _btb_0_bht_T_8 & _btb_163_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_163_bht_T_19 = _btb_0_bht_T_8 & _btb_163_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_163_bht_T_20 = _btb_163_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_21 = _btb_163_bht_T_16 ? 2'h0 : _btb_163_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_22 = _btb_163_bht_T_13 ? 2'h0 : _btb_163_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_23 = _btb_163_bht_T_10 ? 2'h0 : _btb_163_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_24 = _btb_163_bht_T_7 ? 2'h3 : _btb_163_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_25 = _btb_163_bht_T_5 ? 2'h3 : _btb_163_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_26 = _btb_163_bht_T_3 ? 2'h3 : _btb_163_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_163_bht_T_27 = _btb_163_bht_T_1 ? 2'h1 : _btb_163_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9358 = btb_163_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6819
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9360 = btb_163_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_163_bht_T_27 : _GEN_8355; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_164_bht_T = btb_164_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_164_bht_T_1 = io_i_branch_resolve_pack_taken & btb_164_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_164_bht_T_2 = btb_164_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_164_bht_T_3 = io_i_branch_resolve_pack_taken & btb_164_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_164_bht_T_4 = btb_164_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_164_bht_T_5 = io_i_branch_resolve_pack_taken & btb_164_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_164_bht_T_6 = btb_164_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_164_bht_T_7 = io_i_branch_resolve_pack_taken & btb_164_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_164_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_164_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_164_bht_T_13 = _btb_0_bht_T_8 & _btb_164_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_164_bht_T_16 = _btb_0_bht_T_8 & _btb_164_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_164_bht_T_19 = _btb_0_bht_T_8 & _btb_164_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_164_bht_T_20 = _btb_164_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_21 = _btb_164_bht_T_16 ? 2'h0 : _btb_164_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_22 = _btb_164_bht_T_13 ? 2'h0 : _btb_164_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_23 = _btb_164_bht_T_10 ? 2'h0 : _btb_164_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_24 = _btb_164_bht_T_7 ? 2'h3 : _btb_164_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_25 = _btb_164_bht_T_5 ? 2'h3 : _btb_164_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_26 = _btb_164_bht_T_3 ? 2'h3 : _btb_164_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_164_bht_T_27 = _btb_164_bht_T_1 ? 2'h1 : _btb_164_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9361 = btb_164_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_163_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_162_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_161_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_160_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_159_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_158_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_157_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_156_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_155_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_154_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_153_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_152_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_151_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_150_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9301)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9362 = btb_164_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6820
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9364 = btb_164_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_164_bht_T_27 : _GEN_8356; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_165_bht_T = btb_165_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_165_bht_T_1 = io_i_branch_resolve_pack_taken & btb_165_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_165_bht_T_2 = btb_165_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_165_bht_T_3 = io_i_branch_resolve_pack_taken & btb_165_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_165_bht_T_4 = btb_165_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_165_bht_T_5 = io_i_branch_resolve_pack_taken & btb_165_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_165_bht_T_6 = btb_165_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_165_bht_T_7 = io_i_branch_resolve_pack_taken & btb_165_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_165_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_165_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_165_bht_T_13 = _btb_0_bht_T_8 & _btb_165_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_165_bht_T_16 = _btb_0_bht_T_8 & _btb_165_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_165_bht_T_19 = _btb_0_bht_T_8 & _btb_165_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_165_bht_T_20 = _btb_165_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_21 = _btb_165_bht_T_16 ? 2'h0 : _btb_165_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_22 = _btb_165_bht_T_13 ? 2'h0 : _btb_165_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_23 = _btb_165_bht_T_10 ? 2'h0 : _btb_165_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_24 = _btb_165_bht_T_7 ? 2'h3 : _btb_165_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_25 = _btb_165_bht_T_5 ? 2'h3 : _btb_165_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_26 = _btb_165_bht_T_3 ? 2'h3 : _btb_165_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_165_bht_T_27 = _btb_165_bht_T_1 ? 2'h1 : _btb_165_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9366 = btb_165_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6821
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9368 = btb_165_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_165_bht_T_27 : _GEN_8357; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_166_bht_T = btb_166_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_166_bht_T_1 = io_i_branch_resolve_pack_taken & btb_166_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_166_bht_T_2 = btb_166_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_166_bht_T_3 = io_i_branch_resolve_pack_taken & btb_166_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_166_bht_T_4 = btb_166_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_166_bht_T_5 = io_i_branch_resolve_pack_taken & btb_166_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_166_bht_T_6 = btb_166_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_166_bht_T_7 = io_i_branch_resolve_pack_taken & btb_166_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_166_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_166_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_166_bht_T_13 = _btb_0_bht_T_8 & _btb_166_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_166_bht_T_16 = _btb_0_bht_T_8 & _btb_166_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_166_bht_T_19 = _btb_0_bht_T_8 & _btb_166_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_166_bht_T_20 = _btb_166_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_21 = _btb_166_bht_T_16 ? 2'h0 : _btb_166_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_22 = _btb_166_bht_T_13 ? 2'h0 : _btb_166_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_23 = _btb_166_bht_T_10 ? 2'h0 : _btb_166_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_24 = _btb_166_bht_T_7 ? 2'h3 : _btb_166_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_25 = _btb_166_bht_T_5 ? 2'h3 : _btb_166_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_26 = _btb_166_bht_T_3 ? 2'h3 : _btb_166_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_166_bht_T_27 = _btb_166_bht_T_1 ? 2'h1 : _btb_166_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9370 = btb_166_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6822
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9372 = btb_166_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_166_bht_T_27 : _GEN_8358; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_167_bht_T = btb_167_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_167_bht_T_1 = io_i_branch_resolve_pack_taken & btb_167_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_167_bht_T_2 = btb_167_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_167_bht_T_3 = io_i_branch_resolve_pack_taken & btb_167_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_167_bht_T_4 = btb_167_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_167_bht_T_5 = io_i_branch_resolve_pack_taken & btb_167_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_167_bht_T_6 = btb_167_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_167_bht_T_7 = io_i_branch_resolve_pack_taken & btb_167_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_167_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_167_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_167_bht_T_13 = _btb_0_bht_T_8 & _btb_167_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_167_bht_T_16 = _btb_0_bht_T_8 & _btb_167_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_167_bht_T_19 = _btb_0_bht_T_8 & _btb_167_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_167_bht_T_20 = _btb_167_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_21 = _btb_167_bht_T_16 ? 2'h0 : _btb_167_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_22 = _btb_167_bht_T_13 ? 2'h0 : _btb_167_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_23 = _btb_167_bht_T_10 ? 2'h0 : _btb_167_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_24 = _btb_167_bht_T_7 ? 2'h3 : _btb_167_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_25 = _btb_167_bht_T_5 ? 2'h3 : _btb_167_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_26 = _btb_167_bht_T_3 ? 2'h3 : _btb_167_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_167_bht_T_27 = _btb_167_bht_T_1 ? 2'h1 : _btb_167_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9374 = btb_167_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6823
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9376 = btb_167_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_167_bht_T_27 : _GEN_8359; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_168_bht_T = btb_168_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_168_bht_T_1 = io_i_branch_resolve_pack_taken & btb_168_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_168_bht_T_2 = btb_168_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_168_bht_T_3 = io_i_branch_resolve_pack_taken & btb_168_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_168_bht_T_4 = btb_168_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_168_bht_T_5 = io_i_branch_resolve_pack_taken & btb_168_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_168_bht_T_6 = btb_168_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_168_bht_T_7 = io_i_branch_resolve_pack_taken & btb_168_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_168_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_168_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_168_bht_T_13 = _btb_0_bht_T_8 & _btb_168_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_168_bht_T_16 = _btb_0_bht_T_8 & _btb_168_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_168_bht_T_19 = _btb_0_bht_T_8 & _btb_168_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_168_bht_T_20 = _btb_168_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_21 = _btb_168_bht_T_16 ? 2'h0 : _btb_168_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_22 = _btb_168_bht_T_13 ? 2'h0 : _btb_168_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_23 = _btb_168_bht_T_10 ? 2'h0 : _btb_168_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_24 = _btb_168_bht_T_7 ? 2'h3 : _btb_168_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_25 = _btb_168_bht_T_5 ? 2'h3 : _btb_168_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_26 = _btb_168_bht_T_3 ? 2'h3 : _btb_168_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_168_bht_T_27 = _btb_168_bht_T_1 ? 2'h1 : _btb_168_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9378 = btb_168_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6824
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9380 = btb_168_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_168_bht_T_27 : _GEN_8360; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_169_bht_T = btb_169_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_169_bht_T_1 = io_i_branch_resolve_pack_taken & btb_169_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_169_bht_T_2 = btb_169_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_169_bht_T_3 = io_i_branch_resolve_pack_taken & btb_169_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_169_bht_T_4 = btb_169_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_169_bht_T_5 = io_i_branch_resolve_pack_taken & btb_169_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_169_bht_T_6 = btb_169_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_169_bht_T_7 = io_i_branch_resolve_pack_taken & btb_169_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_169_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_169_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_169_bht_T_13 = _btb_0_bht_T_8 & _btb_169_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_169_bht_T_16 = _btb_0_bht_T_8 & _btb_169_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_169_bht_T_19 = _btb_0_bht_T_8 & _btb_169_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_169_bht_T_20 = _btb_169_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_21 = _btb_169_bht_T_16 ? 2'h0 : _btb_169_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_22 = _btb_169_bht_T_13 ? 2'h0 : _btb_169_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_23 = _btb_169_bht_T_10 ? 2'h0 : _btb_169_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_24 = _btb_169_bht_T_7 ? 2'h3 : _btb_169_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_25 = _btb_169_bht_T_5 ? 2'h3 : _btb_169_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_26 = _btb_169_bht_T_3 ? 2'h3 : _btb_169_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_169_bht_T_27 = _btb_169_bht_T_1 ? 2'h1 : _btb_169_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9382 = btb_169_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6825
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9384 = btb_169_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_169_bht_T_27 : _GEN_8361; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_170_bht_T = btb_170_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_170_bht_T_1 = io_i_branch_resolve_pack_taken & btb_170_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_170_bht_T_2 = btb_170_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_170_bht_T_3 = io_i_branch_resolve_pack_taken & btb_170_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_170_bht_T_4 = btb_170_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_170_bht_T_5 = io_i_branch_resolve_pack_taken & btb_170_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_170_bht_T_6 = btb_170_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_170_bht_T_7 = io_i_branch_resolve_pack_taken & btb_170_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_170_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_170_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_170_bht_T_13 = _btb_0_bht_T_8 & _btb_170_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_170_bht_T_16 = _btb_0_bht_T_8 & _btb_170_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_170_bht_T_19 = _btb_0_bht_T_8 & _btb_170_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_170_bht_T_20 = _btb_170_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_21 = _btb_170_bht_T_16 ? 2'h0 : _btb_170_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_22 = _btb_170_bht_T_13 ? 2'h0 : _btb_170_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_23 = _btb_170_bht_T_10 ? 2'h0 : _btb_170_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_24 = _btb_170_bht_T_7 ? 2'h3 : _btb_170_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_25 = _btb_170_bht_T_5 ? 2'h3 : _btb_170_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_26 = _btb_170_bht_T_3 ? 2'h3 : _btb_170_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_170_bht_T_27 = _btb_170_bht_T_1 ? 2'h1 : _btb_170_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9386 = btb_170_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6826
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9388 = btb_170_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_170_bht_T_27 : _GEN_8362; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_171_bht_T = btb_171_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_171_bht_T_1 = io_i_branch_resolve_pack_taken & btb_171_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_171_bht_T_2 = btb_171_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_171_bht_T_3 = io_i_branch_resolve_pack_taken & btb_171_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_171_bht_T_4 = btb_171_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_171_bht_T_5 = io_i_branch_resolve_pack_taken & btb_171_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_171_bht_T_6 = btb_171_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_171_bht_T_7 = io_i_branch_resolve_pack_taken & btb_171_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_171_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_171_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_171_bht_T_13 = _btb_0_bht_T_8 & _btb_171_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_171_bht_T_16 = _btb_0_bht_T_8 & _btb_171_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_171_bht_T_19 = _btb_0_bht_T_8 & _btb_171_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_171_bht_T_20 = _btb_171_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_21 = _btb_171_bht_T_16 ? 2'h0 : _btb_171_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_22 = _btb_171_bht_T_13 ? 2'h0 : _btb_171_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_23 = _btb_171_bht_T_10 ? 2'h0 : _btb_171_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_24 = _btb_171_bht_T_7 ? 2'h3 : _btb_171_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_25 = _btb_171_bht_T_5 ? 2'h3 : _btb_171_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_26 = _btb_171_bht_T_3 ? 2'h3 : _btb_171_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_171_bht_T_27 = _btb_171_bht_T_1 ? 2'h1 : _btb_171_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9390 = btb_171_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6827
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9392 = btb_171_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_171_bht_T_27 : _GEN_8363; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_172_bht_T = btb_172_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_172_bht_T_1 = io_i_branch_resolve_pack_taken & btb_172_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_172_bht_T_2 = btb_172_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_172_bht_T_3 = io_i_branch_resolve_pack_taken & btb_172_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_172_bht_T_4 = btb_172_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_172_bht_T_5 = io_i_branch_resolve_pack_taken & btb_172_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_172_bht_T_6 = btb_172_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_172_bht_T_7 = io_i_branch_resolve_pack_taken & btb_172_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_172_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_172_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_172_bht_T_13 = _btb_0_bht_T_8 & _btb_172_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_172_bht_T_16 = _btb_0_bht_T_8 & _btb_172_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_172_bht_T_19 = _btb_0_bht_T_8 & _btb_172_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_172_bht_T_20 = _btb_172_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_21 = _btb_172_bht_T_16 ? 2'h0 : _btb_172_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_22 = _btb_172_bht_T_13 ? 2'h0 : _btb_172_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_23 = _btb_172_bht_T_10 ? 2'h0 : _btb_172_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_24 = _btb_172_bht_T_7 ? 2'h3 : _btb_172_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_25 = _btb_172_bht_T_5 ? 2'h3 : _btb_172_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_26 = _btb_172_bht_T_3 ? 2'h3 : _btb_172_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_172_bht_T_27 = _btb_172_bht_T_1 ? 2'h1 : _btb_172_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9394 = btb_172_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6828
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9396 = btb_172_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_172_bht_T_27 : _GEN_8364; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_173_bht_T = btb_173_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_173_bht_T_1 = io_i_branch_resolve_pack_taken & btb_173_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_173_bht_T_2 = btb_173_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_173_bht_T_3 = io_i_branch_resolve_pack_taken & btb_173_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_173_bht_T_4 = btb_173_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_173_bht_T_5 = io_i_branch_resolve_pack_taken & btb_173_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_173_bht_T_6 = btb_173_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_173_bht_T_7 = io_i_branch_resolve_pack_taken & btb_173_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_173_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_173_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_173_bht_T_13 = _btb_0_bht_T_8 & _btb_173_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_173_bht_T_16 = _btb_0_bht_T_8 & _btb_173_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_173_bht_T_19 = _btb_0_bht_T_8 & _btb_173_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_173_bht_T_20 = _btb_173_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_21 = _btb_173_bht_T_16 ? 2'h0 : _btb_173_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_22 = _btb_173_bht_T_13 ? 2'h0 : _btb_173_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_23 = _btb_173_bht_T_10 ? 2'h0 : _btb_173_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_24 = _btb_173_bht_T_7 ? 2'h3 : _btb_173_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_25 = _btb_173_bht_T_5 ? 2'h3 : _btb_173_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_26 = _btb_173_bht_T_3 ? 2'h3 : _btb_173_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_173_bht_T_27 = _btb_173_bht_T_1 ? 2'h1 : _btb_173_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9398 = btb_173_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6829
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9400 = btb_173_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_173_bht_T_27 : _GEN_8365; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_174_bht_T = btb_174_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_174_bht_T_1 = io_i_branch_resolve_pack_taken & btb_174_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_174_bht_T_2 = btb_174_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_174_bht_T_3 = io_i_branch_resolve_pack_taken & btb_174_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_174_bht_T_4 = btb_174_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_174_bht_T_5 = io_i_branch_resolve_pack_taken & btb_174_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_174_bht_T_6 = btb_174_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_174_bht_T_7 = io_i_branch_resolve_pack_taken & btb_174_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_174_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_174_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_174_bht_T_13 = _btb_0_bht_T_8 & _btb_174_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_174_bht_T_16 = _btb_0_bht_T_8 & _btb_174_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_174_bht_T_19 = _btb_0_bht_T_8 & _btb_174_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_174_bht_T_20 = _btb_174_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_21 = _btb_174_bht_T_16 ? 2'h0 : _btb_174_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_22 = _btb_174_bht_T_13 ? 2'h0 : _btb_174_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_23 = _btb_174_bht_T_10 ? 2'h0 : _btb_174_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_24 = _btb_174_bht_T_7 ? 2'h3 : _btb_174_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_25 = _btb_174_bht_T_5 ? 2'h3 : _btb_174_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_26 = _btb_174_bht_T_3 ? 2'h3 : _btb_174_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_174_bht_T_27 = _btb_174_bht_T_1 ? 2'h1 : _btb_174_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9402 = btb_174_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6830
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9404 = btb_174_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_174_bht_T_27 : _GEN_8366; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_175_bht_T = btb_175_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_175_bht_T_1 = io_i_branch_resolve_pack_taken & btb_175_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_175_bht_T_2 = btb_175_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_175_bht_T_3 = io_i_branch_resolve_pack_taken & btb_175_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_175_bht_T_4 = btb_175_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_175_bht_T_5 = io_i_branch_resolve_pack_taken & btb_175_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_175_bht_T_6 = btb_175_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_175_bht_T_7 = io_i_branch_resolve_pack_taken & btb_175_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_175_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_175_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_175_bht_T_13 = _btb_0_bht_T_8 & _btb_175_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_175_bht_T_16 = _btb_0_bht_T_8 & _btb_175_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_175_bht_T_19 = _btb_0_bht_T_8 & _btb_175_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_175_bht_T_20 = _btb_175_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_21 = _btb_175_bht_T_16 ? 2'h0 : _btb_175_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_22 = _btb_175_bht_T_13 ? 2'h0 : _btb_175_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_23 = _btb_175_bht_T_10 ? 2'h0 : _btb_175_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_24 = _btb_175_bht_T_7 ? 2'h3 : _btb_175_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_25 = _btb_175_bht_T_5 ? 2'h3 : _btb_175_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_26 = _btb_175_bht_T_3 ? 2'h3 : _btb_175_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_175_bht_T_27 = _btb_175_bht_T_1 ? 2'h1 : _btb_175_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9406 = btb_175_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6831
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9408 = btb_175_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_175_bht_T_27 : _GEN_8367; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_176_bht_T = btb_176_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_176_bht_T_1 = io_i_branch_resolve_pack_taken & btb_176_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_176_bht_T_2 = btb_176_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_176_bht_T_3 = io_i_branch_resolve_pack_taken & btb_176_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_176_bht_T_4 = btb_176_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_176_bht_T_5 = io_i_branch_resolve_pack_taken & btb_176_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_176_bht_T_6 = btb_176_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_176_bht_T_7 = io_i_branch_resolve_pack_taken & btb_176_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_176_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_176_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_176_bht_T_13 = _btb_0_bht_T_8 & _btb_176_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_176_bht_T_16 = _btb_0_bht_T_8 & _btb_176_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_176_bht_T_19 = _btb_0_bht_T_8 & _btb_176_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_176_bht_T_20 = _btb_176_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_21 = _btb_176_bht_T_16 ? 2'h0 : _btb_176_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_22 = _btb_176_bht_T_13 ? 2'h0 : _btb_176_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_23 = _btb_176_bht_T_10 ? 2'h0 : _btb_176_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_24 = _btb_176_bht_T_7 ? 2'h3 : _btb_176_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_25 = _btb_176_bht_T_5 ? 2'h3 : _btb_176_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_26 = _btb_176_bht_T_3 ? 2'h3 : _btb_176_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_176_bht_T_27 = _btb_176_bht_T_1 ? 2'h1 : _btb_176_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9410 = btb_176_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6832
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9412 = btb_176_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_176_bht_T_27 : _GEN_8368; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_177_bht_T = btb_177_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_177_bht_T_1 = io_i_branch_resolve_pack_taken & btb_177_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_177_bht_T_2 = btb_177_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_177_bht_T_3 = io_i_branch_resolve_pack_taken & btb_177_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_177_bht_T_4 = btb_177_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_177_bht_T_5 = io_i_branch_resolve_pack_taken & btb_177_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_177_bht_T_6 = btb_177_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_177_bht_T_7 = io_i_branch_resolve_pack_taken & btb_177_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_177_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_177_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_177_bht_T_13 = _btb_0_bht_T_8 & _btb_177_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_177_bht_T_16 = _btb_0_bht_T_8 & _btb_177_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_177_bht_T_19 = _btb_0_bht_T_8 & _btb_177_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_177_bht_T_20 = _btb_177_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_21 = _btb_177_bht_T_16 ? 2'h0 : _btb_177_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_22 = _btb_177_bht_T_13 ? 2'h0 : _btb_177_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_23 = _btb_177_bht_T_10 ? 2'h0 : _btb_177_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_24 = _btb_177_bht_T_7 ? 2'h3 : _btb_177_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_25 = _btb_177_bht_T_5 ? 2'h3 : _btb_177_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_26 = _btb_177_bht_T_3 ? 2'h3 : _btb_177_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_177_bht_T_27 = _btb_177_bht_T_1 ? 2'h1 : _btb_177_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9414 = btb_177_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6833
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9416 = btb_177_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_177_bht_T_27 : _GEN_8369; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_178_bht_T = btb_178_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_178_bht_T_1 = io_i_branch_resolve_pack_taken & btb_178_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_178_bht_T_2 = btb_178_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_178_bht_T_3 = io_i_branch_resolve_pack_taken & btb_178_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_178_bht_T_4 = btb_178_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_178_bht_T_5 = io_i_branch_resolve_pack_taken & btb_178_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_178_bht_T_6 = btb_178_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_178_bht_T_7 = io_i_branch_resolve_pack_taken & btb_178_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_178_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_178_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_178_bht_T_13 = _btb_0_bht_T_8 & _btb_178_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_178_bht_T_16 = _btb_0_bht_T_8 & _btb_178_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_178_bht_T_19 = _btb_0_bht_T_8 & _btb_178_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_178_bht_T_20 = _btb_178_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_21 = _btb_178_bht_T_16 ? 2'h0 : _btb_178_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_22 = _btb_178_bht_T_13 ? 2'h0 : _btb_178_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_23 = _btb_178_bht_T_10 ? 2'h0 : _btb_178_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_24 = _btb_178_bht_T_7 ? 2'h3 : _btb_178_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_25 = _btb_178_bht_T_5 ? 2'h3 : _btb_178_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_26 = _btb_178_bht_T_3 ? 2'h3 : _btb_178_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_178_bht_T_27 = _btb_178_bht_T_1 ? 2'h1 : _btb_178_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9418 = btb_178_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6834
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9420 = btb_178_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_178_bht_T_27 : _GEN_8370; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_179_bht_T = btb_179_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_179_bht_T_1 = io_i_branch_resolve_pack_taken & btb_179_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_179_bht_T_2 = btb_179_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_179_bht_T_3 = io_i_branch_resolve_pack_taken & btb_179_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_179_bht_T_4 = btb_179_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_179_bht_T_5 = io_i_branch_resolve_pack_taken & btb_179_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_179_bht_T_6 = btb_179_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_179_bht_T_7 = io_i_branch_resolve_pack_taken & btb_179_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_179_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_179_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_179_bht_T_13 = _btb_0_bht_T_8 & _btb_179_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_179_bht_T_16 = _btb_0_bht_T_8 & _btb_179_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_179_bht_T_19 = _btb_0_bht_T_8 & _btb_179_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_179_bht_T_20 = _btb_179_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_21 = _btb_179_bht_T_16 ? 2'h0 : _btb_179_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_22 = _btb_179_bht_T_13 ? 2'h0 : _btb_179_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_23 = _btb_179_bht_T_10 ? 2'h0 : _btb_179_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_24 = _btb_179_bht_T_7 ? 2'h3 : _btb_179_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_25 = _btb_179_bht_T_5 ? 2'h3 : _btb_179_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_26 = _btb_179_bht_T_3 ? 2'h3 : _btb_179_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_179_bht_T_27 = _btb_179_bht_T_1 ? 2'h1 : _btb_179_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9421 = btb_179_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_178_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_177_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_176_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_175_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_174_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_173_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_172_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_171_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_170_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_169_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_168_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_167_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_166_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_165_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9361)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9422 = btb_179_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6835
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9424 = btb_179_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_179_bht_T_27 : _GEN_8371; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_180_bht_T = btb_180_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_180_bht_T_1 = io_i_branch_resolve_pack_taken & btb_180_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_180_bht_T_2 = btb_180_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_180_bht_T_3 = io_i_branch_resolve_pack_taken & btb_180_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_180_bht_T_4 = btb_180_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_180_bht_T_5 = io_i_branch_resolve_pack_taken & btb_180_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_180_bht_T_6 = btb_180_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_180_bht_T_7 = io_i_branch_resolve_pack_taken & btb_180_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_180_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_180_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_180_bht_T_13 = _btb_0_bht_T_8 & _btb_180_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_180_bht_T_16 = _btb_0_bht_T_8 & _btb_180_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_180_bht_T_19 = _btb_0_bht_T_8 & _btb_180_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_180_bht_T_20 = _btb_180_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_21 = _btb_180_bht_T_16 ? 2'h0 : _btb_180_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_22 = _btb_180_bht_T_13 ? 2'h0 : _btb_180_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_23 = _btb_180_bht_T_10 ? 2'h0 : _btb_180_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_24 = _btb_180_bht_T_7 ? 2'h3 : _btb_180_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_25 = _btb_180_bht_T_5 ? 2'h3 : _btb_180_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_26 = _btb_180_bht_T_3 ? 2'h3 : _btb_180_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_180_bht_T_27 = _btb_180_bht_T_1 ? 2'h1 : _btb_180_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9426 = btb_180_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6836
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9428 = btb_180_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_180_bht_T_27 : _GEN_8372; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_181_bht_T = btb_181_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_181_bht_T_1 = io_i_branch_resolve_pack_taken & btb_181_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_181_bht_T_2 = btb_181_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_181_bht_T_3 = io_i_branch_resolve_pack_taken & btb_181_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_181_bht_T_4 = btb_181_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_181_bht_T_5 = io_i_branch_resolve_pack_taken & btb_181_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_181_bht_T_6 = btb_181_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_181_bht_T_7 = io_i_branch_resolve_pack_taken & btb_181_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_181_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_181_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_181_bht_T_13 = _btb_0_bht_T_8 & _btb_181_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_181_bht_T_16 = _btb_0_bht_T_8 & _btb_181_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_181_bht_T_19 = _btb_0_bht_T_8 & _btb_181_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_181_bht_T_20 = _btb_181_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_21 = _btb_181_bht_T_16 ? 2'h0 : _btb_181_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_22 = _btb_181_bht_T_13 ? 2'h0 : _btb_181_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_23 = _btb_181_bht_T_10 ? 2'h0 : _btb_181_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_24 = _btb_181_bht_T_7 ? 2'h3 : _btb_181_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_25 = _btb_181_bht_T_5 ? 2'h3 : _btb_181_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_26 = _btb_181_bht_T_3 ? 2'h3 : _btb_181_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_181_bht_T_27 = _btb_181_bht_T_1 ? 2'h1 : _btb_181_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9430 = btb_181_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6837
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9432 = btb_181_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_181_bht_T_27 : _GEN_8373; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_182_bht_T = btb_182_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_182_bht_T_1 = io_i_branch_resolve_pack_taken & btb_182_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_182_bht_T_2 = btb_182_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_182_bht_T_3 = io_i_branch_resolve_pack_taken & btb_182_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_182_bht_T_4 = btb_182_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_182_bht_T_5 = io_i_branch_resolve_pack_taken & btb_182_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_182_bht_T_6 = btb_182_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_182_bht_T_7 = io_i_branch_resolve_pack_taken & btb_182_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_182_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_182_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_182_bht_T_13 = _btb_0_bht_T_8 & _btb_182_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_182_bht_T_16 = _btb_0_bht_T_8 & _btb_182_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_182_bht_T_19 = _btb_0_bht_T_8 & _btb_182_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_182_bht_T_20 = _btb_182_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_21 = _btb_182_bht_T_16 ? 2'h0 : _btb_182_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_22 = _btb_182_bht_T_13 ? 2'h0 : _btb_182_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_23 = _btb_182_bht_T_10 ? 2'h0 : _btb_182_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_24 = _btb_182_bht_T_7 ? 2'h3 : _btb_182_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_25 = _btb_182_bht_T_5 ? 2'h3 : _btb_182_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_26 = _btb_182_bht_T_3 ? 2'h3 : _btb_182_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_182_bht_T_27 = _btb_182_bht_T_1 ? 2'h1 : _btb_182_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9434 = btb_182_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6838
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9436 = btb_182_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_182_bht_T_27 : _GEN_8374; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_183_bht_T = btb_183_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_183_bht_T_1 = io_i_branch_resolve_pack_taken & btb_183_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_183_bht_T_2 = btb_183_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_183_bht_T_3 = io_i_branch_resolve_pack_taken & btb_183_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_183_bht_T_4 = btb_183_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_183_bht_T_5 = io_i_branch_resolve_pack_taken & btb_183_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_183_bht_T_6 = btb_183_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_183_bht_T_7 = io_i_branch_resolve_pack_taken & btb_183_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_183_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_183_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_183_bht_T_13 = _btb_0_bht_T_8 & _btb_183_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_183_bht_T_16 = _btb_0_bht_T_8 & _btb_183_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_183_bht_T_19 = _btb_0_bht_T_8 & _btb_183_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_183_bht_T_20 = _btb_183_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_21 = _btb_183_bht_T_16 ? 2'h0 : _btb_183_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_22 = _btb_183_bht_T_13 ? 2'h0 : _btb_183_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_23 = _btb_183_bht_T_10 ? 2'h0 : _btb_183_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_24 = _btb_183_bht_T_7 ? 2'h3 : _btb_183_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_25 = _btb_183_bht_T_5 ? 2'h3 : _btb_183_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_26 = _btb_183_bht_T_3 ? 2'h3 : _btb_183_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_183_bht_T_27 = _btb_183_bht_T_1 ? 2'h1 : _btb_183_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9438 = btb_183_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6839
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9440 = btb_183_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_183_bht_T_27 : _GEN_8375; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_184_bht_T = btb_184_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_184_bht_T_1 = io_i_branch_resolve_pack_taken & btb_184_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_184_bht_T_2 = btb_184_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_184_bht_T_3 = io_i_branch_resolve_pack_taken & btb_184_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_184_bht_T_4 = btb_184_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_184_bht_T_5 = io_i_branch_resolve_pack_taken & btb_184_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_184_bht_T_6 = btb_184_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_184_bht_T_7 = io_i_branch_resolve_pack_taken & btb_184_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_184_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_184_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_184_bht_T_13 = _btb_0_bht_T_8 & _btb_184_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_184_bht_T_16 = _btb_0_bht_T_8 & _btb_184_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_184_bht_T_19 = _btb_0_bht_T_8 & _btb_184_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_184_bht_T_20 = _btb_184_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_21 = _btb_184_bht_T_16 ? 2'h0 : _btb_184_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_22 = _btb_184_bht_T_13 ? 2'h0 : _btb_184_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_23 = _btb_184_bht_T_10 ? 2'h0 : _btb_184_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_24 = _btb_184_bht_T_7 ? 2'h3 : _btb_184_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_25 = _btb_184_bht_T_5 ? 2'h3 : _btb_184_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_26 = _btb_184_bht_T_3 ? 2'h3 : _btb_184_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_184_bht_T_27 = _btb_184_bht_T_1 ? 2'h1 : _btb_184_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9442 = btb_184_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6840
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9444 = btb_184_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_184_bht_T_27 : _GEN_8376; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_185_bht_T = btb_185_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_185_bht_T_1 = io_i_branch_resolve_pack_taken & btb_185_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_185_bht_T_2 = btb_185_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_185_bht_T_3 = io_i_branch_resolve_pack_taken & btb_185_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_185_bht_T_4 = btb_185_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_185_bht_T_5 = io_i_branch_resolve_pack_taken & btb_185_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_185_bht_T_6 = btb_185_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_185_bht_T_7 = io_i_branch_resolve_pack_taken & btb_185_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_185_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_185_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_185_bht_T_13 = _btb_0_bht_T_8 & _btb_185_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_185_bht_T_16 = _btb_0_bht_T_8 & _btb_185_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_185_bht_T_19 = _btb_0_bht_T_8 & _btb_185_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_185_bht_T_20 = _btb_185_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_21 = _btb_185_bht_T_16 ? 2'h0 : _btb_185_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_22 = _btb_185_bht_T_13 ? 2'h0 : _btb_185_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_23 = _btb_185_bht_T_10 ? 2'h0 : _btb_185_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_24 = _btb_185_bht_T_7 ? 2'h3 : _btb_185_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_25 = _btb_185_bht_T_5 ? 2'h3 : _btb_185_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_26 = _btb_185_bht_T_3 ? 2'h3 : _btb_185_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_185_bht_T_27 = _btb_185_bht_T_1 ? 2'h1 : _btb_185_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9446 = btb_185_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6841
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9448 = btb_185_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_185_bht_T_27 : _GEN_8377; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_186_bht_T = btb_186_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_186_bht_T_1 = io_i_branch_resolve_pack_taken & btb_186_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_186_bht_T_2 = btb_186_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_186_bht_T_3 = io_i_branch_resolve_pack_taken & btb_186_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_186_bht_T_4 = btb_186_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_186_bht_T_5 = io_i_branch_resolve_pack_taken & btb_186_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_186_bht_T_6 = btb_186_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_186_bht_T_7 = io_i_branch_resolve_pack_taken & btb_186_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_186_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_186_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_186_bht_T_13 = _btb_0_bht_T_8 & _btb_186_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_186_bht_T_16 = _btb_0_bht_T_8 & _btb_186_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_186_bht_T_19 = _btb_0_bht_T_8 & _btb_186_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_186_bht_T_20 = _btb_186_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_21 = _btb_186_bht_T_16 ? 2'h0 : _btb_186_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_22 = _btb_186_bht_T_13 ? 2'h0 : _btb_186_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_23 = _btb_186_bht_T_10 ? 2'h0 : _btb_186_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_24 = _btb_186_bht_T_7 ? 2'h3 : _btb_186_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_25 = _btb_186_bht_T_5 ? 2'h3 : _btb_186_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_26 = _btb_186_bht_T_3 ? 2'h3 : _btb_186_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_186_bht_T_27 = _btb_186_bht_T_1 ? 2'h1 : _btb_186_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9450 = btb_186_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6842
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9452 = btb_186_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_186_bht_T_27 : _GEN_8378; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_187_bht_T = btb_187_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_187_bht_T_1 = io_i_branch_resolve_pack_taken & btb_187_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_187_bht_T_2 = btb_187_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_187_bht_T_3 = io_i_branch_resolve_pack_taken & btb_187_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_187_bht_T_4 = btb_187_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_187_bht_T_5 = io_i_branch_resolve_pack_taken & btb_187_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_187_bht_T_6 = btb_187_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_187_bht_T_7 = io_i_branch_resolve_pack_taken & btb_187_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_187_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_187_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_187_bht_T_13 = _btb_0_bht_T_8 & _btb_187_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_187_bht_T_16 = _btb_0_bht_T_8 & _btb_187_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_187_bht_T_19 = _btb_0_bht_T_8 & _btb_187_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_187_bht_T_20 = _btb_187_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_21 = _btb_187_bht_T_16 ? 2'h0 : _btb_187_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_22 = _btb_187_bht_T_13 ? 2'h0 : _btb_187_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_23 = _btb_187_bht_T_10 ? 2'h0 : _btb_187_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_24 = _btb_187_bht_T_7 ? 2'h3 : _btb_187_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_25 = _btb_187_bht_T_5 ? 2'h3 : _btb_187_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_26 = _btb_187_bht_T_3 ? 2'h3 : _btb_187_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_187_bht_T_27 = _btb_187_bht_T_1 ? 2'h1 : _btb_187_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9454 = btb_187_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6843
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9456 = btb_187_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_187_bht_T_27 : _GEN_8379; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_188_bht_T = btb_188_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_188_bht_T_1 = io_i_branch_resolve_pack_taken & btb_188_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_188_bht_T_2 = btb_188_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_188_bht_T_3 = io_i_branch_resolve_pack_taken & btb_188_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_188_bht_T_4 = btb_188_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_188_bht_T_5 = io_i_branch_resolve_pack_taken & btb_188_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_188_bht_T_6 = btb_188_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_188_bht_T_7 = io_i_branch_resolve_pack_taken & btb_188_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_188_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_188_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_188_bht_T_13 = _btb_0_bht_T_8 & _btb_188_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_188_bht_T_16 = _btb_0_bht_T_8 & _btb_188_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_188_bht_T_19 = _btb_0_bht_T_8 & _btb_188_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_188_bht_T_20 = _btb_188_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_21 = _btb_188_bht_T_16 ? 2'h0 : _btb_188_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_22 = _btb_188_bht_T_13 ? 2'h0 : _btb_188_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_23 = _btb_188_bht_T_10 ? 2'h0 : _btb_188_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_24 = _btb_188_bht_T_7 ? 2'h3 : _btb_188_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_25 = _btb_188_bht_T_5 ? 2'h3 : _btb_188_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_26 = _btb_188_bht_T_3 ? 2'h3 : _btb_188_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_188_bht_T_27 = _btb_188_bht_T_1 ? 2'h1 : _btb_188_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9458 = btb_188_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6844
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9460 = btb_188_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_188_bht_T_27 : _GEN_8380; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_189_bht_T = btb_189_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_189_bht_T_1 = io_i_branch_resolve_pack_taken & btb_189_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_189_bht_T_2 = btb_189_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_189_bht_T_3 = io_i_branch_resolve_pack_taken & btb_189_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_189_bht_T_4 = btb_189_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_189_bht_T_5 = io_i_branch_resolve_pack_taken & btb_189_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_189_bht_T_6 = btb_189_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_189_bht_T_7 = io_i_branch_resolve_pack_taken & btb_189_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_189_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_189_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_189_bht_T_13 = _btb_0_bht_T_8 & _btb_189_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_189_bht_T_16 = _btb_0_bht_T_8 & _btb_189_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_189_bht_T_19 = _btb_0_bht_T_8 & _btb_189_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_189_bht_T_20 = _btb_189_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_21 = _btb_189_bht_T_16 ? 2'h0 : _btb_189_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_22 = _btb_189_bht_T_13 ? 2'h0 : _btb_189_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_23 = _btb_189_bht_T_10 ? 2'h0 : _btb_189_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_24 = _btb_189_bht_T_7 ? 2'h3 : _btb_189_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_25 = _btb_189_bht_T_5 ? 2'h3 : _btb_189_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_26 = _btb_189_bht_T_3 ? 2'h3 : _btb_189_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_189_bht_T_27 = _btb_189_bht_T_1 ? 2'h1 : _btb_189_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9462 = btb_189_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6845
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9464 = btb_189_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_189_bht_T_27 : _GEN_8381; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_190_bht_T = btb_190_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_190_bht_T_1 = io_i_branch_resolve_pack_taken & btb_190_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_190_bht_T_2 = btb_190_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_190_bht_T_3 = io_i_branch_resolve_pack_taken & btb_190_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_190_bht_T_4 = btb_190_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_190_bht_T_5 = io_i_branch_resolve_pack_taken & btb_190_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_190_bht_T_6 = btb_190_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_190_bht_T_7 = io_i_branch_resolve_pack_taken & btb_190_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_190_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_190_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_190_bht_T_13 = _btb_0_bht_T_8 & _btb_190_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_190_bht_T_16 = _btb_0_bht_T_8 & _btb_190_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_190_bht_T_19 = _btb_0_bht_T_8 & _btb_190_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_190_bht_T_20 = _btb_190_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_21 = _btb_190_bht_T_16 ? 2'h0 : _btb_190_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_22 = _btb_190_bht_T_13 ? 2'h0 : _btb_190_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_23 = _btb_190_bht_T_10 ? 2'h0 : _btb_190_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_24 = _btb_190_bht_T_7 ? 2'h3 : _btb_190_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_25 = _btb_190_bht_T_5 ? 2'h3 : _btb_190_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_26 = _btb_190_bht_T_3 ? 2'h3 : _btb_190_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_190_bht_T_27 = _btb_190_bht_T_1 ? 2'h1 : _btb_190_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9466 = btb_190_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6846
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9468 = btb_190_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_190_bht_T_27 : _GEN_8382; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_191_bht_T = btb_191_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_191_bht_T_1 = io_i_branch_resolve_pack_taken & btb_191_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_191_bht_T_2 = btb_191_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_191_bht_T_3 = io_i_branch_resolve_pack_taken & btb_191_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_191_bht_T_4 = btb_191_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_191_bht_T_5 = io_i_branch_resolve_pack_taken & btb_191_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_191_bht_T_6 = btb_191_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_191_bht_T_7 = io_i_branch_resolve_pack_taken & btb_191_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_191_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_191_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_191_bht_T_13 = _btb_0_bht_T_8 & _btb_191_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_191_bht_T_16 = _btb_0_bht_T_8 & _btb_191_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_191_bht_T_19 = _btb_0_bht_T_8 & _btb_191_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_191_bht_T_20 = _btb_191_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_21 = _btb_191_bht_T_16 ? 2'h0 : _btb_191_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_22 = _btb_191_bht_T_13 ? 2'h0 : _btb_191_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_23 = _btb_191_bht_T_10 ? 2'h0 : _btb_191_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_24 = _btb_191_bht_T_7 ? 2'h3 : _btb_191_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_25 = _btb_191_bht_T_5 ? 2'h3 : _btb_191_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_26 = _btb_191_bht_T_3 ? 2'h3 : _btb_191_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_191_bht_T_27 = _btb_191_bht_T_1 ? 2'h1 : _btb_191_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9470 = btb_191_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6847
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9472 = btb_191_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_191_bht_T_27 : _GEN_8383; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_192_bht_T = btb_192_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_192_bht_T_1 = io_i_branch_resolve_pack_taken & btb_192_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_192_bht_T_2 = btb_192_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_192_bht_T_3 = io_i_branch_resolve_pack_taken & btb_192_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_192_bht_T_4 = btb_192_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_192_bht_T_5 = io_i_branch_resolve_pack_taken & btb_192_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_192_bht_T_6 = btb_192_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_192_bht_T_7 = io_i_branch_resolve_pack_taken & btb_192_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_192_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_192_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_192_bht_T_13 = _btb_0_bht_T_8 & _btb_192_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_192_bht_T_16 = _btb_0_bht_T_8 & _btb_192_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_192_bht_T_19 = _btb_0_bht_T_8 & _btb_192_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_192_bht_T_20 = _btb_192_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_21 = _btb_192_bht_T_16 ? 2'h0 : _btb_192_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_22 = _btb_192_bht_T_13 ? 2'h0 : _btb_192_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_23 = _btb_192_bht_T_10 ? 2'h0 : _btb_192_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_24 = _btb_192_bht_T_7 ? 2'h3 : _btb_192_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_25 = _btb_192_bht_T_5 ? 2'h3 : _btb_192_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_26 = _btb_192_bht_T_3 ? 2'h3 : _btb_192_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_192_bht_T_27 = _btb_192_bht_T_1 ? 2'h1 : _btb_192_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9474 = btb_192_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6848
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9476 = btb_192_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_192_bht_T_27 : _GEN_8384; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_193_bht_T = btb_193_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_193_bht_T_1 = io_i_branch_resolve_pack_taken & btb_193_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_193_bht_T_2 = btb_193_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_193_bht_T_3 = io_i_branch_resolve_pack_taken & btb_193_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_193_bht_T_4 = btb_193_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_193_bht_T_5 = io_i_branch_resolve_pack_taken & btb_193_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_193_bht_T_6 = btb_193_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_193_bht_T_7 = io_i_branch_resolve_pack_taken & btb_193_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_193_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_193_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_193_bht_T_13 = _btb_0_bht_T_8 & _btb_193_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_193_bht_T_16 = _btb_0_bht_T_8 & _btb_193_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_193_bht_T_19 = _btb_0_bht_T_8 & _btb_193_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_193_bht_T_20 = _btb_193_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_21 = _btb_193_bht_T_16 ? 2'h0 : _btb_193_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_22 = _btb_193_bht_T_13 ? 2'h0 : _btb_193_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_23 = _btb_193_bht_T_10 ? 2'h0 : _btb_193_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_24 = _btb_193_bht_T_7 ? 2'h3 : _btb_193_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_25 = _btb_193_bht_T_5 ? 2'h3 : _btb_193_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_26 = _btb_193_bht_T_3 ? 2'h3 : _btb_193_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_193_bht_T_27 = _btb_193_bht_T_1 ? 2'h1 : _btb_193_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9478 = btb_193_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6849
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9480 = btb_193_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_193_bht_T_27 : _GEN_8385; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_194_bht_T = btb_194_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_194_bht_T_1 = io_i_branch_resolve_pack_taken & btb_194_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_194_bht_T_2 = btb_194_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_194_bht_T_3 = io_i_branch_resolve_pack_taken & btb_194_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_194_bht_T_4 = btb_194_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_194_bht_T_5 = io_i_branch_resolve_pack_taken & btb_194_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_194_bht_T_6 = btb_194_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_194_bht_T_7 = io_i_branch_resolve_pack_taken & btb_194_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_194_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_194_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_194_bht_T_13 = _btb_0_bht_T_8 & _btb_194_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_194_bht_T_16 = _btb_0_bht_T_8 & _btb_194_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_194_bht_T_19 = _btb_0_bht_T_8 & _btb_194_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_194_bht_T_20 = _btb_194_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_21 = _btb_194_bht_T_16 ? 2'h0 : _btb_194_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_22 = _btb_194_bht_T_13 ? 2'h0 : _btb_194_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_23 = _btb_194_bht_T_10 ? 2'h0 : _btb_194_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_24 = _btb_194_bht_T_7 ? 2'h3 : _btb_194_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_25 = _btb_194_bht_T_5 ? 2'h3 : _btb_194_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_26 = _btb_194_bht_T_3 ? 2'h3 : _btb_194_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_194_bht_T_27 = _btb_194_bht_T_1 ? 2'h1 : _btb_194_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9481 = btb_194_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_193_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_192_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_191_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_190_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_189_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_188_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_187_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_186_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_185_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_184_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_183_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_182_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_181_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_180_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9421)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9482 = btb_194_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6850
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9484 = btb_194_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_194_bht_T_27 : _GEN_8386; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_195_bht_T = btb_195_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_195_bht_T_1 = io_i_branch_resolve_pack_taken & btb_195_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_195_bht_T_2 = btb_195_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_195_bht_T_3 = io_i_branch_resolve_pack_taken & btb_195_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_195_bht_T_4 = btb_195_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_195_bht_T_5 = io_i_branch_resolve_pack_taken & btb_195_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_195_bht_T_6 = btb_195_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_195_bht_T_7 = io_i_branch_resolve_pack_taken & btb_195_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_195_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_195_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_195_bht_T_13 = _btb_0_bht_T_8 & _btb_195_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_195_bht_T_16 = _btb_0_bht_T_8 & _btb_195_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_195_bht_T_19 = _btb_0_bht_T_8 & _btb_195_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_195_bht_T_20 = _btb_195_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_21 = _btb_195_bht_T_16 ? 2'h0 : _btb_195_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_22 = _btb_195_bht_T_13 ? 2'h0 : _btb_195_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_23 = _btb_195_bht_T_10 ? 2'h0 : _btb_195_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_24 = _btb_195_bht_T_7 ? 2'h3 : _btb_195_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_25 = _btb_195_bht_T_5 ? 2'h3 : _btb_195_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_26 = _btb_195_bht_T_3 ? 2'h3 : _btb_195_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_195_bht_T_27 = _btb_195_bht_T_1 ? 2'h1 : _btb_195_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9486 = btb_195_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6851
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9488 = btb_195_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_195_bht_T_27 : _GEN_8387; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_196_bht_T = btb_196_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_196_bht_T_1 = io_i_branch_resolve_pack_taken & btb_196_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_196_bht_T_2 = btb_196_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_196_bht_T_3 = io_i_branch_resolve_pack_taken & btb_196_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_196_bht_T_4 = btb_196_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_196_bht_T_5 = io_i_branch_resolve_pack_taken & btb_196_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_196_bht_T_6 = btb_196_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_196_bht_T_7 = io_i_branch_resolve_pack_taken & btb_196_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_196_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_196_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_196_bht_T_13 = _btb_0_bht_T_8 & _btb_196_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_196_bht_T_16 = _btb_0_bht_T_8 & _btb_196_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_196_bht_T_19 = _btb_0_bht_T_8 & _btb_196_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_196_bht_T_20 = _btb_196_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_21 = _btb_196_bht_T_16 ? 2'h0 : _btb_196_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_22 = _btb_196_bht_T_13 ? 2'h0 : _btb_196_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_23 = _btb_196_bht_T_10 ? 2'h0 : _btb_196_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_24 = _btb_196_bht_T_7 ? 2'h3 : _btb_196_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_25 = _btb_196_bht_T_5 ? 2'h3 : _btb_196_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_26 = _btb_196_bht_T_3 ? 2'h3 : _btb_196_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_196_bht_T_27 = _btb_196_bht_T_1 ? 2'h1 : _btb_196_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9490 = btb_196_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6852
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9492 = btb_196_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_196_bht_T_27 : _GEN_8388; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_197_bht_T = btb_197_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_197_bht_T_1 = io_i_branch_resolve_pack_taken & btb_197_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_197_bht_T_2 = btb_197_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_197_bht_T_3 = io_i_branch_resolve_pack_taken & btb_197_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_197_bht_T_4 = btb_197_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_197_bht_T_5 = io_i_branch_resolve_pack_taken & btb_197_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_197_bht_T_6 = btb_197_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_197_bht_T_7 = io_i_branch_resolve_pack_taken & btb_197_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_197_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_197_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_197_bht_T_13 = _btb_0_bht_T_8 & _btb_197_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_197_bht_T_16 = _btb_0_bht_T_8 & _btb_197_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_197_bht_T_19 = _btb_0_bht_T_8 & _btb_197_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_197_bht_T_20 = _btb_197_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_21 = _btb_197_bht_T_16 ? 2'h0 : _btb_197_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_22 = _btb_197_bht_T_13 ? 2'h0 : _btb_197_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_23 = _btb_197_bht_T_10 ? 2'h0 : _btb_197_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_24 = _btb_197_bht_T_7 ? 2'h3 : _btb_197_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_25 = _btb_197_bht_T_5 ? 2'h3 : _btb_197_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_26 = _btb_197_bht_T_3 ? 2'h3 : _btb_197_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_197_bht_T_27 = _btb_197_bht_T_1 ? 2'h1 : _btb_197_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9494 = btb_197_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6853
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9496 = btb_197_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_197_bht_T_27 : _GEN_8389; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_198_bht_T = btb_198_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_198_bht_T_1 = io_i_branch_resolve_pack_taken & btb_198_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_198_bht_T_2 = btb_198_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_198_bht_T_3 = io_i_branch_resolve_pack_taken & btb_198_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_198_bht_T_4 = btb_198_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_198_bht_T_5 = io_i_branch_resolve_pack_taken & btb_198_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_198_bht_T_6 = btb_198_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_198_bht_T_7 = io_i_branch_resolve_pack_taken & btb_198_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_198_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_198_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_198_bht_T_13 = _btb_0_bht_T_8 & _btb_198_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_198_bht_T_16 = _btb_0_bht_T_8 & _btb_198_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_198_bht_T_19 = _btb_0_bht_T_8 & _btb_198_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_198_bht_T_20 = _btb_198_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_21 = _btb_198_bht_T_16 ? 2'h0 : _btb_198_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_22 = _btb_198_bht_T_13 ? 2'h0 : _btb_198_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_23 = _btb_198_bht_T_10 ? 2'h0 : _btb_198_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_24 = _btb_198_bht_T_7 ? 2'h3 : _btb_198_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_25 = _btb_198_bht_T_5 ? 2'h3 : _btb_198_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_26 = _btb_198_bht_T_3 ? 2'h3 : _btb_198_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_198_bht_T_27 = _btb_198_bht_T_1 ? 2'h1 : _btb_198_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9498 = btb_198_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6854
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9500 = btb_198_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_198_bht_T_27 : _GEN_8390; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_199_bht_T = btb_199_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_199_bht_T_1 = io_i_branch_resolve_pack_taken & btb_199_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_199_bht_T_2 = btb_199_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_199_bht_T_3 = io_i_branch_resolve_pack_taken & btb_199_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_199_bht_T_4 = btb_199_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_199_bht_T_5 = io_i_branch_resolve_pack_taken & btb_199_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_199_bht_T_6 = btb_199_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_199_bht_T_7 = io_i_branch_resolve_pack_taken & btb_199_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_199_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_199_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_199_bht_T_13 = _btb_0_bht_T_8 & _btb_199_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_199_bht_T_16 = _btb_0_bht_T_8 & _btb_199_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_199_bht_T_19 = _btb_0_bht_T_8 & _btb_199_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_199_bht_T_20 = _btb_199_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_21 = _btb_199_bht_T_16 ? 2'h0 : _btb_199_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_22 = _btb_199_bht_T_13 ? 2'h0 : _btb_199_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_23 = _btb_199_bht_T_10 ? 2'h0 : _btb_199_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_24 = _btb_199_bht_T_7 ? 2'h3 : _btb_199_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_25 = _btb_199_bht_T_5 ? 2'h3 : _btb_199_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_26 = _btb_199_bht_T_3 ? 2'h3 : _btb_199_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_199_bht_T_27 = _btb_199_bht_T_1 ? 2'h1 : _btb_199_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9502 = btb_199_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6855
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9504 = btb_199_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_199_bht_T_27 : _GEN_8391; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_200_bht_T = btb_200_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_200_bht_T_1 = io_i_branch_resolve_pack_taken & btb_200_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_200_bht_T_2 = btb_200_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_200_bht_T_3 = io_i_branch_resolve_pack_taken & btb_200_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_200_bht_T_4 = btb_200_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_200_bht_T_5 = io_i_branch_resolve_pack_taken & btb_200_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_200_bht_T_6 = btb_200_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_200_bht_T_7 = io_i_branch_resolve_pack_taken & btb_200_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_200_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_200_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_200_bht_T_13 = _btb_0_bht_T_8 & _btb_200_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_200_bht_T_16 = _btb_0_bht_T_8 & _btb_200_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_200_bht_T_19 = _btb_0_bht_T_8 & _btb_200_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_200_bht_T_20 = _btb_200_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_21 = _btb_200_bht_T_16 ? 2'h0 : _btb_200_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_22 = _btb_200_bht_T_13 ? 2'h0 : _btb_200_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_23 = _btb_200_bht_T_10 ? 2'h0 : _btb_200_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_24 = _btb_200_bht_T_7 ? 2'h3 : _btb_200_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_25 = _btb_200_bht_T_5 ? 2'h3 : _btb_200_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_26 = _btb_200_bht_T_3 ? 2'h3 : _btb_200_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_200_bht_T_27 = _btb_200_bht_T_1 ? 2'h1 : _btb_200_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9506 = btb_200_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6856
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9508 = btb_200_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_200_bht_T_27 : _GEN_8392; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_201_bht_T = btb_201_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_201_bht_T_1 = io_i_branch_resolve_pack_taken & btb_201_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_201_bht_T_2 = btb_201_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_201_bht_T_3 = io_i_branch_resolve_pack_taken & btb_201_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_201_bht_T_4 = btb_201_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_201_bht_T_5 = io_i_branch_resolve_pack_taken & btb_201_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_201_bht_T_6 = btb_201_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_201_bht_T_7 = io_i_branch_resolve_pack_taken & btb_201_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_201_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_201_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_201_bht_T_13 = _btb_0_bht_T_8 & _btb_201_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_201_bht_T_16 = _btb_0_bht_T_8 & _btb_201_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_201_bht_T_19 = _btb_0_bht_T_8 & _btb_201_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_201_bht_T_20 = _btb_201_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_21 = _btb_201_bht_T_16 ? 2'h0 : _btb_201_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_22 = _btb_201_bht_T_13 ? 2'h0 : _btb_201_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_23 = _btb_201_bht_T_10 ? 2'h0 : _btb_201_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_24 = _btb_201_bht_T_7 ? 2'h3 : _btb_201_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_25 = _btb_201_bht_T_5 ? 2'h3 : _btb_201_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_26 = _btb_201_bht_T_3 ? 2'h3 : _btb_201_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_201_bht_T_27 = _btb_201_bht_T_1 ? 2'h1 : _btb_201_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9510 = btb_201_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6857
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9512 = btb_201_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_201_bht_T_27 : _GEN_8393; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_202_bht_T = btb_202_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_202_bht_T_1 = io_i_branch_resolve_pack_taken & btb_202_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_202_bht_T_2 = btb_202_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_202_bht_T_3 = io_i_branch_resolve_pack_taken & btb_202_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_202_bht_T_4 = btb_202_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_202_bht_T_5 = io_i_branch_resolve_pack_taken & btb_202_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_202_bht_T_6 = btb_202_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_202_bht_T_7 = io_i_branch_resolve_pack_taken & btb_202_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_202_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_202_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_202_bht_T_13 = _btb_0_bht_T_8 & _btb_202_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_202_bht_T_16 = _btb_0_bht_T_8 & _btb_202_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_202_bht_T_19 = _btb_0_bht_T_8 & _btb_202_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_202_bht_T_20 = _btb_202_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_21 = _btb_202_bht_T_16 ? 2'h0 : _btb_202_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_22 = _btb_202_bht_T_13 ? 2'h0 : _btb_202_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_23 = _btb_202_bht_T_10 ? 2'h0 : _btb_202_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_24 = _btb_202_bht_T_7 ? 2'h3 : _btb_202_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_25 = _btb_202_bht_T_5 ? 2'h3 : _btb_202_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_26 = _btb_202_bht_T_3 ? 2'h3 : _btb_202_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_202_bht_T_27 = _btb_202_bht_T_1 ? 2'h1 : _btb_202_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9514 = btb_202_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6858
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9516 = btb_202_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_202_bht_T_27 : _GEN_8394; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_203_bht_T = btb_203_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_203_bht_T_1 = io_i_branch_resolve_pack_taken & btb_203_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_203_bht_T_2 = btb_203_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_203_bht_T_3 = io_i_branch_resolve_pack_taken & btb_203_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_203_bht_T_4 = btb_203_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_203_bht_T_5 = io_i_branch_resolve_pack_taken & btb_203_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_203_bht_T_6 = btb_203_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_203_bht_T_7 = io_i_branch_resolve_pack_taken & btb_203_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_203_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_203_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_203_bht_T_13 = _btb_0_bht_T_8 & _btb_203_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_203_bht_T_16 = _btb_0_bht_T_8 & _btb_203_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_203_bht_T_19 = _btb_0_bht_T_8 & _btb_203_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_203_bht_T_20 = _btb_203_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_21 = _btb_203_bht_T_16 ? 2'h0 : _btb_203_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_22 = _btb_203_bht_T_13 ? 2'h0 : _btb_203_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_23 = _btb_203_bht_T_10 ? 2'h0 : _btb_203_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_24 = _btb_203_bht_T_7 ? 2'h3 : _btb_203_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_25 = _btb_203_bht_T_5 ? 2'h3 : _btb_203_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_26 = _btb_203_bht_T_3 ? 2'h3 : _btb_203_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_203_bht_T_27 = _btb_203_bht_T_1 ? 2'h1 : _btb_203_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9518 = btb_203_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6859
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9520 = btb_203_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_203_bht_T_27 : _GEN_8395; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_204_bht_T = btb_204_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_204_bht_T_1 = io_i_branch_resolve_pack_taken & btb_204_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_204_bht_T_2 = btb_204_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_204_bht_T_3 = io_i_branch_resolve_pack_taken & btb_204_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_204_bht_T_4 = btb_204_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_204_bht_T_5 = io_i_branch_resolve_pack_taken & btb_204_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_204_bht_T_6 = btb_204_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_204_bht_T_7 = io_i_branch_resolve_pack_taken & btb_204_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_204_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_204_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_204_bht_T_13 = _btb_0_bht_T_8 & _btb_204_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_204_bht_T_16 = _btb_0_bht_T_8 & _btb_204_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_204_bht_T_19 = _btb_0_bht_T_8 & _btb_204_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_204_bht_T_20 = _btb_204_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_21 = _btb_204_bht_T_16 ? 2'h0 : _btb_204_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_22 = _btb_204_bht_T_13 ? 2'h0 : _btb_204_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_23 = _btb_204_bht_T_10 ? 2'h0 : _btb_204_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_24 = _btb_204_bht_T_7 ? 2'h3 : _btb_204_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_25 = _btb_204_bht_T_5 ? 2'h3 : _btb_204_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_26 = _btb_204_bht_T_3 ? 2'h3 : _btb_204_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_204_bht_T_27 = _btb_204_bht_T_1 ? 2'h1 : _btb_204_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9522 = btb_204_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6860
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9524 = btb_204_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_204_bht_T_27 : _GEN_8396; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_205_bht_T = btb_205_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_205_bht_T_1 = io_i_branch_resolve_pack_taken & btb_205_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_205_bht_T_2 = btb_205_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_205_bht_T_3 = io_i_branch_resolve_pack_taken & btb_205_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_205_bht_T_4 = btb_205_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_205_bht_T_5 = io_i_branch_resolve_pack_taken & btb_205_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_205_bht_T_6 = btb_205_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_205_bht_T_7 = io_i_branch_resolve_pack_taken & btb_205_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_205_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_205_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_205_bht_T_13 = _btb_0_bht_T_8 & _btb_205_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_205_bht_T_16 = _btb_0_bht_T_8 & _btb_205_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_205_bht_T_19 = _btb_0_bht_T_8 & _btb_205_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_205_bht_T_20 = _btb_205_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_21 = _btb_205_bht_T_16 ? 2'h0 : _btb_205_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_22 = _btb_205_bht_T_13 ? 2'h0 : _btb_205_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_23 = _btb_205_bht_T_10 ? 2'h0 : _btb_205_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_24 = _btb_205_bht_T_7 ? 2'h3 : _btb_205_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_25 = _btb_205_bht_T_5 ? 2'h3 : _btb_205_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_26 = _btb_205_bht_T_3 ? 2'h3 : _btb_205_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_205_bht_T_27 = _btb_205_bht_T_1 ? 2'h1 : _btb_205_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9526 = btb_205_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6861
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9528 = btb_205_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_205_bht_T_27 : _GEN_8397; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_206_bht_T = btb_206_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_206_bht_T_1 = io_i_branch_resolve_pack_taken & btb_206_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_206_bht_T_2 = btb_206_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_206_bht_T_3 = io_i_branch_resolve_pack_taken & btb_206_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_206_bht_T_4 = btb_206_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_206_bht_T_5 = io_i_branch_resolve_pack_taken & btb_206_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_206_bht_T_6 = btb_206_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_206_bht_T_7 = io_i_branch_resolve_pack_taken & btb_206_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_206_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_206_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_206_bht_T_13 = _btb_0_bht_T_8 & _btb_206_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_206_bht_T_16 = _btb_0_bht_T_8 & _btb_206_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_206_bht_T_19 = _btb_0_bht_T_8 & _btb_206_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_206_bht_T_20 = _btb_206_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_21 = _btb_206_bht_T_16 ? 2'h0 : _btb_206_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_22 = _btb_206_bht_T_13 ? 2'h0 : _btb_206_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_23 = _btb_206_bht_T_10 ? 2'h0 : _btb_206_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_24 = _btb_206_bht_T_7 ? 2'h3 : _btb_206_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_25 = _btb_206_bht_T_5 ? 2'h3 : _btb_206_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_26 = _btb_206_bht_T_3 ? 2'h3 : _btb_206_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_206_bht_T_27 = _btb_206_bht_T_1 ? 2'h1 : _btb_206_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9530 = btb_206_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6862
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9532 = btb_206_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_206_bht_T_27 : _GEN_8398; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_207_bht_T = btb_207_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_207_bht_T_1 = io_i_branch_resolve_pack_taken & btb_207_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_207_bht_T_2 = btb_207_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_207_bht_T_3 = io_i_branch_resolve_pack_taken & btb_207_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_207_bht_T_4 = btb_207_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_207_bht_T_5 = io_i_branch_resolve_pack_taken & btb_207_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_207_bht_T_6 = btb_207_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_207_bht_T_7 = io_i_branch_resolve_pack_taken & btb_207_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_207_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_207_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_207_bht_T_13 = _btb_0_bht_T_8 & _btb_207_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_207_bht_T_16 = _btb_0_bht_T_8 & _btb_207_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_207_bht_T_19 = _btb_0_bht_T_8 & _btb_207_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_207_bht_T_20 = _btb_207_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_21 = _btb_207_bht_T_16 ? 2'h0 : _btb_207_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_22 = _btb_207_bht_T_13 ? 2'h0 : _btb_207_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_23 = _btb_207_bht_T_10 ? 2'h0 : _btb_207_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_24 = _btb_207_bht_T_7 ? 2'h3 : _btb_207_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_25 = _btb_207_bht_T_5 ? 2'h3 : _btb_207_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_26 = _btb_207_bht_T_3 ? 2'h3 : _btb_207_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_207_bht_T_27 = _btb_207_bht_T_1 ? 2'h1 : _btb_207_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9534 = btb_207_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6863
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9536 = btb_207_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_207_bht_T_27 : _GEN_8399; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_208_bht_T = btb_208_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_208_bht_T_1 = io_i_branch_resolve_pack_taken & btb_208_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_208_bht_T_2 = btb_208_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_208_bht_T_3 = io_i_branch_resolve_pack_taken & btb_208_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_208_bht_T_4 = btb_208_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_208_bht_T_5 = io_i_branch_resolve_pack_taken & btb_208_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_208_bht_T_6 = btb_208_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_208_bht_T_7 = io_i_branch_resolve_pack_taken & btb_208_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_208_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_208_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_208_bht_T_13 = _btb_0_bht_T_8 & _btb_208_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_208_bht_T_16 = _btb_0_bht_T_8 & _btb_208_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_208_bht_T_19 = _btb_0_bht_T_8 & _btb_208_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_208_bht_T_20 = _btb_208_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_21 = _btb_208_bht_T_16 ? 2'h0 : _btb_208_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_22 = _btb_208_bht_T_13 ? 2'h0 : _btb_208_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_23 = _btb_208_bht_T_10 ? 2'h0 : _btb_208_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_24 = _btb_208_bht_T_7 ? 2'h3 : _btb_208_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_25 = _btb_208_bht_T_5 ? 2'h3 : _btb_208_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_26 = _btb_208_bht_T_3 ? 2'h3 : _btb_208_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_208_bht_T_27 = _btb_208_bht_T_1 ? 2'h1 : _btb_208_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9538 = btb_208_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6864
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9540 = btb_208_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_208_bht_T_27 : _GEN_8400; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_209_bht_T = btb_209_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_209_bht_T_1 = io_i_branch_resolve_pack_taken & btb_209_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_209_bht_T_2 = btb_209_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_209_bht_T_3 = io_i_branch_resolve_pack_taken & btb_209_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_209_bht_T_4 = btb_209_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_209_bht_T_5 = io_i_branch_resolve_pack_taken & btb_209_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_209_bht_T_6 = btb_209_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_209_bht_T_7 = io_i_branch_resolve_pack_taken & btb_209_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_209_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_209_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_209_bht_T_13 = _btb_0_bht_T_8 & _btb_209_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_209_bht_T_16 = _btb_0_bht_T_8 & _btb_209_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_209_bht_T_19 = _btb_0_bht_T_8 & _btb_209_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_209_bht_T_20 = _btb_209_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_21 = _btb_209_bht_T_16 ? 2'h0 : _btb_209_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_22 = _btb_209_bht_T_13 ? 2'h0 : _btb_209_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_23 = _btb_209_bht_T_10 ? 2'h0 : _btb_209_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_24 = _btb_209_bht_T_7 ? 2'h3 : _btb_209_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_25 = _btb_209_bht_T_5 ? 2'h3 : _btb_209_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_26 = _btb_209_bht_T_3 ? 2'h3 : _btb_209_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_209_bht_T_27 = _btb_209_bht_T_1 ? 2'h1 : _btb_209_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9541 = btb_209_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_208_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_207_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_206_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_205_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_204_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_203_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_202_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_201_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_200_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_199_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_198_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_197_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_196_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_195_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9481)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9542 = btb_209_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6865
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9544 = btb_209_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_209_bht_T_27 : _GEN_8401; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_210_bht_T = btb_210_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_210_bht_T_1 = io_i_branch_resolve_pack_taken & btb_210_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_210_bht_T_2 = btb_210_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_210_bht_T_3 = io_i_branch_resolve_pack_taken & btb_210_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_210_bht_T_4 = btb_210_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_210_bht_T_5 = io_i_branch_resolve_pack_taken & btb_210_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_210_bht_T_6 = btb_210_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_210_bht_T_7 = io_i_branch_resolve_pack_taken & btb_210_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_210_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_210_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_210_bht_T_13 = _btb_0_bht_T_8 & _btb_210_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_210_bht_T_16 = _btb_0_bht_T_8 & _btb_210_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_210_bht_T_19 = _btb_0_bht_T_8 & _btb_210_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_210_bht_T_20 = _btb_210_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_21 = _btb_210_bht_T_16 ? 2'h0 : _btb_210_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_22 = _btb_210_bht_T_13 ? 2'h0 : _btb_210_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_23 = _btb_210_bht_T_10 ? 2'h0 : _btb_210_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_24 = _btb_210_bht_T_7 ? 2'h3 : _btb_210_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_25 = _btb_210_bht_T_5 ? 2'h3 : _btb_210_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_26 = _btb_210_bht_T_3 ? 2'h3 : _btb_210_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_210_bht_T_27 = _btb_210_bht_T_1 ? 2'h1 : _btb_210_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9546 = btb_210_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6866
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9548 = btb_210_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_210_bht_T_27 : _GEN_8402; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_211_bht_T = btb_211_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_211_bht_T_1 = io_i_branch_resolve_pack_taken & btb_211_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_211_bht_T_2 = btb_211_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_211_bht_T_3 = io_i_branch_resolve_pack_taken & btb_211_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_211_bht_T_4 = btb_211_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_211_bht_T_5 = io_i_branch_resolve_pack_taken & btb_211_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_211_bht_T_6 = btb_211_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_211_bht_T_7 = io_i_branch_resolve_pack_taken & btb_211_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_211_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_211_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_211_bht_T_13 = _btb_0_bht_T_8 & _btb_211_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_211_bht_T_16 = _btb_0_bht_T_8 & _btb_211_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_211_bht_T_19 = _btb_0_bht_T_8 & _btb_211_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_211_bht_T_20 = _btb_211_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_21 = _btb_211_bht_T_16 ? 2'h0 : _btb_211_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_22 = _btb_211_bht_T_13 ? 2'h0 : _btb_211_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_23 = _btb_211_bht_T_10 ? 2'h0 : _btb_211_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_24 = _btb_211_bht_T_7 ? 2'h3 : _btb_211_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_25 = _btb_211_bht_T_5 ? 2'h3 : _btb_211_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_26 = _btb_211_bht_T_3 ? 2'h3 : _btb_211_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_211_bht_T_27 = _btb_211_bht_T_1 ? 2'h1 : _btb_211_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9550 = btb_211_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6867
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9552 = btb_211_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_211_bht_T_27 : _GEN_8403; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_212_bht_T = btb_212_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_212_bht_T_1 = io_i_branch_resolve_pack_taken & btb_212_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_212_bht_T_2 = btb_212_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_212_bht_T_3 = io_i_branch_resolve_pack_taken & btb_212_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_212_bht_T_4 = btb_212_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_212_bht_T_5 = io_i_branch_resolve_pack_taken & btb_212_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_212_bht_T_6 = btb_212_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_212_bht_T_7 = io_i_branch_resolve_pack_taken & btb_212_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_212_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_212_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_212_bht_T_13 = _btb_0_bht_T_8 & _btb_212_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_212_bht_T_16 = _btb_0_bht_T_8 & _btb_212_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_212_bht_T_19 = _btb_0_bht_T_8 & _btb_212_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_212_bht_T_20 = _btb_212_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_21 = _btb_212_bht_T_16 ? 2'h0 : _btb_212_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_22 = _btb_212_bht_T_13 ? 2'h0 : _btb_212_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_23 = _btb_212_bht_T_10 ? 2'h0 : _btb_212_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_24 = _btb_212_bht_T_7 ? 2'h3 : _btb_212_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_25 = _btb_212_bht_T_5 ? 2'h3 : _btb_212_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_26 = _btb_212_bht_T_3 ? 2'h3 : _btb_212_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_212_bht_T_27 = _btb_212_bht_T_1 ? 2'h1 : _btb_212_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9554 = btb_212_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6868
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9556 = btb_212_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_212_bht_T_27 : _GEN_8404; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_213_bht_T = btb_213_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_213_bht_T_1 = io_i_branch_resolve_pack_taken & btb_213_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_213_bht_T_2 = btb_213_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_213_bht_T_3 = io_i_branch_resolve_pack_taken & btb_213_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_213_bht_T_4 = btb_213_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_213_bht_T_5 = io_i_branch_resolve_pack_taken & btb_213_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_213_bht_T_6 = btb_213_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_213_bht_T_7 = io_i_branch_resolve_pack_taken & btb_213_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_213_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_213_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_213_bht_T_13 = _btb_0_bht_T_8 & _btb_213_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_213_bht_T_16 = _btb_0_bht_T_8 & _btb_213_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_213_bht_T_19 = _btb_0_bht_T_8 & _btb_213_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_213_bht_T_20 = _btb_213_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_21 = _btb_213_bht_T_16 ? 2'h0 : _btb_213_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_22 = _btb_213_bht_T_13 ? 2'h0 : _btb_213_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_23 = _btb_213_bht_T_10 ? 2'h0 : _btb_213_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_24 = _btb_213_bht_T_7 ? 2'h3 : _btb_213_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_25 = _btb_213_bht_T_5 ? 2'h3 : _btb_213_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_26 = _btb_213_bht_T_3 ? 2'h3 : _btb_213_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_213_bht_T_27 = _btb_213_bht_T_1 ? 2'h1 : _btb_213_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9558 = btb_213_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6869
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9560 = btb_213_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_213_bht_T_27 : _GEN_8405; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_214_bht_T = btb_214_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_214_bht_T_1 = io_i_branch_resolve_pack_taken & btb_214_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_214_bht_T_2 = btb_214_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_214_bht_T_3 = io_i_branch_resolve_pack_taken & btb_214_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_214_bht_T_4 = btb_214_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_214_bht_T_5 = io_i_branch_resolve_pack_taken & btb_214_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_214_bht_T_6 = btb_214_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_214_bht_T_7 = io_i_branch_resolve_pack_taken & btb_214_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_214_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_214_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_214_bht_T_13 = _btb_0_bht_T_8 & _btb_214_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_214_bht_T_16 = _btb_0_bht_T_8 & _btb_214_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_214_bht_T_19 = _btb_0_bht_T_8 & _btb_214_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_214_bht_T_20 = _btb_214_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_21 = _btb_214_bht_T_16 ? 2'h0 : _btb_214_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_22 = _btb_214_bht_T_13 ? 2'h0 : _btb_214_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_23 = _btb_214_bht_T_10 ? 2'h0 : _btb_214_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_24 = _btb_214_bht_T_7 ? 2'h3 : _btb_214_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_25 = _btb_214_bht_T_5 ? 2'h3 : _btb_214_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_26 = _btb_214_bht_T_3 ? 2'h3 : _btb_214_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_214_bht_T_27 = _btb_214_bht_T_1 ? 2'h1 : _btb_214_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9562 = btb_214_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6870
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9564 = btb_214_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_214_bht_T_27 : _GEN_8406; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_215_bht_T = btb_215_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_215_bht_T_1 = io_i_branch_resolve_pack_taken & btb_215_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_215_bht_T_2 = btb_215_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_215_bht_T_3 = io_i_branch_resolve_pack_taken & btb_215_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_215_bht_T_4 = btb_215_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_215_bht_T_5 = io_i_branch_resolve_pack_taken & btb_215_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_215_bht_T_6 = btb_215_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_215_bht_T_7 = io_i_branch_resolve_pack_taken & btb_215_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_215_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_215_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_215_bht_T_13 = _btb_0_bht_T_8 & _btb_215_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_215_bht_T_16 = _btb_0_bht_T_8 & _btb_215_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_215_bht_T_19 = _btb_0_bht_T_8 & _btb_215_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_215_bht_T_20 = _btb_215_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_21 = _btb_215_bht_T_16 ? 2'h0 : _btb_215_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_22 = _btb_215_bht_T_13 ? 2'h0 : _btb_215_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_23 = _btb_215_bht_T_10 ? 2'h0 : _btb_215_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_24 = _btb_215_bht_T_7 ? 2'h3 : _btb_215_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_25 = _btb_215_bht_T_5 ? 2'h3 : _btb_215_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_26 = _btb_215_bht_T_3 ? 2'h3 : _btb_215_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_215_bht_T_27 = _btb_215_bht_T_1 ? 2'h1 : _btb_215_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9566 = btb_215_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6871
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9568 = btb_215_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_215_bht_T_27 : _GEN_8407; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_216_bht_T = btb_216_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_216_bht_T_1 = io_i_branch_resolve_pack_taken & btb_216_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_216_bht_T_2 = btb_216_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_216_bht_T_3 = io_i_branch_resolve_pack_taken & btb_216_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_216_bht_T_4 = btb_216_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_216_bht_T_5 = io_i_branch_resolve_pack_taken & btb_216_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_216_bht_T_6 = btb_216_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_216_bht_T_7 = io_i_branch_resolve_pack_taken & btb_216_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_216_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_216_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_216_bht_T_13 = _btb_0_bht_T_8 & _btb_216_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_216_bht_T_16 = _btb_0_bht_T_8 & _btb_216_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_216_bht_T_19 = _btb_0_bht_T_8 & _btb_216_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_216_bht_T_20 = _btb_216_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_21 = _btb_216_bht_T_16 ? 2'h0 : _btb_216_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_22 = _btb_216_bht_T_13 ? 2'h0 : _btb_216_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_23 = _btb_216_bht_T_10 ? 2'h0 : _btb_216_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_24 = _btb_216_bht_T_7 ? 2'h3 : _btb_216_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_25 = _btb_216_bht_T_5 ? 2'h3 : _btb_216_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_26 = _btb_216_bht_T_3 ? 2'h3 : _btb_216_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_216_bht_T_27 = _btb_216_bht_T_1 ? 2'h1 : _btb_216_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9570 = btb_216_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6872
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9572 = btb_216_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_216_bht_T_27 : _GEN_8408; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_217_bht_T = btb_217_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_217_bht_T_1 = io_i_branch_resolve_pack_taken & btb_217_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_217_bht_T_2 = btb_217_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_217_bht_T_3 = io_i_branch_resolve_pack_taken & btb_217_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_217_bht_T_4 = btb_217_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_217_bht_T_5 = io_i_branch_resolve_pack_taken & btb_217_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_217_bht_T_6 = btb_217_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_217_bht_T_7 = io_i_branch_resolve_pack_taken & btb_217_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_217_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_217_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_217_bht_T_13 = _btb_0_bht_T_8 & _btb_217_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_217_bht_T_16 = _btb_0_bht_T_8 & _btb_217_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_217_bht_T_19 = _btb_0_bht_T_8 & _btb_217_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_217_bht_T_20 = _btb_217_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_21 = _btb_217_bht_T_16 ? 2'h0 : _btb_217_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_22 = _btb_217_bht_T_13 ? 2'h0 : _btb_217_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_23 = _btb_217_bht_T_10 ? 2'h0 : _btb_217_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_24 = _btb_217_bht_T_7 ? 2'h3 : _btb_217_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_25 = _btb_217_bht_T_5 ? 2'h3 : _btb_217_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_26 = _btb_217_bht_T_3 ? 2'h3 : _btb_217_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_217_bht_T_27 = _btb_217_bht_T_1 ? 2'h1 : _btb_217_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9574 = btb_217_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6873
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9576 = btb_217_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_217_bht_T_27 : _GEN_8409; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_218_bht_T = btb_218_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_218_bht_T_1 = io_i_branch_resolve_pack_taken & btb_218_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_218_bht_T_2 = btb_218_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_218_bht_T_3 = io_i_branch_resolve_pack_taken & btb_218_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_218_bht_T_4 = btb_218_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_218_bht_T_5 = io_i_branch_resolve_pack_taken & btb_218_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_218_bht_T_6 = btb_218_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_218_bht_T_7 = io_i_branch_resolve_pack_taken & btb_218_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_218_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_218_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_218_bht_T_13 = _btb_0_bht_T_8 & _btb_218_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_218_bht_T_16 = _btb_0_bht_T_8 & _btb_218_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_218_bht_T_19 = _btb_0_bht_T_8 & _btb_218_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_218_bht_T_20 = _btb_218_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_21 = _btb_218_bht_T_16 ? 2'h0 : _btb_218_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_22 = _btb_218_bht_T_13 ? 2'h0 : _btb_218_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_23 = _btb_218_bht_T_10 ? 2'h0 : _btb_218_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_24 = _btb_218_bht_T_7 ? 2'h3 : _btb_218_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_25 = _btb_218_bht_T_5 ? 2'h3 : _btb_218_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_26 = _btb_218_bht_T_3 ? 2'h3 : _btb_218_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_218_bht_T_27 = _btb_218_bht_T_1 ? 2'h1 : _btb_218_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9578 = btb_218_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6874
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9580 = btb_218_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_218_bht_T_27 : _GEN_8410; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_219_bht_T = btb_219_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_219_bht_T_1 = io_i_branch_resolve_pack_taken & btb_219_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_219_bht_T_2 = btb_219_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_219_bht_T_3 = io_i_branch_resolve_pack_taken & btb_219_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_219_bht_T_4 = btb_219_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_219_bht_T_5 = io_i_branch_resolve_pack_taken & btb_219_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_219_bht_T_6 = btb_219_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_219_bht_T_7 = io_i_branch_resolve_pack_taken & btb_219_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_219_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_219_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_219_bht_T_13 = _btb_0_bht_T_8 & _btb_219_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_219_bht_T_16 = _btb_0_bht_T_8 & _btb_219_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_219_bht_T_19 = _btb_0_bht_T_8 & _btb_219_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_219_bht_T_20 = _btb_219_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_21 = _btb_219_bht_T_16 ? 2'h0 : _btb_219_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_22 = _btb_219_bht_T_13 ? 2'h0 : _btb_219_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_23 = _btb_219_bht_T_10 ? 2'h0 : _btb_219_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_24 = _btb_219_bht_T_7 ? 2'h3 : _btb_219_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_25 = _btb_219_bht_T_5 ? 2'h3 : _btb_219_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_26 = _btb_219_bht_T_3 ? 2'h3 : _btb_219_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_219_bht_T_27 = _btb_219_bht_T_1 ? 2'h1 : _btb_219_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9582 = btb_219_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6875
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9584 = btb_219_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_219_bht_T_27 : _GEN_8411; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_220_bht_T = btb_220_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_220_bht_T_1 = io_i_branch_resolve_pack_taken & btb_220_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_220_bht_T_2 = btb_220_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_220_bht_T_3 = io_i_branch_resolve_pack_taken & btb_220_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_220_bht_T_4 = btb_220_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_220_bht_T_5 = io_i_branch_resolve_pack_taken & btb_220_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_220_bht_T_6 = btb_220_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_220_bht_T_7 = io_i_branch_resolve_pack_taken & btb_220_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_220_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_220_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_220_bht_T_13 = _btb_0_bht_T_8 & _btb_220_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_220_bht_T_16 = _btb_0_bht_T_8 & _btb_220_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_220_bht_T_19 = _btb_0_bht_T_8 & _btb_220_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_220_bht_T_20 = _btb_220_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_21 = _btb_220_bht_T_16 ? 2'h0 : _btb_220_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_22 = _btb_220_bht_T_13 ? 2'h0 : _btb_220_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_23 = _btb_220_bht_T_10 ? 2'h0 : _btb_220_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_24 = _btb_220_bht_T_7 ? 2'h3 : _btb_220_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_25 = _btb_220_bht_T_5 ? 2'h3 : _btb_220_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_26 = _btb_220_bht_T_3 ? 2'h3 : _btb_220_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_220_bht_T_27 = _btb_220_bht_T_1 ? 2'h1 : _btb_220_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9586 = btb_220_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6876
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9588 = btb_220_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_220_bht_T_27 : _GEN_8412; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_221_bht_T = btb_221_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_221_bht_T_1 = io_i_branch_resolve_pack_taken & btb_221_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_221_bht_T_2 = btb_221_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_221_bht_T_3 = io_i_branch_resolve_pack_taken & btb_221_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_221_bht_T_4 = btb_221_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_221_bht_T_5 = io_i_branch_resolve_pack_taken & btb_221_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_221_bht_T_6 = btb_221_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_221_bht_T_7 = io_i_branch_resolve_pack_taken & btb_221_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_221_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_221_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_221_bht_T_13 = _btb_0_bht_T_8 & _btb_221_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_221_bht_T_16 = _btb_0_bht_T_8 & _btb_221_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_221_bht_T_19 = _btb_0_bht_T_8 & _btb_221_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_221_bht_T_20 = _btb_221_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_21 = _btb_221_bht_T_16 ? 2'h0 : _btb_221_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_22 = _btb_221_bht_T_13 ? 2'h0 : _btb_221_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_23 = _btb_221_bht_T_10 ? 2'h0 : _btb_221_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_24 = _btb_221_bht_T_7 ? 2'h3 : _btb_221_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_25 = _btb_221_bht_T_5 ? 2'h3 : _btb_221_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_26 = _btb_221_bht_T_3 ? 2'h3 : _btb_221_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_221_bht_T_27 = _btb_221_bht_T_1 ? 2'h1 : _btb_221_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9590 = btb_221_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6877
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9592 = btb_221_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_221_bht_T_27 : _GEN_8413; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_222_bht_T = btb_222_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_222_bht_T_1 = io_i_branch_resolve_pack_taken & btb_222_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_222_bht_T_2 = btb_222_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_222_bht_T_3 = io_i_branch_resolve_pack_taken & btb_222_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_222_bht_T_4 = btb_222_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_222_bht_T_5 = io_i_branch_resolve_pack_taken & btb_222_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_222_bht_T_6 = btb_222_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_222_bht_T_7 = io_i_branch_resolve_pack_taken & btb_222_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_222_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_222_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_222_bht_T_13 = _btb_0_bht_T_8 & _btb_222_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_222_bht_T_16 = _btb_0_bht_T_8 & _btb_222_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_222_bht_T_19 = _btb_0_bht_T_8 & _btb_222_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_222_bht_T_20 = _btb_222_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_21 = _btb_222_bht_T_16 ? 2'h0 : _btb_222_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_22 = _btb_222_bht_T_13 ? 2'h0 : _btb_222_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_23 = _btb_222_bht_T_10 ? 2'h0 : _btb_222_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_24 = _btb_222_bht_T_7 ? 2'h3 : _btb_222_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_25 = _btb_222_bht_T_5 ? 2'h3 : _btb_222_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_26 = _btb_222_bht_T_3 ? 2'h3 : _btb_222_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_222_bht_T_27 = _btb_222_bht_T_1 ? 2'h1 : _btb_222_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9594 = btb_222_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6878
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9596 = btb_222_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_222_bht_T_27 : _GEN_8414; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_223_bht_T = btb_223_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_223_bht_T_1 = io_i_branch_resolve_pack_taken & btb_223_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_223_bht_T_2 = btb_223_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_223_bht_T_3 = io_i_branch_resolve_pack_taken & btb_223_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_223_bht_T_4 = btb_223_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_223_bht_T_5 = io_i_branch_resolve_pack_taken & btb_223_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_223_bht_T_6 = btb_223_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_223_bht_T_7 = io_i_branch_resolve_pack_taken & btb_223_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_223_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_223_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_223_bht_T_13 = _btb_0_bht_T_8 & _btb_223_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_223_bht_T_16 = _btb_0_bht_T_8 & _btb_223_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_223_bht_T_19 = _btb_0_bht_T_8 & _btb_223_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_223_bht_T_20 = _btb_223_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_21 = _btb_223_bht_T_16 ? 2'h0 : _btb_223_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_22 = _btb_223_bht_T_13 ? 2'h0 : _btb_223_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_23 = _btb_223_bht_T_10 ? 2'h0 : _btb_223_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_24 = _btb_223_bht_T_7 ? 2'h3 : _btb_223_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_25 = _btb_223_bht_T_5 ? 2'h3 : _btb_223_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_26 = _btb_223_bht_T_3 ? 2'h3 : _btb_223_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_223_bht_T_27 = _btb_223_bht_T_1 ? 2'h1 : _btb_223_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9598 = btb_223_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6879
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9600 = btb_223_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_223_bht_T_27 : _GEN_8415; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_224_bht_T = btb_224_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_224_bht_T_1 = io_i_branch_resolve_pack_taken & btb_224_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_224_bht_T_2 = btb_224_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_224_bht_T_3 = io_i_branch_resolve_pack_taken & btb_224_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_224_bht_T_4 = btb_224_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_224_bht_T_5 = io_i_branch_resolve_pack_taken & btb_224_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_224_bht_T_6 = btb_224_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_224_bht_T_7 = io_i_branch_resolve_pack_taken & btb_224_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_224_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_224_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_224_bht_T_13 = _btb_0_bht_T_8 & _btb_224_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_224_bht_T_16 = _btb_0_bht_T_8 & _btb_224_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_224_bht_T_19 = _btb_0_bht_T_8 & _btb_224_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_224_bht_T_20 = _btb_224_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_21 = _btb_224_bht_T_16 ? 2'h0 : _btb_224_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_22 = _btb_224_bht_T_13 ? 2'h0 : _btb_224_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_23 = _btb_224_bht_T_10 ? 2'h0 : _btb_224_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_24 = _btb_224_bht_T_7 ? 2'h3 : _btb_224_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_25 = _btb_224_bht_T_5 ? 2'h3 : _btb_224_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_26 = _btb_224_bht_T_3 ? 2'h3 : _btb_224_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_224_bht_T_27 = _btb_224_bht_T_1 ? 2'h1 : _btb_224_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9601 = btb_224_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_223_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_222_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_221_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_220_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_219_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_218_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_217_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_216_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_215_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_214_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_213_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_212_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_211_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_210_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9541)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9602 = btb_224_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6880
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9604 = btb_224_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_224_bht_T_27 : _GEN_8416; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_225_bht_T = btb_225_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_225_bht_T_1 = io_i_branch_resolve_pack_taken & btb_225_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_225_bht_T_2 = btb_225_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_225_bht_T_3 = io_i_branch_resolve_pack_taken & btb_225_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_225_bht_T_4 = btb_225_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_225_bht_T_5 = io_i_branch_resolve_pack_taken & btb_225_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_225_bht_T_6 = btb_225_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_225_bht_T_7 = io_i_branch_resolve_pack_taken & btb_225_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_225_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_225_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_225_bht_T_13 = _btb_0_bht_T_8 & _btb_225_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_225_bht_T_16 = _btb_0_bht_T_8 & _btb_225_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_225_bht_T_19 = _btb_0_bht_T_8 & _btb_225_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_225_bht_T_20 = _btb_225_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_21 = _btb_225_bht_T_16 ? 2'h0 : _btb_225_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_22 = _btb_225_bht_T_13 ? 2'h0 : _btb_225_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_23 = _btb_225_bht_T_10 ? 2'h0 : _btb_225_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_24 = _btb_225_bht_T_7 ? 2'h3 : _btb_225_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_25 = _btb_225_bht_T_5 ? 2'h3 : _btb_225_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_26 = _btb_225_bht_T_3 ? 2'h3 : _btb_225_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_225_bht_T_27 = _btb_225_bht_T_1 ? 2'h1 : _btb_225_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9606 = btb_225_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6881
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9608 = btb_225_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_225_bht_T_27 : _GEN_8417; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_226_bht_T = btb_226_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_226_bht_T_1 = io_i_branch_resolve_pack_taken & btb_226_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_226_bht_T_2 = btb_226_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_226_bht_T_3 = io_i_branch_resolve_pack_taken & btb_226_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_226_bht_T_4 = btb_226_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_226_bht_T_5 = io_i_branch_resolve_pack_taken & btb_226_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_226_bht_T_6 = btb_226_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_226_bht_T_7 = io_i_branch_resolve_pack_taken & btb_226_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_226_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_226_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_226_bht_T_13 = _btb_0_bht_T_8 & _btb_226_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_226_bht_T_16 = _btb_0_bht_T_8 & _btb_226_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_226_bht_T_19 = _btb_0_bht_T_8 & _btb_226_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_226_bht_T_20 = _btb_226_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_21 = _btb_226_bht_T_16 ? 2'h0 : _btb_226_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_22 = _btb_226_bht_T_13 ? 2'h0 : _btb_226_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_23 = _btb_226_bht_T_10 ? 2'h0 : _btb_226_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_24 = _btb_226_bht_T_7 ? 2'h3 : _btb_226_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_25 = _btb_226_bht_T_5 ? 2'h3 : _btb_226_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_26 = _btb_226_bht_T_3 ? 2'h3 : _btb_226_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_226_bht_T_27 = _btb_226_bht_T_1 ? 2'h1 : _btb_226_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9610 = btb_226_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6882
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9612 = btb_226_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_226_bht_T_27 : _GEN_8418; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_227_bht_T = btb_227_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_227_bht_T_1 = io_i_branch_resolve_pack_taken & btb_227_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_227_bht_T_2 = btb_227_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_227_bht_T_3 = io_i_branch_resolve_pack_taken & btb_227_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_227_bht_T_4 = btb_227_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_227_bht_T_5 = io_i_branch_resolve_pack_taken & btb_227_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_227_bht_T_6 = btb_227_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_227_bht_T_7 = io_i_branch_resolve_pack_taken & btb_227_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_227_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_227_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_227_bht_T_13 = _btb_0_bht_T_8 & _btb_227_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_227_bht_T_16 = _btb_0_bht_T_8 & _btb_227_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_227_bht_T_19 = _btb_0_bht_T_8 & _btb_227_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_227_bht_T_20 = _btb_227_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_21 = _btb_227_bht_T_16 ? 2'h0 : _btb_227_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_22 = _btb_227_bht_T_13 ? 2'h0 : _btb_227_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_23 = _btb_227_bht_T_10 ? 2'h0 : _btb_227_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_24 = _btb_227_bht_T_7 ? 2'h3 : _btb_227_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_25 = _btb_227_bht_T_5 ? 2'h3 : _btb_227_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_26 = _btb_227_bht_T_3 ? 2'h3 : _btb_227_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_227_bht_T_27 = _btb_227_bht_T_1 ? 2'h1 : _btb_227_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9614 = btb_227_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6883
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9616 = btb_227_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_227_bht_T_27 : _GEN_8419; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_228_bht_T = btb_228_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_228_bht_T_1 = io_i_branch_resolve_pack_taken & btb_228_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_228_bht_T_2 = btb_228_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_228_bht_T_3 = io_i_branch_resolve_pack_taken & btb_228_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_228_bht_T_4 = btb_228_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_228_bht_T_5 = io_i_branch_resolve_pack_taken & btb_228_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_228_bht_T_6 = btb_228_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_228_bht_T_7 = io_i_branch_resolve_pack_taken & btb_228_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_228_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_228_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_228_bht_T_13 = _btb_0_bht_T_8 & _btb_228_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_228_bht_T_16 = _btb_0_bht_T_8 & _btb_228_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_228_bht_T_19 = _btb_0_bht_T_8 & _btb_228_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_228_bht_T_20 = _btb_228_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_21 = _btb_228_bht_T_16 ? 2'h0 : _btb_228_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_22 = _btb_228_bht_T_13 ? 2'h0 : _btb_228_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_23 = _btb_228_bht_T_10 ? 2'h0 : _btb_228_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_24 = _btb_228_bht_T_7 ? 2'h3 : _btb_228_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_25 = _btb_228_bht_T_5 ? 2'h3 : _btb_228_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_26 = _btb_228_bht_T_3 ? 2'h3 : _btb_228_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_228_bht_T_27 = _btb_228_bht_T_1 ? 2'h1 : _btb_228_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9618 = btb_228_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6884
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9620 = btb_228_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_228_bht_T_27 : _GEN_8420; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_229_bht_T = btb_229_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_229_bht_T_1 = io_i_branch_resolve_pack_taken & btb_229_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_229_bht_T_2 = btb_229_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_229_bht_T_3 = io_i_branch_resolve_pack_taken & btb_229_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_229_bht_T_4 = btb_229_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_229_bht_T_5 = io_i_branch_resolve_pack_taken & btb_229_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_229_bht_T_6 = btb_229_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_229_bht_T_7 = io_i_branch_resolve_pack_taken & btb_229_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_229_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_229_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_229_bht_T_13 = _btb_0_bht_T_8 & _btb_229_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_229_bht_T_16 = _btb_0_bht_T_8 & _btb_229_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_229_bht_T_19 = _btb_0_bht_T_8 & _btb_229_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_229_bht_T_20 = _btb_229_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_21 = _btb_229_bht_T_16 ? 2'h0 : _btb_229_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_22 = _btb_229_bht_T_13 ? 2'h0 : _btb_229_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_23 = _btb_229_bht_T_10 ? 2'h0 : _btb_229_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_24 = _btb_229_bht_T_7 ? 2'h3 : _btb_229_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_25 = _btb_229_bht_T_5 ? 2'h3 : _btb_229_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_26 = _btb_229_bht_T_3 ? 2'h3 : _btb_229_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_229_bht_T_27 = _btb_229_bht_T_1 ? 2'h1 : _btb_229_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9622 = btb_229_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6885
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9624 = btb_229_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_229_bht_T_27 : _GEN_8421; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_230_bht_T = btb_230_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_230_bht_T_1 = io_i_branch_resolve_pack_taken & btb_230_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_230_bht_T_2 = btb_230_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_230_bht_T_3 = io_i_branch_resolve_pack_taken & btb_230_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_230_bht_T_4 = btb_230_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_230_bht_T_5 = io_i_branch_resolve_pack_taken & btb_230_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_230_bht_T_6 = btb_230_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_230_bht_T_7 = io_i_branch_resolve_pack_taken & btb_230_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_230_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_230_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_230_bht_T_13 = _btb_0_bht_T_8 & _btb_230_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_230_bht_T_16 = _btb_0_bht_T_8 & _btb_230_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_230_bht_T_19 = _btb_0_bht_T_8 & _btb_230_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_230_bht_T_20 = _btb_230_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_21 = _btb_230_bht_T_16 ? 2'h0 : _btb_230_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_22 = _btb_230_bht_T_13 ? 2'h0 : _btb_230_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_23 = _btb_230_bht_T_10 ? 2'h0 : _btb_230_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_24 = _btb_230_bht_T_7 ? 2'h3 : _btb_230_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_25 = _btb_230_bht_T_5 ? 2'h3 : _btb_230_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_26 = _btb_230_bht_T_3 ? 2'h3 : _btb_230_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_230_bht_T_27 = _btb_230_bht_T_1 ? 2'h1 : _btb_230_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9626 = btb_230_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6886
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9628 = btb_230_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_230_bht_T_27 : _GEN_8422; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_231_bht_T = btb_231_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_231_bht_T_1 = io_i_branch_resolve_pack_taken & btb_231_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_231_bht_T_2 = btb_231_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_231_bht_T_3 = io_i_branch_resolve_pack_taken & btb_231_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_231_bht_T_4 = btb_231_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_231_bht_T_5 = io_i_branch_resolve_pack_taken & btb_231_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_231_bht_T_6 = btb_231_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_231_bht_T_7 = io_i_branch_resolve_pack_taken & btb_231_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_231_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_231_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_231_bht_T_13 = _btb_0_bht_T_8 & _btb_231_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_231_bht_T_16 = _btb_0_bht_T_8 & _btb_231_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_231_bht_T_19 = _btb_0_bht_T_8 & _btb_231_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_231_bht_T_20 = _btb_231_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_21 = _btb_231_bht_T_16 ? 2'h0 : _btb_231_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_22 = _btb_231_bht_T_13 ? 2'h0 : _btb_231_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_23 = _btb_231_bht_T_10 ? 2'h0 : _btb_231_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_24 = _btb_231_bht_T_7 ? 2'h3 : _btb_231_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_25 = _btb_231_bht_T_5 ? 2'h3 : _btb_231_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_26 = _btb_231_bht_T_3 ? 2'h3 : _btb_231_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_231_bht_T_27 = _btb_231_bht_T_1 ? 2'h1 : _btb_231_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9630 = btb_231_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6887
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9632 = btb_231_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_231_bht_T_27 : _GEN_8423; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_232_bht_T = btb_232_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_232_bht_T_1 = io_i_branch_resolve_pack_taken & btb_232_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_232_bht_T_2 = btb_232_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_232_bht_T_3 = io_i_branch_resolve_pack_taken & btb_232_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_232_bht_T_4 = btb_232_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_232_bht_T_5 = io_i_branch_resolve_pack_taken & btb_232_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_232_bht_T_6 = btb_232_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_232_bht_T_7 = io_i_branch_resolve_pack_taken & btb_232_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_232_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_232_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_232_bht_T_13 = _btb_0_bht_T_8 & _btb_232_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_232_bht_T_16 = _btb_0_bht_T_8 & _btb_232_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_232_bht_T_19 = _btb_0_bht_T_8 & _btb_232_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_232_bht_T_20 = _btb_232_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_21 = _btb_232_bht_T_16 ? 2'h0 : _btb_232_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_22 = _btb_232_bht_T_13 ? 2'h0 : _btb_232_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_23 = _btb_232_bht_T_10 ? 2'h0 : _btb_232_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_24 = _btb_232_bht_T_7 ? 2'h3 : _btb_232_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_25 = _btb_232_bht_T_5 ? 2'h3 : _btb_232_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_26 = _btb_232_bht_T_3 ? 2'h3 : _btb_232_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_232_bht_T_27 = _btb_232_bht_T_1 ? 2'h1 : _btb_232_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9634 = btb_232_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6888
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9636 = btb_232_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_232_bht_T_27 : _GEN_8424; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_233_bht_T = btb_233_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_233_bht_T_1 = io_i_branch_resolve_pack_taken & btb_233_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_233_bht_T_2 = btb_233_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_233_bht_T_3 = io_i_branch_resolve_pack_taken & btb_233_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_233_bht_T_4 = btb_233_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_233_bht_T_5 = io_i_branch_resolve_pack_taken & btb_233_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_233_bht_T_6 = btb_233_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_233_bht_T_7 = io_i_branch_resolve_pack_taken & btb_233_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_233_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_233_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_233_bht_T_13 = _btb_0_bht_T_8 & _btb_233_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_233_bht_T_16 = _btb_0_bht_T_8 & _btb_233_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_233_bht_T_19 = _btb_0_bht_T_8 & _btb_233_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_233_bht_T_20 = _btb_233_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_21 = _btb_233_bht_T_16 ? 2'h0 : _btb_233_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_22 = _btb_233_bht_T_13 ? 2'h0 : _btb_233_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_23 = _btb_233_bht_T_10 ? 2'h0 : _btb_233_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_24 = _btb_233_bht_T_7 ? 2'h3 : _btb_233_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_25 = _btb_233_bht_T_5 ? 2'h3 : _btb_233_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_26 = _btb_233_bht_T_3 ? 2'h3 : _btb_233_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_233_bht_T_27 = _btb_233_bht_T_1 ? 2'h1 : _btb_233_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9638 = btb_233_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6889
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9640 = btb_233_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_233_bht_T_27 : _GEN_8425; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_234_bht_T = btb_234_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_234_bht_T_1 = io_i_branch_resolve_pack_taken & btb_234_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_234_bht_T_2 = btb_234_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_234_bht_T_3 = io_i_branch_resolve_pack_taken & btb_234_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_234_bht_T_4 = btb_234_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_234_bht_T_5 = io_i_branch_resolve_pack_taken & btb_234_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_234_bht_T_6 = btb_234_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_234_bht_T_7 = io_i_branch_resolve_pack_taken & btb_234_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_234_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_234_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_234_bht_T_13 = _btb_0_bht_T_8 & _btb_234_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_234_bht_T_16 = _btb_0_bht_T_8 & _btb_234_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_234_bht_T_19 = _btb_0_bht_T_8 & _btb_234_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_234_bht_T_20 = _btb_234_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_21 = _btb_234_bht_T_16 ? 2'h0 : _btb_234_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_22 = _btb_234_bht_T_13 ? 2'h0 : _btb_234_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_23 = _btb_234_bht_T_10 ? 2'h0 : _btb_234_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_24 = _btb_234_bht_T_7 ? 2'h3 : _btb_234_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_25 = _btb_234_bht_T_5 ? 2'h3 : _btb_234_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_26 = _btb_234_bht_T_3 ? 2'h3 : _btb_234_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_234_bht_T_27 = _btb_234_bht_T_1 ? 2'h1 : _btb_234_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9642 = btb_234_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6890
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9644 = btb_234_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_234_bht_T_27 : _GEN_8426; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_235_bht_T = btb_235_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_235_bht_T_1 = io_i_branch_resolve_pack_taken & btb_235_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_235_bht_T_2 = btb_235_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_235_bht_T_3 = io_i_branch_resolve_pack_taken & btb_235_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_235_bht_T_4 = btb_235_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_235_bht_T_5 = io_i_branch_resolve_pack_taken & btb_235_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_235_bht_T_6 = btb_235_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_235_bht_T_7 = io_i_branch_resolve_pack_taken & btb_235_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_235_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_235_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_235_bht_T_13 = _btb_0_bht_T_8 & _btb_235_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_235_bht_T_16 = _btb_0_bht_T_8 & _btb_235_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_235_bht_T_19 = _btb_0_bht_T_8 & _btb_235_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_235_bht_T_20 = _btb_235_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_21 = _btb_235_bht_T_16 ? 2'h0 : _btb_235_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_22 = _btb_235_bht_T_13 ? 2'h0 : _btb_235_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_23 = _btb_235_bht_T_10 ? 2'h0 : _btb_235_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_24 = _btb_235_bht_T_7 ? 2'h3 : _btb_235_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_25 = _btb_235_bht_T_5 ? 2'h3 : _btb_235_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_26 = _btb_235_bht_T_3 ? 2'h3 : _btb_235_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_235_bht_T_27 = _btb_235_bht_T_1 ? 2'h1 : _btb_235_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9646 = btb_235_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6891
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9648 = btb_235_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_235_bht_T_27 : _GEN_8427; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_236_bht_T = btb_236_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_236_bht_T_1 = io_i_branch_resolve_pack_taken & btb_236_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_236_bht_T_2 = btb_236_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_236_bht_T_3 = io_i_branch_resolve_pack_taken & btb_236_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_236_bht_T_4 = btb_236_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_236_bht_T_5 = io_i_branch_resolve_pack_taken & btb_236_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_236_bht_T_6 = btb_236_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_236_bht_T_7 = io_i_branch_resolve_pack_taken & btb_236_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_236_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_236_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_236_bht_T_13 = _btb_0_bht_T_8 & _btb_236_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_236_bht_T_16 = _btb_0_bht_T_8 & _btb_236_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_236_bht_T_19 = _btb_0_bht_T_8 & _btb_236_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_236_bht_T_20 = _btb_236_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_21 = _btb_236_bht_T_16 ? 2'h0 : _btb_236_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_22 = _btb_236_bht_T_13 ? 2'h0 : _btb_236_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_23 = _btb_236_bht_T_10 ? 2'h0 : _btb_236_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_24 = _btb_236_bht_T_7 ? 2'h3 : _btb_236_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_25 = _btb_236_bht_T_5 ? 2'h3 : _btb_236_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_26 = _btb_236_bht_T_3 ? 2'h3 : _btb_236_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_236_bht_T_27 = _btb_236_bht_T_1 ? 2'h1 : _btb_236_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9650 = btb_236_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6892
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9652 = btb_236_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_236_bht_T_27 : _GEN_8428; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_237_bht_T = btb_237_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_237_bht_T_1 = io_i_branch_resolve_pack_taken & btb_237_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_237_bht_T_2 = btb_237_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_237_bht_T_3 = io_i_branch_resolve_pack_taken & btb_237_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_237_bht_T_4 = btb_237_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_237_bht_T_5 = io_i_branch_resolve_pack_taken & btb_237_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_237_bht_T_6 = btb_237_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_237_bht_T_7 = io_i_branch_resolve_pack_taken & btb_237_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_237_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_237_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_237_bht_T_13 = _btb_0_bht_T_8 & _btb_237_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_237_bht_T_16 = _btb_0_bht_T_8 & _btb_237_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_237_bht_T_19 = _btb_0_bht_T_8 & _btb_237_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_237_bht_T_20 = _btb_237_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_21 = _btb_237_bht_T_16 ? 2'h0 : _btb_237_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_22 = _btb_237_bht_T_13 ? 2'h0 : _btb_237_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_23 = _btb_237_bht_T_10 ? 2'h0 : _btb_237_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_24 = _btb_237_bht_T_7 ? 2'h3 : _btb_237_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_25 = _btb_237_bht_T_5 ? 2'h3 : _btb_237_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_26 = _btb_237_bht_T_3 ? 2'h3 : _btb_237_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_237_bht_T_27 = _btb_237_bht_T_1 ? 2'h1 : _btb_237_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9654 = btb_237_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6893
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9656 = btb_237_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_237_bht_T_27 : _GEN_8429; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_238_bht_T = btb_238_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_238_bht_T_1 = io_i_branch_resolve_pack_taken & btb_238_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_238_bht_T_2 = btb_238_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_238_bht_T_3 = io_i_branch_resolve_pack_taken & btb_238_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_238_bht_T_4 = btb_238_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_238_bht_T_5 = io_i_branch_resolve_pack_taken & btb_238_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_238_bht_T_6 = btb_238_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_238_bht_T_7 = io_i_branch_resolve_pack_taken & btb_238_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_238_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_238_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_238_bht_T_13 = _btb_0_bht_T_8 & _btb_238_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_238_bht_T_16 = _btb_0_bht_T_8 & _btb_238_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_238_bht_T_19 = _btb_0_bht_T_8 & _btb_238_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_238_bht_T_20 = _btb_238_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_21 = _btb_238_bht_T_16 ? 2'h0 : _btb_238_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_22 = _btb_238_bht_T_13 ? 2'h0 : _btb_238_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_23 = _btb_238_bht_T_10 ? 2'h0 : _btb_238_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_24 = _btb_238_bht_T_7 ? 2'h3 : _btb_238_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_25 = _btb_238_bht_T_5 ? 2'h3 : _btb_238_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_26 = _btb_238_bht_T_3 ? 2'h3 : _btb_238_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_238_bht_T_27 = _btb_238_bht_T_1 ? 2'h1 : _btb_238_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9658 = btb_238_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6894
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9660 = btb_238_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_238_bht_T_27 : _GEN_8430; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_239_bht_T = btb_239_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_239_bht_T_1 = io_i_branch_resolve_pack_taken & btb_239_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_239_bht_T_2 = btb_239_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_239_bht_T_3 = io_i_branch_resolve_pack_taken & btb_239_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_239_bht_T_4 = btb_239_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_239_bht_T_5 = io_i_branch_resolve_pack_taken & btb_239_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_239_bht_T_6 = btb_239_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_239_bht_T_7 = io_i_branch_resolve_pack_taken & btb_239_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_239_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_239_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_239_bht_T_13 = _btb_0_bht_T_8 & _btb_239_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_239_bht_T_16 = _btb_0_bht_T_8 & _btb_239_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_239_bht_T_19 = _btb_0_bht_T_8 & _btb_239_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_239_bht_T_20 = _btb_239_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_21 = _btb_239_bht_T_16 ? 2'h0 : _btb_239_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_22 = _btb_239_bht_T_13 ? 2'h0 : _btb_239_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_23 = _btb_239_bht_T_10 ? 2'h0 : _btb_239_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_24 = _btb_239_bht_T_7 ? 2'h3 : _btb_239_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_25 = _btb_239_bht_T_5 ? 2'h3 : _btb_239_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_26 = _btb_239_bht_T_3 ? 2'h3 : _btb_239_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_239_bht_T_27 = _btb_239_bht_T_1 ? 2'h1 : _btb_239_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9661 = btb_239_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_238_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_237_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_236_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_235_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_234_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_233_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_232_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_231_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_230_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_229_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_228_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_227_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_226_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_225_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9601)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9662 = btb_239_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6895
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9664 = btb_239_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_239_bht_T_27 : _GEN_8431; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_240_bht_T = btb_240_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_240_bht_T_1 = io_i_branch_resolve_pack_taken & btb_240_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_240_bht_T_2 = btb_240_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_240_bht_T_3 = io_i_branch_resolve_pack_taken & btb_240_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_240_bht_T_4 = btb_240_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_240_bht_T_5 = io_i_branch_resolve_pack_taken & btb_240_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_240_bht_T_6 = btb_240_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_240_bht_T_7 = io_i_branch_resolve_pack_taken & btb_240_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_240_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_240_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_240_bht_T_13 = _btb_0_bht_T_8 & _btb_240_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_240_bht_T_16 = _btb_0_bht_T_8 & _btb_240_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_240_bht_T_19 = _btb_0_bht_T_8 & _btb_240_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_240_bht_T_20 = _btb_240_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_21 = _btb_240_bht_T_16 ? 2'h0 : _btb_240_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_22 = _btb_240_bht_T_13 ? 2'h0 : _btb_240_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_23 = _btb_240_bht_T_10 ? 2'h0 : _btb_240_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_24 = _btb_240_bht_T_7 ? 2'h3 : _btb_240_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_25 = _btb_240_bht_T_5 ? 2'h3 : _btb_240_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_26 = _btb_240_bht_T_3 ? 2'h3 : _btb_240_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_240_bht_T_27 = _btb_240_bht_T_1 ? 2'h1 : _btb_240_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9666 = btb_240_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6896
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9668 = btb_240_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_240_bht_T_27 : _GEN_8432; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_241_bht_T = btb_241_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_241_bht_T_1 = io_i_branch_resolve_pack_taken & btb_241_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_241_bht_T_2 = btb_241_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_241_bht_T_3 = io_i_branch_resolve_pack_taken & btb_241_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_241_bht_T_4 = btb_241_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_241_bht_T_5 = io_i_branch_resolve_pack_taken & btb_241_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_241_bht_T_6 = btb_241_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_241_bht_T_7 = io_i_branch_resolve_pack_taken & btb_241_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_241_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_241_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_241_bht_T_13 = _btb_0_bht_T_8 & _btb_241_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_241_bht_T_16 = _btb_0_bht_T_8 & _btb_241_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_241_bht_T_19 = _btb_0_bht_T_8 & _btb_241_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_241_bht_T_20 = _btb_241_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_21 = _btb_241_bht_T_16 ? 2'h0 : _btb_241_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_22 = _btb_241_bht_T_13 ? 2'h0 : _btb_241_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_23 = _btb_241_bht_T_10 ? 2'h0 : _btb_241_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_24 = _btb_241_bht_T_7 ? 2'h3 : _btb_241_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_25 = _btb_241_bht_T_5 ? 2'h3 : _btb_241_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_26 = _btb_241_bht_T_3 ? 2'h3 : _btb_241_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_241_bht_T_27 = _btb_241_bht_T_1 ? 2'h1 : _btb_241_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9670 = btb_241_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6897
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9672 = btb_241_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_241_bht_T_27 : _GEN_8433; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_242_bht_T = btb_242_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_242_bht_T_1 = io_i_branch_resolve_pack_taken & btb_242_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_242_bht_T_2 = btb_242_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_242_bht_T_3 = io_i_branch_resolve_pack_taken & btb_242_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_242_bht_T_4 = btb_242_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_242_bht_T_5 = io_i_branch_resolve_pack_taken & btb_242_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_242_bht_T_6 = btb_242_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_242_bht_T_7 = io_i_branch_resolve_pack_taken & btb_242_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_242_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_242_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_242_bht_T_13 = _btb_0_bht_T_8 & _btb_242_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_242_bht_T_16 = _btb_0_bht_T_8 & _btb_242_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_242_bht_T_19 = _btb_0_bht_T_8 & _btb_242_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_242_bht_T_20 = _btb_242_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_21 = _btb_242_bht_T_16 ? 2'h0 : _btb_242_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_22 = _btb_242_bht_T_13 ? 2'h0 : _btb_242_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_23 = _btb_242_bht_T_10 ? 2'h0 : _btb_242_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_24 = _btb_242_bht_T_7 ? 2'h3 : _btb_242_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_25 = _btb_242_bht_T_5 ? 2'h3 : _btb_242_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_26 = _btb_242_bht_T_3 ? 2'h3 : _btb_242_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_242_bht_T_27 = _btb_242_bht_T_1 ? 2'h1 : _btb_242_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9674 = btb_242_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6898
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9676 = btb_242_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_242_bht_T_27 : _GEN_8434; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_243_bht_T = btb_243_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_243_bht_T_1 = io_i_branch_resolve_pack_taken & btb_243_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_243_bht_T_2 = btb_243_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_243_bht_T_3 = io_i_branch_resolve_pack_taken & btb_243_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_243_bht_T_4 = btb_243_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_243_bht_T_5 = io_i_branch_resolve_pack_taken & btb_243_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_243_bht_T_6 = btb_243_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_243_bht_T_7 = io_i_branch_resolve_pack_taken & btb_243_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_243_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_243_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_243_bht_T_13 = _btb_0_bht_T_8 & _btb_243_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_243_bht_T_16 = _btb_0_bht_T_8 & _btb_243_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_243_bht_T_19 = _btb_0_bht_T_8 & _btb_243_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_243_bht_T_20 = _btb_243_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_21 = _btb_243_bht_T_16 ? 2'h0 : _btb_243_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_22 = _btb_243_bht_T_13 ? 2'h0 : _btb_243_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_23 = _btb_243_bht_T_10 ? 2'h0 : _btb_243_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_24 = _btb_243_bht_T_7 ? 2'h3 : _btb_243_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_25 = _btb_243_bht_T_5 ? 2'h3 : _btb_243_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_26 = _btb_243_bht_T_3 ? 2'h3 : _btb_243_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_243_bht_T_27 = _btb_243_bht_T_1 ? 2'h1 : _btb_243_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9678 = btb_243_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6899
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9680 = btb_243_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_243_bht_T_27 : _GEN_8435; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_244_bht_T = btb_244_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_244_bht_T_1 = io_i_branch_resolve_pack_taken & btb_244_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_244_bht_T_2 = btb_244_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_244_bht_T_3 = io_i_branch_resolve_pack_taken & btb_244_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_244_bht_T_4 = btb_244_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_244_bht_T_5 = io_i_branch_resolve_pack_taken & btb_244_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_244_bht_T_6 = btb_244_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_244_bht_T_7 = io_i_branch_resolve_pack_taken & btb_244_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_244_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_244_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_244_bht_T_13 = _btb_0_bht_T_8 & _btb_244_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_244_bht_T_16 = _btb_0_bht_T_8 & _btb_244_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_244_bht_T_19 = _btb_0_bht_T_8 & _btb_244_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_244_bht_T_20 = _btb_244_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_21 = _btb_244_bht_T_16 ? 2'h0 : _btb_244_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_22 = _btb_244_bht_T_13 ? 2'h0 : _btb_244_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_23 = _btb_244_bht_T_10 ? 2'h0 : _btb_244_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_24 = _btb_244_bht_T_7 ? 2'h3 : _btb_244_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_25 = _btb_244_bht_T_5 ? 2'h3 : _btb_244_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_26 = _btb_244_bht_T_3 ? 2'h3 : _btb_244_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_244_bht_T_27 = _btb_244_bht_T_1 ? 2'h1 : _btb_244_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9682 = btb_244_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6900
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9684 = btb_244_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_244_bht_T_27 : _GEN_8436; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_245_bht_T = btb_245_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_245_bht_T_1 = io_i_branch_resolve_pack_taken & btb_245_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_245_bht_T_2 = btb_245_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_245_bht_T_3 = io_i_branch_resolve_pack_taken & btb_245_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_245_bht_T_4 = btb_245_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_245_bht_T_5 = io_i_branch_resolve_pack_taken & btb_245_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_245_bht_T_6 = btb_245_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_245_bht_T_7 = io_i_branch_resolve_pack_taken & btb_245_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_245_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_245_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_245_bht_T_13 = _btb_0_bht_T_8 & _btb_245_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_245_bht_T_16 = _btb_0_bht_T_8 & _btb_245_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_245_bht_T_19 = _btb_0_bht_T_8 & _btb_245_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_245_bht_T_20 = _btb_245_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_21 = _btb_245_bht_T_16 ? 2'h0 : _btb_245_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_22 = _btb_245_bht_T_13 ? 2'h0 : _btb_245_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_23 = _btb_245_bht_T_10 ? 2'h0 : _btb_245_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_24 = _btb_245_bht_T_7 ? 2'h3 : _btb_245_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_25 = _btb_245_bht_T_5 ? 2'h3 : _btb_245_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_26 = _btb_245_bht_T_3 ? 2'h3 : _btb_245_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_245_bht_T_27 = _btb_245_bht_T_1 ? 2'h1 : _btb_245_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9686 = btb_245_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6901
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9688 = btb_245_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_245_bht_T_27 : _GEN_8437; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_246_bht_T = btb_246_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_246_bht_T_1 = io_i_branch_resolve_pack_taken & btb_246_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_246_bht_T_2 = btb_246_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_246_bht_T_3 = io_i_branch_resolve_pack_taken & btb_246_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_246_bht_T_4 = btb_246_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_246_bht_T_5 = io_i_branch_resolve_pack_taken & btb_246_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_246_bht_T_6 = btb_246_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_246_bht_T_7 = io_i_branch_resolve_pack_taken & btb_246_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_246_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_246_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_246_bht_T_13 = _btb_0_bht_T_8 & _btb_246_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_246_bht_T_16 = _btb_0_bht_T_8 & _btb_246_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_246_bht_T_19 = _btb_0_bht_T_8 & _btb_246_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_246_bht_T_20 = _btb_246_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_21 = _btb_246_bht_T_16 ? 2'h0 : _btb_246_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_22 = _btb_246_bht_T_13 ? 2'h0 : _btb_246_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_23 = _btb_246_bht_T_10 ? 2'h0 : _btb_246_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_24 = _btb_246_bht_T_7 ? 2'h3 : _btb_246_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_25 = _btb_246_bht_T_5 ? 2'h3 : _btb_246_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_26 = _btb_246_bht_T_3 ? 2'h3 : _btb_246_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_246_bht_T_27 = _btb_246_bht_T_1 ? 2'h1 : _btb_246_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9690 = btb_246_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6902
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9692 = btb_246_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_246_bht_T_27 : _GEN_8438; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_247_bht_T = btb_247_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_247_bht_T_1 = io_i_branch_resolve_pack_taken & btb_247_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_247_bht_T_2 = btb_247_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_247_bht_T_3 = io_i_branch_resolve_pack_taken & btb_247_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_247_bht_T_4 = btb_247_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_247_bht_T_5 = io_i_branch_resolve_pack_taken & btb_247_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_247_bht_T_6 = btb_247_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_247_bht_T_7 = io_i_branch_resolve_pack_taken & btb_247_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_247_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_247_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_247_bht_T_13 = _btb_0_bht_T_8 & _btb_247_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_247_bht_T_16 = _btb_0_bht_T_8 & _btb_247_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_247_bht_T_19 = _btb_0_bht_T_8 & _btb_247_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_247_bht_T_20 = _btb_247_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_21 = _btb_247_bht_T_16 ? 2'h0 : _btb_247_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_22 = _btb_247_bht_T_13 ? 2'h0 : _btb_247_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_23 = _btb_247_bht_T_10 ? 2'h0 : _btb_247_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_24 = _btb_247_bht_T_7 ? 2'h3 : _btb_247_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_25 = _btb_247_bht_T_5 ? 2'h3 : _btb_247_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_26 = _btb_247_bht_T_3 ? 2'h3 : _btb_247_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_247_bht_T_27 = _btb_247_bht_T_1 ? 2'h1 : _btb_247_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9694 = btb_247_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6903
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9696 = btb_247_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_247_bht_T_27 : _GEN_8439; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_248_bht_T = btb_248_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_248_bht_T_1 = io_i_branch_resolve_pack_taken & btb_248_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_248_bht_T_2 = btb_248_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_248_bht_T_3 = io_i_branch_resolve_pack_taken & btb_248_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_248_bht_T_4 = btb_248_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_248_bht_T_5 = io_i_branch_resolve_pack_taken & btb_248_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_248_bht_T_6 = btb_248_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_248_bht_T_7 = io_i_branch_resolve_pack_taken & btb_248_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_248_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_248_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_248_bht_T_13 = _btb_0_bht_T_8 & _btb_248_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_248_bht_T_16 = _btb_0_bht_T_8 & _btb_248_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_248_bht_T_19 = _btb_0_bht_T_8 & _btb_248_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_248_bht_T_20 = _btb_248_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_21 = _btb_248_bht_T_16 ? 2'h0 : _btb_248_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_22 = _btb_248_bht_T_13 ? 2'h0 : _btb_248_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_23 = _btb_248_bht_T_10 ? 2'h0 : _btb_248_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_24 = _btb_248_bht_T_7 ? 2'h3 : _btb_248_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_25 = _btb_248_bht_T_5 ? 2'h3 : _btb_248_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_26 = _btb_248_bht_T_3 ? 2'h3 : _btb_248_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_248_bht_T_27 = _btb_248_bht_T_1 ? 2'h1 : _btb_248_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9698 = btb_248_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6904
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9700 = btb_248_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_248_bht_T_27 : _GEN_8440; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_249_bht_T = btb_249_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_249_bht_T_1 = io_i_branch_resolve_pack_taken & btb_249_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_249_bht_T_2 = btb_249_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_249_bht_T_3 = io_i_branch_resolve_pack_taken & btb_249_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_249_bht_T_4 = btb_249_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_249_bht_T_5 = io_i_branch_resolve_pack_taken & btb_249_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_249_bht_T_6 = btb_249_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_249_bht_T_7 = io_i_branch_resolve_pack_taken & btb_249_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_249_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_249_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_249_bht_T_13 = _btb_0_bht_T_8 & _btb_249_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_249_bht_T_16 = _btb_0_bht_T_8 & _btb_249_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_249_bht_T_19 = _btb_0_bht_T_8 & _btb_249_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_249_bht_T_20 = _btb_249_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_21 = _btb_249_bht_T_16 ? 2'h0 : _btb_249_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_22 = _btb_249_bht_T_13 ? 2'h0 : _btb_249_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_23 = _btb_249_bht_T_10 ? 2'h0 : _btb_249_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_24 = _btb_249_bht_T_7 ? 2'h3 : _btb_249_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_25 = _btb_249_bht_T_5 ? 2'h3 : _btb_249_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_26 = _btb_249_bht_T_3 ? 2'h3 : _btb_249_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_249_bht_T_27 = _btb_249_bht_T_1 ? 2'h1 : _btb_249_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9702 = btb_249_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6905
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9704 = btb_249_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_249_bht_T_27 : _GEN_8441; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_250_bht_T = btb_250_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_250_bht_T_1 = io_i_branch_resolve_pack_taken & btb_250_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_250_bht_T_2 = btb_250_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_250_bht_T_3 = io_i_branch_resolve_pack_taken & btb_250_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_250_bht_T_4 = btb_250_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_250_bht_T_5 = io_i_branch_resolve_pack_taken & btb_250_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_250_bht_T_6 = btb_250_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_250_bht_T_7 = io_i_branch_resolve_pack_taken & btb_250_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_250_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_250_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_250_bht_T_13 = _btb_0_bht_T_8 & _btb_250_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_250_bht_T_16 = _btb_0_bht_T_8 & _btb_250_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_250_bht_T_19 = _btb_0_bht_T_8 & _btb_250_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_250_bht_T_20 = _btb_250_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_21 = _btb_250_bht_T_16 ? 2'h0 : _btb_250_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_22 = _btb_250_bht_T_13 ? 2'h0 : _btb_250_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_23 = _btb_250_bht_T_10 ? 2'h0 : _btb_250_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_24 = _btb_250_bht_T_7 ? 2'h3 : _btb_250_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_25 = _btb_250_bht_T_5 ? 2'h3 : _btb_250_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_26 = _btb_250_bht_T_3 ? 2'h3 : _btb_250_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_250_bht_T_27 = _btb_250_bht_T_1 ? 2'h1 : _btb_250_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9706 = btb_250_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6906
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9708 = btb_250_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_250_bht_T_27 : _GEN_8442; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_251_bht_T = btb_251_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_251_bht_T_1 = io_i_branch_resolve_pack_taken & btb_251_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_251_bht_T_2 = btb_251_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_251_bht_T_3 = io_i_branch_resolve_pack_taken & btb_251_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_251_bht_T_4 = btb_251_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_251_bht_T_5 = io_i_branch_resolve_pack_taken & btb_251_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_251_bht_T_6 = btb_251_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_251_bht_T_7 = io_i_branch_resolve_pack_taken & btb_251_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_251_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_251_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_251_bht_T_13 = _btb_0_bht_T_8 & _btb_251_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_251_bht_T_16 = _btb_0_bht_T_8 & _btb_251_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_251_bht_T_19 = _btb_0_bht_T_8 & _btb_251_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_251_bht_T_20 = _btb_251_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_21 = _btb_251_bht_T_16 ? 2'h0 : _btb_251_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_22 = _btb_251_bht_T_13 ? 2'h0 : _btb_251_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_23 = _btb_251_bht_T_10 ? 2'h0 : _btb_251_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_24 = _btb_251_bht_T_7 ? 2'h3 : _btb_251_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_25 = _btb_251_bht_T_5 ? 2'h3 : _btb_251_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_26 = _btb_251_bht_T_3 ? 2'h3 : _btb_251_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_251_bht_T_27 = _btb_251_bht_T_1 ? 2'h1 : _btb_251_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9710 = btb_251_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6907
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9712 = btb_251_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_251_bht_T_27 : _GEN_8443; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_252_bht_T = btb_252_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_252_bht_T_1 = io_i_branch_resolve_pack_taken & btb_252_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_252_bht_T_2 = btb_252_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_252_bht_T_3 = io_i_branch_resolve_pack_taken & btb_252_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_252_bht_T_4 = btb_252_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_252_bht_T_5 = io_i_branch_resolve_pack_taken & btb_252_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_252_bht_T_6 = btb_252_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_252_bht_T_7 = io_i_branch_resolve_pack_taken & btb_252_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_252_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_252_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_252_bht_T_13 = _btb_0_bht_T_8 & _btb_252_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_252_bht_T_16 = _btb_0_bht_T_8 & _btb_252_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_252_bht_T_19 = _btb_0_bht_T_8 & _btb_252_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_252_bht_T_20 = _btb_252_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_21 = _btb_252_bht_T_16 ? 2'h0 : _btb_252_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_22 = _btb_252_bht_T_13 ? 2'h0 : _btb_252_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_23 = _btb_252_bht_T_10 ? 2'h0 : _btb_252_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_24 = _btb_252_bht_T_7 ? 2'h3 : _btb_252_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_25 = _btb_252_bht_T_5 ? 2'h3 : _btb_252_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_26 = _btb_252_bht_T_3 ? 2'h3 : _btb_252_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_252_bht_T_27 = _btb_252_bht_T_1 ? 2'h1 : _btb_252_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9714 = btb_252_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6908
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9716 = btb_252_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_252_bht_T_27 : _GEN_8444; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_253_bht_T = btb_253_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_253_bht_T_1 = io_i_branch_resolve_pack_taken & btb_253_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_253_bht_T_2 = btb_253_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_253_bht_T_3 = io_i_branch_resolve_pack_taken & btb_253_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_253_bht_T_4 = btb_253_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_253_bht_T_5 = io_i_branch_resolve_pack_taken & btb_253_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_253_bht_T_6 = btb_253_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_253_bht_T_7 = io_i_branch_resolve_pack_taken & btb_253_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_253_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_253_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_253_bht_T_13 = _btb_0_bht_T_8 & _btb_253_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_253_bht_T_16 = _btb_0_bht_T_8 & _btb_253_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_253_bht_T_19 = _btb_0_bht_T_8 & _btb_253_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_253_bht_T_20 = _btb_253_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_21 = _btb_253_bht_T_16 ? 2'h0 : _btb_253_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_22 = _btb_253_bht_T_13 ? 2'h0 : _btb_253_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_23 = _btb_253_bht_T_10 ? 2'h0 : _btb_253_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_24 = _btb_253_bht_T_7 ? 2'h3 : _btb_253_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_25 = _btb_253_bht_T_5 ? 2'h3 : _btb_253_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_26 = _btb_253_bht_T_3 ? 2'h3 : _btb_253_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_253_bht_T_27 = _btb_253_bht_T_1 ? 2'h1 : _btb_253_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9718 = btb_253_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6909
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9720 = btb_253_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_253_bht_T_27 : _GEN_8445; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_254_bht_T = btb_254_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_254_bht_T_1 = io_i_branch_resolve_pack_taken & btb_254_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_254_bht_T_2 = btb_254_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_254_bht_T_3 = io_i_branch_resolve_pack_taken & btb_254_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_254_bht_T_4 = btb_254_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_254_bht_T_5 = io_i_branch_resolve_pack_taken & btb_254_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_254_bht_T_6 = btb_254_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_254_bht_T_7 = io_i_branch_resolve_pack_taken & btb_254_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_254_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_254_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_254_bht_T_13 = _btb_0_bht_T_8 & _btb_254_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_254_bht_T_16 = _btb_0_bht_T_8 & _btb_254_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_254_bht_T_19 = _btb_0_bht_T_8 & _btb_254_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_254_bht_T_20 = _btb_254_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_21 = _btb_254_bht_T_16 ? 2'h0 : _btb_254_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_22 = _btb_254_bht_T_13 ? 2'h0 : _btb_254_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_23 = _btb_254_bht_T_10 ? 2'h0 : _btb_254_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_24 = _btb_254_bht_T_7 ? 2'h3 : _btb_254_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_25 = _btb_254_bht_T_5 ? 2'h3 : _btb_254_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_26 = _btb_254_bht_T_3 ? 2'h3 : _btb_254_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_254_bht_T_27 = _btb_254_bht_T_1 ? 2'h1 : _btb_254_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9721 = btb_254_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_253_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_252_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_251_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_250_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_249_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_248_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_247_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_246_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_245_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_244_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_243_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_242_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_241_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_240_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9661)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9722 = btb_254_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6910
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9724 = btb_254_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_254_bht_T_27 : _GEN_8446; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_255_bht_T = btb_255_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_255_bht_T_1 = io_i_branch_resolve_pack_taken & btb_255_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_255_bht_T_2 = btb_255_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_255_bht_T_3 = io_i_branch_resolve_pack_taken & btb_255_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_255_bht_T_4 = btb_255_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_255_bht_T_5 = io_i_branch_resolve_pack_taken & btb_255_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_255_bht_T_6 = btb_255_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_255_bht_T_7 = io_i_branch_resolve_pack_taken & btb_255_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_255_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_255_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_255_bht_T_13 = _btb_0_bht_T_8 & _btb_255_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_255_bht_T_16 = _btb_0_bht_T_8 & _btb_255_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_255_bht_T_19 = _btb_0_bht_T_8 & _btb_255_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_255_bht_T_20 = _btb_255_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_21 = _btb_255_bht_T_16 ? 2'h0 : _btb_255_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_22 = _btb_255_bht_T_13 ? 2'h0 : _btb_255_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_23 = _btb_255_bht_T_10 ? 2'h0 : _btb_255_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_24 = _btb_255_bht_T_7 ? 2'h3 : _btb_255_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_25 = _btb_255_bht_T_5 ? 2'h3 : _btb_255_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_26 = _btb_255_bht_T_3 ? 2'h3 : _btb_255_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_255_bht_T_27 = _btb_255_bht_T_1 ? 2'h1 : _btb_255_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9726 = btb_255_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6911
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9728 = btb_255_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_255_bht_T_27 : _GEN_8447; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_256_bht_T = btb_256_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_256_bht_T_1 = io_i_branch_resolve_pack_taken & btb_256_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_256_bht_T_2 = btb_256_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_256_bht_T_3 = io_i_branch_resolve_pack_taken & btb_256_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_256_bht_T_4 = btb_256_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_256_bht_T_5 = io_i_branch_resolve_pack_taken & btb_256_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_256_bht_T_6 = btb_256_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_256_bht_T_7 = io_i_branch_resolve_pack_taken & btb_256_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_256_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_256_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_256_bht_T_13 = _btb_0_bht_T_8 & _btb_256_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_256_bht_T_16 = _btb_0_bht_T_8 & _btb_256_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_256_bht_T_19 = _btb_0_bht_T_8 & _btb_256_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_256_bht_T_20 = _btb_256_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_21 = _btb_256_bht_T_16 ? 2'h0 : _btb_256_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_22 = _btb_256_bht_T_13 ? 2'h0 : _btb_256_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_23 = _btb_256_bht_T_10 ? 2'h0 : _btb_256_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_24 = _btb_256_bht_T_7 ? 2'h3 : _btb_256_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_25 = _btb_256_bht_T_5 ? 2'h3 : _btb_256_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_26 = _btb_256_bht_T_3 ? 2'h3 : _btb_256_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_256_bht_T_27 = _btb_256_bht_T_1 ? 2'h1 : _btb_256_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9730 = btb_256_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6912
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9732 = btb_256_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_256_bht_T_27 : _GEN_8448; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_257_bht_T = btb_257_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_257_bht_T_1 = io_i_branch_resolve_pack_taken & btb_257_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_257_bht_T_2 = btb_257_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_257_bht_T_3 = io_i_branch_resolve_pack_taken & btb_257_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_257_bht_T_4 = btb_257_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_257_bht_T_5 = io_i_branch_resolve_pack_taken & btb_257_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_257_bht_T_6 = btb_257_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_257_bht_T_7 = io_i_branch_resolve_pack_taken & btb_257_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_257_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_257_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_257_bht_T_13 = _btb_0_bht_T_8 & _btb_257_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_257_bht_T_16 = _btb_0_bht_T_8 & _btb_257_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_257_bht_T_19 = _btb_0_bht_T_8 & _btb_257_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_257_bht_T_20 = _btb_257_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_21 = _btb_257_bht_T_16 ? 2'h0 : _btb_257_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_22 = _btb_257_bht_T_13 ? 2'h0 : _btb_257_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_23 = _btb_257_bht_T_10 ? 2'h0 : _btb_257_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_24 = _btb_257_bht_T_7 ? 2'h3 : _btb_257_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_25 = _btb_257_bht_T_5 ? 2'h3 : _btb_257_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_26 = _btb_257_bht_T_3 ? 2'h3 : _btb_257_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_257_bht_T_27 = _btb_257_bht_T_1 ? 2'h1 : _btb_257_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9734 = btb_257_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6913
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9736 = btb_257_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_257_bht_T_27 : _GEN_8449; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_258_bht_T = btb_258_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_258_bht_T_1 = io_i_branch_resolve_pack_taken & btb_258_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_258_bht_T_2 = btb_258_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_258_bht_T_3 = io_i_branch_resolve_pack_taken & btb_258_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_258_bht_T_4 = btb_258_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_258_bht_T_5 = io_i_branch_resolve_pack_taken & btb_258_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_258_bht_T_6 = btb_258_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_258_bht_T_7 = io_i_branch_resolve_pack_taken & btb_258_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_258_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_258_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_258_bht_T_13 = _btb_0_bht_T_8 & _btb_258_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_258_bht_T_16 = _btb_0_bht_T_8 & _btb_258_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_258_bht_T_19 = _btb_0_bht_T_8 & _btb_258_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_258_bht_T_20 = _btb_258_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_21 = _btb_258_bht_T_16 ? 2'h0 : _btb_258_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_22 = _btb_258_bht_T_13 ? 2'h0 : _btb_258_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_23 = _btb_258_bht_T_10 ? 2'h0 : _btb_258_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_24 = _btb_258_bht_T_7 ? 2'h3 : _btb_258_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_25 = _btb_258_bht_T_5 ? 2'h3 : _btb_258_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_26 = _btb_258_bht_T_3 ? 2'h3 : _btb_258_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_258_bht_T_27 = _btb_258_bht_T_1 ? 2'h1 : _btb_258_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9738 = btb_258_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6914
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9740 = btb_258_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_258_bht_T_27 : _GEN_8450; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_259_bht_T = btb_259_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_259_bht_T_1 = io_i_branch_resolve_pack_taken & btb_259_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_259_bht_T_2 = btb_259_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_259_bht_T_3 = io_i_branch_resolve_pack_taken & btb_259_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_259_bht_T_4 = btb_259_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_259_bht_T_5 = io_i_branch_resolve_pack_taken & btb_259_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_259_bht_T_6 = btb_259_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_259_bht_T_7 = io_i_branch_resolve_pack_taken & btb_259_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_259_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_259_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_259_bht_T_13 = _btb_0_bht_T_8 & _btb_259_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_259_bht_T_16 = _btb_0_bht_T_8 & _btb_259_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_259_bht_T_19 = _btb_0_bht_T_8 & _btb_259_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_259_bht_T_20 = _btb_259_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_21 = _btb_259_bht_T_16 ? 2'h0 : _btb_259_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_22 = _btb_259_bht_T_13 ? 2'h0 : _btb_259_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_23 = _btb_259_bht_T_10 ? 2'h0 : _btb_259_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_24 = _btb_259_bht_T_7 ? 2'h3 : _btb_259_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_25 = _btb_259_bht_T_5 ? 2'h3 : _btb_259_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_26 = _btb_259_bht_T_3 ? 2'h3 : _btb_259_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_259_bht_T_27 = _btb_259_bht_T_1 ? 2'h1 : _btb_259_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9742 = btb_259_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6915
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9744 = btb_259_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_259_bht_T_27 : _GEN_8451; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_260_bht_T = btb_260_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_260_bht_T_1 = io_i_branch_resolve_pack_taken & btb_260_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_260_bht_T_2 = btb_260_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_260_bht_T_3 = io_i_branch_resolve_pack_taken & btb_260_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_260_bht_T_4 = btb_260_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_260_bht_T_5 = io_i_branch_resolve_pack_taken & btb_260_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_260_bht_T_6 = btb_260_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_260_bht_T_7 = io_i_branch_resolve_pack_taken & btb_260_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_260_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_260_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_260_bht_T_13 = _btb_0_bht_T_8 & _btb_260_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_260_bht_T_16 = _btb_0_bht_T_8 & _btb_260_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_260_bht_T_19 = _btb_0_bht_T_8 & _btb_260_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_260_bht_T_20 = _btb_260_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_21 = _btb_260_bht_T_16 ? 2'h0 : _btb_260_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_22 = _btb_260_bht_T_13 ? 2'h0 : _btb_260_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_23 = _btb_260_bht_T_10 ? 2'h0 : _btb_260_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_24 = _btb_260_bht_T_7 ? 2'h3 : _btb_260_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_25 = _btb_260_bht_T_5 ? 2'h3 : _btb_260_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_26 = _btb_260_bht_T_3 ? 2'h3 : _btb_260_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_260_bht_T_27 = _btb_260_bht_T_1 ? 2'h1 : _btb_260_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9746 = btb_260_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6916
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9748 = btb_260_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_260_bht_T_27 : _GEN_8452; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_261_bht_T = btb_261_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_261_bht_T_1 = io_i_branch_resolve_pack_taken & btb_261_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_261_bht_T_2 = btb_261_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_261_bht_T_3 = io_i_branch_resolve_pack_taken & btb_261_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_261_bht_T_4 = btb_261_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_261_bht_T_5 = io_i_branch_resolve_pack_taken & btb_261_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_261_bht_T_6 = btb_261_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_261_bht_T_7 = io_i_branch_resolve_pack_taken & btb_261_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_261_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_261_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_261_bht_T_13 = _btb_0_bht_T_8 & _btb_261_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_261_bht_T_16 = _btb_0_bht_T_8 & _btb_261_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_261_bht_T_19 = _btb_0_bht_T_8 & _btb_261_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_261_bht_T_20 = _btb_261_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_21 = _btb_261_bht_T_16 ? 2'h0 : _btb_261_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_22 = _btb_261_bht_T_13 ? 2'h0 : _btb_261_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_23 = _btb_261_bht_T_10 ? 2'h0 : _btb_261_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_24 = _btb_261_bht_T_7 ? 2'h3 : _btb_261_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_25 = _btb_261_bht_T_5 ? 2'h3 : _btb_261_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_26 = _btb_261_bht_T_3 ? 2'h3 : _btb_261_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_261_bht_T_27 = _btb_261_bht_T_1 ? 2'h1 : _btb_261_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9750 = btb_261_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6917
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9752 = btb_261_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_261_bht_T_27 : _GEN_8453; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_262_bht_T = btb_262_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_262_bht_T_1 = io_i_branch_resolve_pack_taken & btb_262_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_262_bht_T_2 = btb_262_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_262_bht_T_3 = io_i_branch_resolve_pack_taken & btb_262_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_262_bht_T_4 = btb_262_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_262_bht_T_5 = io_i_branch_resolve_pack_taken & btb_262_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_262_bht_T_6 = btb_262_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_262_bht_T_7 = io_i_branch_resolve_pack_taken & btb_262_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_262_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_262_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_262_bht_T_13 = _btb_0_bht_T_8 & _btb_262_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_262_bht_T_16 = _btb_0_bht_T_8 & _btb_262_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_262_bht_T_19 = _btb_0_bht_T_8 & _btb_262_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_262_bht_T_20 = _btb_262_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_21 = _btb_262_bht_T_16 ? 2'h0 : _btb_262_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_22 = _btb_262_bht_T_13 ? 2'h0 : _btb_262_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_23 = _btb_262_bht_T_10 ? 2'h0 : _btb_262_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_24 = _btb_262_bht_T_7 ? 2'h3 : _btb_262_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_25 = _btb_262_bht_T_5 ? 2'h3 : _btb_262_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_26 = _btb_262_bht_T_3 ? 2'h3 : _btb_262_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_262_bht_T_27 = _btb_262_bht_T_1 ? 2'h1 : _btb_262_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9754 = btb_262_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6918
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9756 = btb_262_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_262_bht_T_27 : _GEN_8454; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_263_bht_T = btb_263_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_263_bht_T_1 = io_i_branch_resolve_pack_taken & btb_263_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_263_bht_T_2 = btb_263_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_263_bht_T_3 = io_i_branch_resolve_pack_taken & btb_263_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_263_bht_T_4 = btb_263_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_263_bht_T_5 = io_i_branch_resolve_pack_taken & btb_263_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_263_bht_T_6 = btb_263_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_263_bht_T_7 = io_i_branch_resolve_pack_taken & btb_263_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_263_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_263_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_263_bht_T_13 = _btb_0_bht_T_8 & _btb_263_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_263_bht_T_16 = _btb_0_bht_T_8 & _btb_263_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_263_bht_T_19 = _btb_0_bht_T_8 & _btb_263_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_263_bht_T_20 = _btb_263_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_21 = _btb_263_bht_T_16 ? 2'h0 : _btb_263_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_22 = _btb_263_bht_T_13 ? 2'h0 : _btb_263_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_23 = _btb_263_bht_T_10 ? 2'h0 : _btb_263_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_24 = _btb_263_bht_T_7 ? 2'h3 : _btb_263_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_25 = _btb_263_bht_T_5 ? 2'h3 : _btb_263_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_26 = _btb_263_bht_T_3 ? 2'h3 : _btb_263_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_263_bht_T_27 = _btb_263_bht_T_1 ? 2'h1 : _btb_263_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9758 = btb_263_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6919
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9760 = btb_263_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_263_bht_T_27 : _GEN_8455; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_264_bht_T = btb_264_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_264_bht_T_1 = io_i_branch_resolve_pack_taken & btb_264_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_264_bht_T_2 = btb_264_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_264_bht_T_3 = io_i_branch_resolve_pack_taken & btb_264_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_264_bht_T_4 = btb_264_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_264_bht_T_5 = io_i_branch_resolve_pack_taken & btb_264_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_264_bht_T_6 = btb_264_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_264_bht_T_7 = io_i_branch_resolve_pack_taken & btb_264_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_264_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_264_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_264_bht_T_13 = _btb_0_bht_T_8 & _btb_264_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_264_bht_T_16 = _btb_0_bht_T_8 & _btb_264_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_264_bht_T_19 = _btb_0_bht_T_8 & _btb_264_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_264_bht_T_20 = _btb_264_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_21 = _btb_264_bht_T_16 ? 2'h0 : _btb_264_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_22 = _btb_264_bht_T_13 ? 2'h0 : _btb_264_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_23 = _btb_264_bht_T_10 ? 2'h0 : _btb_264_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_24 = _btb_264_bht_T_7 ? 2'h3 : _btb_264_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_25 = _btb_264_bht_T_5 ? 2'h3 : _btb_264_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_26 = _btb_264_bht_T_3 ? 2'h3 : _btb_264_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_264_bht_T_27 = _btb_264_bht_T_1 ? 2'h1 : _btb_264_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9762 = btb_264_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6920
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9764 = btb_264_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_264_bht_T_27 : _GEN_8456; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_265_bht_T = btb_265_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_265_bht_T_1 = io_i_branch_resolve_pack_taken & btb_265_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_265_bht_T_2 = btb_265_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_265_bht_T_3 = io_i_branch_resolve_pack_taken & btb_265_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_265_bht_T_4 = btb_265_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_265_bht_T_5 = io_i_branch_resolve_pack_taken & btb_265_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_265_bht_T_6 = btb_265_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_265_bht_T_7 = io_i_branch_resolve_pack_taken & btb_265_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_265_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_265_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_265_bht_T_13 = _btb_0_bht_T_8 & _btb_265_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_265_bht_T_16 = _btb_0_bht_T_8 & _btb_265_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_265_bht_T_19 = _btb_0_bht_T_8 & _btb_265_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_265_bht_T_20 = _btb_265_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_21 = _btb_265_bht_T_16 ? 2'h0 : _btb_265_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_22 = _btb_265_bht_T_13 ? 2'h0 : _btb_265_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_23 = _btb_265_bht_T_10 ? 2'h0 : _btb_265_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_24 = _btb_265_bht_T_7 ? 2'h3 : _btb_265_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_25 = _btb_265_bht_T_5 ? 2'h3 : _btb_265_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_26 = _btb_265_bht_T_3 ? 2'h3 : _btb_265_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_265_bht_T_27 = _btb_265_bht_T_1 ? 2'h1 : _btb_265_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9766 = btb_265_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6921
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9768 = btb_265_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_265_bht_T_27 : _GEN_8457; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_266_bht_T = btb_266_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_266_bht_T_1 = io_i_branch_resolve_pack_taken & btb_266_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_266_bht_T_2 = btb_266_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_266_bht_T_3 = io_i_branch_resolve_pack_taken & btb_266_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_266_bht_T_4 = btb_266_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_266_bht_T_5 = io_i_branch_resolve_pack_taken & btb_266_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_266_bht_T_6 = btb_266_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_266_bht_T_7 = io_i_branch_resolve_pack_taken & btb_266_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_266_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_266_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_266_bht_T_13 = _btb_0_bht_T_8 & _btb_266_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_266_bht_T_16 = _btb_0_bht_T_8 & _btb_266_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_266_bht_T_19 = _btb_0_bht_T_8 & _btb_266_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_266_bht_T_20 = _btb_266_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_21 = _btb_266_bht_T_16 ? 2'h0 : _btb_266_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_22 = _btb_266_bht_T_13 ? 2'h0 : _btb_266_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_23 = _btb_266_bht_T_10 ? 2'h0 : _btb_266_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_24 = _btb_266_bht_T_7 ? 2'h3 : _btb_266_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_25 = _btb_266_bht_T_5 ? 2'h3 : _btb_266_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_26 = _btb_266_bht_T_3 ? 2'h3 : _btb_266_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_266_bht_T_27 = _btb_266_bht_T_1 ? 2'h1 : _btb_266_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9770 = btb_266_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6922
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9772 = btb_266_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_266_bht_T_27 : _GEN_8458; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_267_bht_T = btb_267_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_267_bht_T_1 = io_i_branch_resolve_pack_taken & btb_267_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_267_bht_T_2 = btb_267_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_267_bht_T_3 = io_i_branch_resolve_pack_taken & btb_267_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_267_bht_T_4 = btb_267_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_267_bht_T_5 = io_i_branch_resolve_pack_taken & btb_267_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_267_bht_T_6 = btb_267_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_267_bht_T_7 = io_i_branch_resolve_pack_taken & btb_267_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_267_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_267_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_267_bht_T_13 = _btb_0_bht_T_8 & _btb_267_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_267_bht_T_16 = _btb_0_bht_T_8 & _btb_267_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_267_bht_T_19 = _btb_0_bht_T_8 & _btb_267_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_267_bht_T_20 = _btb_267_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_21 = _btb_267_bht_T_16 ? 2'h0 : _btb_267_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_22 = _btb_267_bht_T_13 ? 2'h0 : _btb_267_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_23 = _btb_267_bht_T_10 ? 2'h0 : _btb_267_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_24 = _btb_267_bht_T_7 ? 2'h3 : _btb_267_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_25 = _btb_267_bht_T_5 ? 2'h3 : _btb_267_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_26 = _btb_267_bht_T_3 ? 2'h3 : _btb_267_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_267_bht_T_27 = _btb_267_bht_T_1 ? 2'h1 : _btb_267_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9774 = btb_267_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6923
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9776 = btb_267_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_267_bht_T_27 : _GEN_8459; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_268_bht_T = btb_268_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_268_bht_T_1 = io_i_branch_resolve_pack_taken & btb_268_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_268_bht_T_2 = btb_268_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_268_bht_T_3 = io_i_branch_resolve_pack_taken & btb_268_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_268_bht_T_4 = btb_268_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_268_bht_T_5 = io_i_branch_resolve_pack_taken & btb_268_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_268_bht_T_6 = btb_268_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_268_bht_T_7 = io_i_branch_resolve_pack_taken & btb_268_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_268_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_268_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_268_bht_T_13 = _btb_0_bht_T_8 & _btb_268_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_268_bht_T_16 = _btb_0_bht_T_8 & _btb_268_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_268_bht_T_19 = _btb_0_bht_T_8 & _btb_268_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_268_bht_T_20 = _btb_268_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_21 = _btb_268_bht_T_16 ? 2'h0 : _btb_268_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_22 = _btb_268_bht_T_13 ? 2'h0 : _btb_268_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_23 = _btb_268_bht_T_10 ? 2'h0 : _btb_268_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_24 = _btb_268_bht_T_7 ? 2'h3 : _btb_268_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_25 = _btb_268_bht_T_5 ? 2'h3 : _btb_268_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_26 = _btb_268_bht_T_3 ? 2'h3 : _btb_268_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_268_bht_T_27 = _btb_268_bht_T_1 ? 2'h1 : _btb_268_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9778 = btb_268_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6924
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9780 = btb_268_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_268_bht_T_27 : _GEN_8460; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_269_bht_T = btb_269_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_269_bht_T_1 = io_i_branch_resolve_pack_taken & btb_269_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_269_bht_T_2 = btb_269_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_269_bht_T_3 = io_i_branch_resolve_pack_taken & btb_269_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_269_bht_T_4 = btb_269_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_269_bht_T_5 = io_i_branch_resolve_pack_taken & btb_269_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_269_bht_T_6 = btb_269_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_269_bht_T_7 = io_i_branch_resolve_pack_taken & btb_269_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_269_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_269_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_269_bht_T_13 = _btb_0_bht_T_8 & _btb_269_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_269_bht_T_16 = _btb_0_bht_T_8 & _btb_269_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_269_bht_T_19 = _btb_0_bht_T_8 & _btb_269_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_269_bht_T_20 = _btb_269_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_21 = _btb_269_bht_T_16 ? 2'h0 : _btb_269_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_22 = _btb_269_bht_T_13 ? 2'h0 : _btb_269_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_23 = _btb_269_bht_T_10 ? 2'h0 : _btb_269_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_24 = _btb_269_bht_T_7 ? 2'h3 : _btb_269_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_25 = _btb_269_bht_T_5 ? 2'h3 : _btb_269_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_26 = _btb_269_bht_T_3 ? 2'h3 : _btb_269_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_269_bht_T_27 = _btb_269_bht_T_1 ? 2'h1 : _btb_269_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9781 = btb_269_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_268_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_267_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_266_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_265_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_264_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_263_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_262_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_261_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_260_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_259_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_258_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_257_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_256_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_255_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9721)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9782 = btb_269_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6925
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9784 = btb_269_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_269_bht_T_27 : _GEN_8461; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_270_bht_T = btb_270_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_270_bht_T_1 = io_i_branch_resolve_pack_taken & btb_270_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_270_bht_T_2 = btb_270_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_270_bht_T_3 = io_i_branch_resolve_pack_taken & btb_270_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_270_bht_T_4 = btb_270_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_270_bht_T_5 = io_i_branch_resolve_pack_taken & btb_270_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_270_bht_T_6 = btb_270_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_270_bht_T_7 = io_i_branch_resolve_pack_taken & btb_270_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_270_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_270_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_270_bht_T_13 = _btb_0_bht_T_8 & _btb_270_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_270_bht_T_16 = _btb_0_bht_T_8 & _btb_270_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_270_bht_T_19 = _btb_0_bht_T_8 & _btb_270_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_270_bht_T_20 = _btb_270_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_21 = _btb_270_bht_T_16 ? 2'h0 : _btb_270_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_22 = _btb_270_bht_T_13 ? 2'h0 : _btb_270_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_23 = _btb_270_bht_T_10 ? 2'h0 : _btb_270_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_24 = _btb_270_bht_T_7 ? 2'h3 : _btb_270_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_25 = _btb_270_bht_T_5 ? 2'h3 : _btb_270_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_26 = _btb_270_bht_T_3 ? 2'h3 : _btb_270_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_270_bht_T_27 = _btb_270_bht_T_1 ? 2'h1 : _btb_270_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9786 = btb_270_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6926
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9788 = btb_270_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_270_bht_T_27 : _GEN_8462; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_271_bht_T = btb_271_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_271_bht_T_1 = io_i_branch_resolve_pack_taken & btb_271_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_271_bht_T_2 = btb_271_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_271_bht_T_3 = io_i_branch_resolve_pack_taken & btb_271_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_271_bht_T_4 = btb_271_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_271_bht_T_5 = io_i_branch_resolve_pack_taken & btb_271_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_271_bht_T_6 = btb_271_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_271_bht_T_7 = io_i_branch_resolve_pack_taken & btb_271_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_271_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_271_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_271_bht_T_13 = _btb_0_bht_T_8 & _btb_271_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_271_bht_T_16 = _btb_0_bht_T_8 & _btb_271_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_271_bht_T_19 = _btb_0_bht_T_8 & _btb_271_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_271_bht_T_20 = _btb_271_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_21 = _btb_271_bht_T_16 ? 2'h0 : _btb_271_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_22 = _btb_271_bht_T_13 ? 2'h0 : _btb_271_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_23 = _btb_271_bht_T_10 ? 2'h0 : _btb_271_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_24 = _btb_271_bht_T_7 ? 2'h3 : _btb_271_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_25 = _btb_271_bht_T_5 ? 2'h3 : _btb_271_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_26 = _btb_271_bht_T_3 ? 2'h3 : _btb_271_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_271_bht_T_27 = _btb_271_bht_T_1 ? 2'h1 : _btb_271_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9790 = btb_271_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6927
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9792 = btb_271_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_271_bht_T_27 : _GEN_8463; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_272_bht_T = btb_272_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_272_bht_T_1 = io_i_branch_resolve_pack_taken & btb_272_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_272_bht_T_2 = btb_272_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_272_bht_T_3 = io_i_branch_resolve_pack_taken & btb_272_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_272_bht_T_4 = btb_272_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_272_bht_T_5 = io_i_branch_resolve_pack_taken & btb_272_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_272_bht_T_6 = btb_272_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_272_bht_T_7 = io_i_branch_resolve_pack_taken & btb_272_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_272_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_272_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_272_bht_T_13 = _btb_0_bht_T_8 & _btb_272_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_272_bht_T_16 = _btb_0_bht_T_8 & _btb_272_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_272_bht_T_19 = _btb_0_bht_T_8 & _btb_272_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_272_bht_T_20 = _btb_272_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_21 = _btb_272_bht_T_16 ? 2'h0 : _btb_272_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_22 = _btb_272_bht_T_13 ? 2'h0 : _btb_272_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_23 = _btb_272_bht_T_10 ? 2'h0 : _btb_272_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_24 = _btb_272_bht_T_7 ? 2'h3 : _btb_272_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_25 = _btb_272_bht_T_5 ? 2'h3 : _btb_272_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_26 = _btb_272_bht_T_3 ? 2'h3 : _btb_272_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_272_bht_T_27 = _btb_272_bht_T_1 ? 2'h1 : _btb_272_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9794 = btb_272_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6928
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9796 = btb_272_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_272_bht_T_27 : _GEN_8464; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_273_bht_T = btb_273_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_273_bht_T_1 = io_i_branch_resolve_pack_taken & btb_273_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_273_bht_T_2 = btb_273_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_273_bht_T_3 = io_i_branch_resolve_pack_taken & btb_273_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_273_bht_T_4 = btb_273_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_273_bht_T_5 = io_i_branch_resolve_pack_taken & btb_273_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_273_bht_T_6 = btb_273_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_273_bht_T_7 = io_i_branch_resolve_pack_taken & btb_273_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_273_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_273_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_273_bht_T_13 = _btb_0_bht_T_8 & _btb_273_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_273_bht_T_16 = _btb_0_bht_T_8 & _btb_273_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_273_bht_T_19 = _btb_0_bht_T_8 & _btb_273_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_273_bht_T_20 = _btb_273_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_21 = _btb_273_bht_T_16 ? 2'h0 : _btb_273_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_22 = _btb_273_bht_T_13 ? 2'h0 : _btb_273_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_23 = _btb_273_bht_T_10 ? 2'h0 : _btb_273_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_24 = _btb_273_bht_T_7 ? 2'h3 : _btb_273_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_25 = _btb_273_bht_T_5 ? 2'h3 : _btb_273_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_26 = _btb_273_bht_T_3 ? 2'h3 : _btb_273_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_273_bht_T_27 = _btb_273_bht_T_1 ? 2'h1 : _btb_273_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9798 = btb_273_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6929
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9800 = btb_273_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_273_bht_T_27 : _GEN_8465; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_274_bht_T = btb_274_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_274_bht_T_1 = io_i_branch_resolve_pack_taken & btb_274_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_274_bht_T_2 = btb_274_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_274_bht_T_3 = io_i_branch_resolve_pack_taken & btb_274_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_274_bht_T_4 = btb_274_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_274_bht_T_5 = io_i_branch_resolve_pack_taken & btb_274_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_274_bht_T_6 = btb_274_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_274_bht_T_7 = io_i_branch_resolve_pack_taken & btb_274_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_274_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_274_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_274_bht_T_13 = _btb_0_bht_T_8 & _btb_274_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_274_bht_T_16 = _btb_0_bht_T_8 & _btb_274_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_274_bht_T_19 = _btb_0_bht_T_8 & _btb_274_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_274_bht_T_20 = _btb_274_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_21 = _btb_274_bht_T_16 ? 2'h0 : _btb_274_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_22 = _btb_274_bht_T_13 ? 2'h0 : _btb_274_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_23 = _btb_274_bht_T_10 ? 2'h0 : _btb_274_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_24 = _btb_274_bht_T_7 ? 2'h3 : _btb_274_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_25 = _btb_274_bht_T_5 ? 2'h3 : _btb_274_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_26 = _btb_274_bht_T_3 ? 2'h3 : _btb_274_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_274_bht_T_27 = _btb_274_bht_T_1 ? 2'h1 : _btb_274_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9802 = btb_274_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6930
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9804 = btb_274_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_274_bht_T_27 : _GEN_8466; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_275_bht_T = btb_275_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_275_bht_T_1 = io_i_branch_resolve_pack_taken & btb_275_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_275_bht_T_2 = btb_275_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_275_bht_T_3 = io_i_branch_resolve_pack_taken & btb_275_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_275_bht_T_4 = btb_275_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_275_bht_T_5 = io_i_branch_resolve_pack_taken & btb_275_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_275_bht_T_6 = btb_275_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_275_bht_T_7 = io_i_branch_resolve_pack_taken & btb_275_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_275_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_275_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_275_bht_T_13 = _btb_0_bht_T_8 & _btb_275_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_275_bht_T_16 = _btb_0_bht_T_8 & _btb_275_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_275_bht_T_19 = _btb_0_bht_T_8 & _btb_275_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_275_bht_T_20 = _btb_275_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_21 = _btb_275_bht_T_16 ? 2'h0 : _btb_275_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_22 = _btb_275_bht_T_13 ? 2'h0 : _btb_275_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_23 = _btb_275_bht_T_10 ? 2'h0 : _btb_275_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_24 = _btb_275_bht_T_7 ? 2'h3 : _btb_275_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_25 = _btb_275_bht_T_5 ? 2'h3 : _btb_275_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_26 = _btb_275_bht_T_3 ? 2'h3 : _btb_275_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_275_bht_T_27 = _btb_275_bht_T_1 ? 2'h1 : _btb_275_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9806 = btb_275_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6931
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9808 = btb_275_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_275_bht_T_27 : _GEN_8467; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_276_bht_T = btb_276_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_276_bht_T_1 = io_i_branch_resolve_pack_taken & btb_276_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_276_bht_T_2 = btb_276_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_276_bht_T_3 = io_i_branch_resolve_pack_taken & btb_276_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_276_bht_T_4 = btb_276_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_276_bht_T_5 = io_i_branch_resolve_pack_taken & btb_276_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_276_bht_T_6 = btb_276_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_276_bht_T_7 = io_i_branch_resolve_pack_taken & btb_276_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_276_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_276_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_276_bht_T_13 = _btb_0_bht_T_8 & _btb_276_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_276_bht_T_16 = _btb_0_bht_T_8 & _btb_276_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_276_bht_T_19 = _btb_0_bht_T_8 & _btb_276_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_276_bht_T_20 = _btb_276_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_21 = _btb_276_bht_T_16 ? 2'h0 : _btb_276_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_22 = _btb_276_bht_T_13 ? 2'h0 : _btb_276_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_23 = _btb_276_bht_T_10 ? 2'h0 : _btb_276_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_24 = _btb_276_bht_T_7 ? 2'h3 : _btb_276_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_25 = _btb_276_bht_T_5 ? 2'h3 : _btb_276_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_26 = _btb_276_bht_T_3 ? 2'h3 : _btb_276_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_276_bht_T_27 = _btb_276_bht_T_1 ? 2'h1 : _btb_276_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9810 = btb_276_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6932
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9812 = btb_276_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_276_bht_T_27 : _GEN_8468; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_277_bht_T = btb_277_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_277_bht_T_1 = io_i_branch_resolve_pack_taken & btb_277_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_277_bht_T_2 = btb_277_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_277_bht_T_3 = io_i_branch_resolve_pack_taken & btb_277_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_277_bht_T_4 = btb_277_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_277_bht_T_5 = io_i_branch_resolve_pack_taken & btb_277_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_277_bht_T_6 = btb_277_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_277_bht_T_7 = io_i_branch_resolve_pack_taken & btb_277_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_277_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_277_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_277_bht_T_13 = _btb_0_bht_T_8 & _btb_277_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_277_bht_T_16 = _btb_0_bht_T_8 & _btb_277_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_277_bht_T_19 = _btb_0_bht_T_8 & _btb_277_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_277_bht_T_20 = _btb_277_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_21 = _btb_277_bht_T_16 ? 2'h0 : _btb_277_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_22 = _btb_277_bht_T_13 ? 2'h0 : _btb_277_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_23 = _btb_277_bht_T_10 ? 2'h0 : _btb_277_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_24 = _btb_277_bht_T_7 ? 2'h3 : _btb_277_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_25 = _btb_277_bht_T_5 ? 2'h3 : _btb_277_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_26 = _btb_277_bht_T_3 ? 2'h3 : _btb_277_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_277_bht_T_27 = _btb_277_bht_T_1 ? 2'h1 : _btb_277_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9814 = btb_277_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6933
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9816 = btb_277_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_277_bht_T_27 : _GEN_8469; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_278_bht_T = btb_278_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_278_bht_T_1 = io_i_branch_resolve_pack_taken & btb_278_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_278_bht_T_2 = btb_278_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_278_bht_T_3 = io_i_branch_resolve_pack_taken & btb_278_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_278_bht_T_4 = btb_278_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_278_bht_T_5 = io_i_branch_resolve_pack_taken & btb_278_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_278_bht_T_6 = btb_278_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_278_bht_T_7 = io_i_branch_resolve_pack_taken & btb_278_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_278_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_278_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_278_bht_T_13 = _btb_0_bht_T_8 & _btb_278_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_278_bht_T_16 = _btb_0_bht_T_8 & _btb_278_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_278_bht_T_19 = _btb_0_bht_T_8 & _btb_278_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_278_bht_T_20 = _btb_278_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_21 = _btb_278_bht_T_16 ? 2'h0 : _btb_278_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_22 = _btb_278_bht_T_13 ? 2'h0 : _btb_278_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_23 = _btb_278_bht_T_10 ? 2'h0 : _btb_278_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_24 = _btb_278_bht_T_7 ? 2'h3 : _btb_278_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_25 = _btb_278_bht_T_5 ? 2'h3 : _btb_278_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_26 = _btb_278_bht_T_3 ? 2'h3 : _btb_278_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_278_bht_T_27 = _btb_278_bht_T_1 ? 2'h1 : _btb_278_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9818 = btb_278_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6934
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9820 = btb_278_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_278_bht_T_27 : _GEN_8470; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_279_bht_T = btb_279_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_279_bht_T_1 = io_i_branch_resolve_pack_taken & btb_279_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_279_bht_T_2 = btb_279_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_279_bht_T_3 = io_i_branch_resolve_pack_taken & btb_279_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_279_bht_T_4 = btb_279_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_279_bht_T_5 = io_i_branch_resolve_pack_taken & btb_279_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_279_bht_T_6 = btb_279_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_279_bht_T_7 = io_i_branch_resolve_pack_taken & btb_279_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_279_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_279_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_279_bht_T_13 = _btb_0_bht_T_8 & _btb_279_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_279_bht_T_16 = _btb_0_bht_T_8 & _btb_279_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_279_bht_T_19 = _btb_0_bht_T_8 & _btb_279_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_279_bht_T_20 = _btb_279_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_21 = _btb_279_bht_T_16 ? 2'h0 : _btb_279_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_22 = _btb_279_bht_T_13 ? 2'h0 : _btb_279_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_23 = _btb_279_bht_T_10 ? 2'h0 : _btb_279_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_24 = _btb_279_bht_T_7 ? 2'h3 : _btb_279_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_25 = _btb_279_bht_T_5 ? 2'h3 : _btb_279_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_26 = _btb_279_bht_T_3 ? 2'h3 : _btb_279_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_279_bht_T_27 = _btb_279_bht_T_1 ? 2'h1 : _btb_279_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9822 = btb_279_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6935
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9824 = btb_279_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_279_bht_T_27 : _GEN_8471; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_280_bht_T = btb_280_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_280_bht_T_1 = io_i_branch_resolve_pack_taken & btb_280_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_280_bht_T_2 = btb_280_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_280_bht_T_3 = io_i_branch_resolve_pack_taken & btb_280_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_280_bht_T_4 = btb_280_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_280_bht_T_5 = io_i_branch_resolve_pack_taken & btb_280_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_280_bht_T_6 = btb_280_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_280_bht_T_7 = io_i_branch_resolve_pack_taken & btb_280_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_280_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_280_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_280_bht_T_13 = _btb_0_bht_T_8 & _btb_280_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_280_bht_T_16 = _btb_0_bht_T_8 & _btb_280_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_280_bht_T_19 = _btb_0_bht_T_8 & _btb_280_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_280_bht_T_20 = _btb_280_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_21 = _btb_280_bht_T_16 ? 2'h0 : _btb_280_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_22 = _btb_280_bht_T_13 ? 2'h0 : _btb_280_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_23 = _btb_280_bht_T_10 ? 2'h0 : _btb_280_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_24 = _btb_280_bht_T_7 ? 2'h3 : _btb_280_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_25 = _btb_280_bht_T_5 ? 2'h3 : _btb_280_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_26 = _btb_280_bht_T_3 ? 2'h3 : _btb_280_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_280_bht_T_27 = _btb_280_bht_T_1 ? 2'h1 : _btb_280_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9826 = btb_280_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6936
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9828 = btb_280_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_280_bht_T_27 : _GEN_8472; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_281_bht_T = btb_281_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_281_bht_T_1 = io_i_branch_resolve_pack_taken & btb_281_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_281_bht_T_2 = btb_281_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_281_bht_T_3 = io_i_branch_resolve_pack_taken & btb_281_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_281_bht_T_4 = btb_281_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_281_bht_T_5 = io_i_branch_resolve_pack_taken & btb_281_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_281_bht_T_6 = btb_281_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_281_bht_T_7 = io_i_branch_resolve_pack_taken & btb_281_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_281_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_281_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_281_bht_T_13 = _btb_0_bht_T_8 & _btb_281_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_281_bht_T_16 = _btb_0_bht_T_8 & _btb_281_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_281_bht_T_19 = _btb_0_bht_T_8 & _btb_281_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_281_bht_T_20 = _btb_281_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_21 = _btb_281_bht_T_16 ? 2'h0 : _btb_281_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_22 = _btb_281_bht_T_13 ? 2'h0 : _btb_281_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_23 = _btb_281_bht_T_10 ? 2'h0 : _btb_281_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_24 = _btb_281_bht_T_7 ? 2'h3 : _btb_281_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_25 = _btb_281_bht_T_5 ? 2'h3 : _btb_281_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_26 = _btb_281_bht_T_3 ? 2'h3 : _btb_281_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_281_bht_T_27 = _btb_281_bht_T_1 ? 2'h1 : _btb_281_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9830 = btb_281_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6937
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9832 = btb_281_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_281_bht_T_27 : _GEN_8473; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_282_bht_T = btb_282_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_282_bht_T_1 = io_i_branch_resolve_pack_taken & btb_282_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_282_bht_T_2 = btb_282_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_282_bht_T_3 = io_i_branch_resolve_pack_taken & btb_282_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_282_bht_T_4 = btb_282_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_282_bht_T_5 = io_i_branch_resolve_pack_taken & btb_282_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_282_bht_T_6 = btb_282_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_282_bht_T_7 = io_i_branch_resolve_pack_taken & btb_282_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_282_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_282_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_282_bht_T_13 = _btb_0_bht_T_8 & _btb_282_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_282_bht_T_16 = _btb_0_bht_T_8 & _btb_282_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_282_bht_T_19 = _btb_0_bht_T_8 & _btb_282_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_282_bht_T_20 = _btb_282_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_21 = _btb_282_bht_T_16 ? 2'h0 : _btb_282_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_22 = _btb_282_bht_T_13 ? 2'h0 : _btb_282_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_23 = _btb_282_bht_T_10 ? 2'h0 : _btb_282_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_24 = _btb_282_bht_T_7 ? 2'h3 : _btb_282_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_25 = _btb_282_bht_T_5 ? 2'h3 : _btb_282_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_26 = _btb_282_bht_T_3 ? 2'h3 : _btb_282_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_282_bht_T_27 = _btb_282_bht_T_1 ? 2'h1 : _btb_282_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9834 = btb_282_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6938
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9836 = btb_282_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_282_bht_T_27 : _GEN_8474; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_283_bht_T = btb_283_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_283_bht_T_1 = io_i_branch_resolve_pack_taken & btb_283_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_283_bht_T_2 = btb_283_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_283_bht_T_3 = io_i_branch_resolve_pack_taken & btb_283_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_283_bht_T_4 = btb_283_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_283_bht_T_5 = io_i_branch_resolve_pack_taken & btb_283_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_283_bht_T_6 = btb_283_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_283_bht_T_7 = io_i_branch_resolve_pack_taken & btb_283_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_283_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_283_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_283_bht_T_13 = _btb_0_bht_T_8 & _btb_283_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_283_bht_T_16 = _btb_0_bht_T_8 & _btb_283_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_283_bht_T_19 = _btb_0_bht_T_8 & _btb_283_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_283_bht_T_20 = _btb_283_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_21 = _btb_283_bht_T_16 ? 2'h0 : _btb_283_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_22 = _btb_283_bht_T_13 ? 2'h0 : _btb_283_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_23 = _btb_283_bht_T_10 ? 2'h0 : _btb_283_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_24 = _btb_283_bht_T_7 ? 2'h3 : _btb_283_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_25 = _btb_283_bht_T_5 ? 2'h3 : _btb_283_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_26 = _btb_283_bht_T_3 ? 2'h3 : _btb_283_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_283_bht_T_27 = _btb_283_bht_T_1 ? 2'h1 : _btb_283_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9838 = btb_283_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6939
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9840 = btb_283_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_283_bht_T_27 : _GEN_8475; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_284_bht_T = btb_284_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_284_bht_T_1 = io_i_branch_resolve_pack_taken & btb_284_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_284_bht_T_2 = btb_284_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_284_bht_T_3 = io_i_branch_resolve_pack_taken & btb_284_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_284_bht_T_4 = btb_284_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_284_bht_T_5 = io_i_branch_resolve_pack_taken & btb_284_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_284_bht_T_6 = btb_284_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_284_bht_T_7 = io_i_branch_resolve_pack_taken & btb_284_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_284_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_284_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_284_bht_T_13 = _btb_0_bht_T_8 & _btb_284_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_284_bht_T_16 = _btb_0_bht_T_8 & _btb_284_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_284_bht_T_19 = _btb_0_bht_T_8 & _btb_284_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_284_bht_T_20 = _btb_284_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_21 = _btb_284_bht_T_16 ? 2'h0 : _btb_284_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_22 = _btb_284_bht_T_13 ? 2'h0 : _btb_284_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_23 = _btb_284_bht_T_10 ? 2'h0 : _btb_284_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_24 = _btb_284_bht_T_7 ? 2'h3 : _btb_284_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_25 = _btb_284_bht_T_5 ? 2'h3 : _btb_284_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_26 = _btb_284_bht_T_3 ? 2'h3 : _btb_284_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_284_bht_T_27 = _btb_284_bht_T_1 ? 2'h1 : _btb_284_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9841 = btb_284_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_283_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_282_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_281_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_280_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_279_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_278_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_277_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_276_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_275_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_274_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_273_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_272_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_271_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_270_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9781)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9842 = btb_284_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6940
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9844 = btb_284_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_284_bht_T_27 : _GEN_8476; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_285_bht_T = btb_285_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_285_bht_T_1 = io_i_branch_resolve_pack_taken & btb_285_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_285_bht_T_2 = btb_285_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_285_bht_T_3 = io_i_branch_resolve_pack_taken & btb_285_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_285_bht_T_4 = btb_285_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_285_bht_T_5 = io_i_branch_resolve_pack_taken & btb_285_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_285_bht_T_6 = btb_285_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_285_bht_T_7 = io_i_branch_resolve_pack_taken & btb_285_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_285_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_285_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_285_bht_T_13 = _btb_0_bht_T_8 & _btb_285_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_285_bht_T_16 = _btb_0_bht_T_8 & _btb_285_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_285_bht_T_19 = _btb_0_bht_T_8 & _btb_285_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_285_bht_T_20 = _btb_285_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_21 = _btb_285_bht_T_16 ? 2'h0 : _btb_285_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_22 = _btb_285_bht_T_13 ? 2'h0 : _btb_285_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_23 = _btb_285_bht_T_10 ? 2'h0 : _btb_285_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_24 = _btb_285_bht_T_7 ? 2'h3 : _btb_285_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_25 = _btb_285_bht_T_5 ? 2'h3 : _btb_285_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_26 = _btb_285_bht_T_3 ? 2'h3 : _btb_285_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_285_bht_T_27 = _btb_285_bht_T_1 ? 2'h1 : _btb_285_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9846 = btb_285_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6941
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9848 = btb_285_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_285_bht_T_27 : _GEN_8477; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_286_bht_T = btb_286_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_286_bht_T_1 = io_i_branch_resolve_pack_taken & btb_286_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_286_bht_T_2 = btb_286_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_286_bht_T_3 = io_i_branch_resolve_pack_taken & btb_286_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_286_bht_T_4 = btb_286_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_286_bht_T_5 = io_i_branch_resolve_pack_taken & btb_286_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_286_bht_T_6 = btb_286_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_286_bht_T_7 = io_i_branch_resolve_pack_taken & btb_286_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_286_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_286_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_286_bht_T_13 = _btb_0_bht_T_8 & _btb_286_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_286_bht_T_16 = _btb_0_bht_T_8 & _btb_286_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_286_bht_T_19 = _btb_0_bht_T_8 & _btb_286_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_286_bht_T_20 = _btb_286_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_21 = _btb_286_bht_T_16 ? 2'h0 : _btb_286_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_22 = _btb_286_bht_T_13 ? 2'h0 : _btb_286_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_23 = _btb_286_bht_T_10 ? 2'h0 : _btb_286_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_24 = _btb_286_bht_T_7 ? 2'h3 : _btb_286_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_25 = _btb_286_bht_T_5 ? 2'h3 : _btb_286_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_26 = _btb_286_bht_T_3 ? 2'h3 : _btb_286_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_286_bht_T_27 = _btb_286_bht_T_1 ? 2'h1 : _btb_286_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9850 = btb_286_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6942
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9852 = btb_286_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_286_bht_T_27 : _GEN_8478; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_287_bht_T = btb_287_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_287_bht_T_1 = io_i_branch_resolve_pack_taken & btb_287_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_287_bht_T_2 = btb_287_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_287_bht_T_3 = io_i_branch_resolve_pack_taken & btb_287_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_287_bht_T_4 = btb_287_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_287_bht_T_5 = io_i_branch_resolve_pack_taken & btb_287_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_287_bht_T_6 = btb_287_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_287_bht_T_7 = io_i_branch_resolve_pack_taken & btb_287_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_287_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_287_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_287_bht_T_13 = _btb_0_bht_T_8 & _btb_287_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_287_bht_T_16 = _btb_0_bht_T_8 & _btb_287_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_287_bht_T_19 = _btb_0_bht_T_8 & _btb_287_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_287_bht_T_20 = _btb_287_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_21 = _btb_287_bht_T_16 ? 2'h0 : _btb_287_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_22 = _btb_287_bht_T_13 ? 2'h0 : _btb_287_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_23 = _btb_287_bht_T_10 ? 2'h0 : _btb_287_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_24 = _btb_287_bht_T_7 ? 2'h3 : _btb_287_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_25 = _btb_287_bht_T_5 ? 2'h3 : _btb_287_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_26 = _btb_287_bht_T_3 ? 2'h3 : _btb_287_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_287_bht_T_27 = _btb_287_bht_T_1 ? 2'h1 : _btb_287_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9854 = btb_287_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6943
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9856 = btb_287_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_287_bht_T_27 : _GEN_8479; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_288_bht_T = btb_288_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_288_bht_T_1 = io_i_branch_resolve_pack_taken & btb_288_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_288_bht_T_2 = btb_288_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_288_bht_T_3 = io_i_branch_resolve_pack_taken & btb_288_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_288_bht_T_4 = btb_288_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_288_bht_T_5 = io_i_branch_resolve_pack_taken & btb_288_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_288_bht_T_6 = btb_288_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_288_bht_T_7 = io_i_branch_resolve_pack_taken & btb_288_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_288_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_288_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_288_bht_T_13 = _btb_0_bht_T_8 & _btb_288_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_288_bht_T_16 = _btb_0_bht_T_8 & _btb_288_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_288_bht_T_19 = _btb_0_bht_T_8 & _btb_288_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_288_bht_T_20 = _btb_288_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_21 = _btb_288_bht_T_16 ? 2'h0 : _btb_288_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_22 = _btb_288_bht_T_13 ? 2'h0 : _btb_288_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_23 = _btb_288_bht_T_10 ? 2'h0 : _btb_288_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_24 = _btb_288_bht_T_7 ? 2'h3 : _btb_288_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_25 = _btb_288_bht_T_5 ? 2'h3 : _btb_288_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_26 = _btb_288_bht_T_3 ? 2'h3 : _btb_288_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_288_bht_T_27 = _btb_288_bht_T_1 ? 2'h1 : _btb_288_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9858 = btb_288_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6944
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9860 = btb_288_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_288_bht_T_27 : _GEN_8480; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_289_bht_T = btb_289_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_289_bht_T_1 = io_i_branch_resolve_pack_taken & btb_289_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_289_bht_T_2 = btb_289_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_289_bht_T_3 = io_i_branch_resolve_pack_taken & btb_289_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_289_bht_T_4 = btb_289_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_289_bht_T_5 = io_i_branch_resolve_pack_taken & btb_289_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_289_bht_T_6 = btb_289_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_289_bht_T_7 = io_i_branch_resolve_pack_taken & btb_289_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_289_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_289_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_289_bht_T_13 = _btb_0_bht_T_8 & _btb_289_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_289_bht_T_16 = _btb_0_bht_T_8 & _btb_289_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_289_bht_T_19 = _btb_0_bht_T_8 & _btb_289_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_289_bht_T_20 = _btb_289_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_21 = _btb_289_bht_T_16 ? 2'h0 : _btb_289_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_22 = _btb_289_bht_T_13 ? 2'h0 : _btb_289_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_23 = _btb_289_bht_T_10 ? 2'h0 : _btb_289_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_24 = _btb_289_bht_T_7 ? 2'h3 : _btb_289_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_25 = _btb_289_bht_T_5 ? 2'h3 : _btb_289_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_26 = _btb_289_bht_T_3 ? 2'h3 : _btb_289_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_289_bht_T_27 = _btb_289_bht_T_1 ? 2'h1 : _btb_289_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9862 = btb_289_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6945
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9864 = btb_289_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_289_bht_T_27 : _GEN_8481; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_290_bht_T = btb_290_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_290_bht_T_1 = io_i_branch_resolve_pack_taken & btb_290_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_290_bht_T_2 = btb_290_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_290_bht_T_3 = io_i_branch_resolve_pack_taken & btb_290_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_290_bht_T_4 = btb_290_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_290_bht_T_5 = io_i_branch_resolve_pack_taken & btb_290_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_290_bht_T_6 = btb_290_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_290_bht_T_7 = io_i_branch_resolve_pack_taken & btb_290_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_290_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_290_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_290_bht_T_13 = _btb_0_bht_T_8 & _btb_290_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_290_bht_T_16 = _btb_0_bht_T_8 & _btb_290_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_290_bht_T_19 = _btb_0_bht_T_8 & _btb_290_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_290_bht_T_20 = _btb_290_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_21 = _btb_290_bht_T_16 ? 2'h0 : _btb_290_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_22 = _btb_290_bht_T_13 ? 2'h0 : _btb_290_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_23 = _btb_290_bht_T_10 ? 2'h0 : _btb_290_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_24 = _btb_290_bht_T_7 ? 2'h3 : _btb_290_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_25 = _btb_290_bht_T_5 ? 2'h3 : _btb_290_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_26 = _btb_290_bht_T_3 ? 2'h3 : _btb_290_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_290_bht_T_27 = _btb_290_bht_T_1 ? 2'h1 : _btb_290_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9866 = btb_290_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6946
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9868 = btb_290_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_290_bht_T_27 : _GEN_8482; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_291_bht_T = btb_291_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_291_bht_T_1 = io_i_branch_resolve_pack_taken & btb_291_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_291_bht_T_2 = btb_291_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_291_bht_T_3 = io_i_branch_resolve_pack_taken & btb_291_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_291_bht_T_4 = btb_291_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_291_bht_T_5 = io_i_branch_resolve_pack_taken & btb_291_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_291_bht_T_6 = btb_291_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_291_bht_T_7 = io_i_branch_resolve_pack_taken & btb_291_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_291_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_291_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_291_bht_T_13 = _btb_0_bht_T_8 & _btb_291_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_291_bht_T_16 = _btb_0_bht_T_8 & _btb_291_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_291_bht_T_19 = _btb_0_bht_T_8 & _btb_291_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_291_bht_T_20 = _btb_291_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_21 = _btb_291_bht_T_16 ? 2'h0 : _btb_291_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_22 = _btb_291_bht_T_13 ? 2'h0 : _btb_291_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_23 = _btb_291_bht_T_10 ? 2'h0 : _btb_291_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_24 = _btb_291_bht_T_7 ? 2'h3 : _btb_291_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_25 = _btb_291_bht_T_5 ? 2'h3 : _btb_291_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_26 = _btb_291_bht_T_3 ? 2'h3 : _btb_291_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_291_bht_T_27 = _btb_291_bht_T_1 ? 2'h1 : _btb_291_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9870 = btb_291_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6947
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9872 = btb_291_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_291_bht_T_27 : _GEN_8483; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_292_bht_T = btb_292_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_292_bht_T_1 = io_i_branch_resolve_pack_taken & btb_292_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_292_bht_T_2 = btb_292_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_292_bht_T_3 = io_i_branch_resolve_pack_taken & btb_292_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_292_bht_T_4 = btb_292_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_292_bht_T_5 = io_i_branch_resolve_pack_taken & btb_292_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_292_bht_T_6 = btb_292_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_292_bht_T_7 = io_i_branch_resolve_pack_taken & btb_292_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_292_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_292_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_292_bht_T_13 = _btb_0_bht_T_8 & _btb_292_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_292_bht_T_16 = _btb_0_bht_T_8 & _btb_292_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_292_bht_T_19 = _btb_0_bht_T_8 & _btb_292_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_292_bht_T_20 = _btb_292_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_21 = _btb_292_bht_T_16 ? 2'h0 : _btb_292_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_22 = _btb_292_bht_T_13 ? 2'h0 : _btb_292_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_23 = _btb_292_bht_T_10 ? 2'h0 : _btb_292_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_24 = _btb_292_bht_T_7 ? 2'h3 : _btb_292_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_25 = _btb_292_bht_T_5 ? 2'h3 : _btb_292_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_26 = _btb_292_bht_T_3 ? 2'h3 : _btb_292_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_292_bht_T_27 = _btb_292_bht_T_1 ? 2'h1 : _btb_292_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9874 = btb_292_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6948
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9876 = btb_292_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_292_bht_T_27 : _GEN_8484; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_293_bht_T = btb_293_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_293_bht_T_1 = io_i_branch_resolve_pack_taken & btb_293_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_293_bht_T_2 = btb_293_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_293_bht_T_3 = io_i_branch_resolve_pack_taken & btb_293_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_293_bht_T_4 = btb_293_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_293_bht_T_5 = io_i_branch_resolve_pack_taken & btb_293_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_293_bht_T_6 = btb_293_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_293_bht_T_7 = io_i_branch_resolve_pack_taken & btb_293_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_293_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_293_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_293_bht_T_13 = _btb_0_bht_T_8 & _btb_293_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_293_bht_T_16 = _btb_0_bht_T_8 & _btb_293_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_293_bht_T_19 = _btb_0_bht_T_8 & _btb_293_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_293_bht_T_20 = _btb_293_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_21 = _btb_293_bht_T_16 ? 2'h0 : _btb_293_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_22 = _btb_293_bht_T_13 ? 2'h0 : _btb_293_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_23 = _btb_293_bht_T_10 ? 2'h0 : _btb_293_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_24 = _btb_293_bht_T_7 ? 2'h3 : _btb_293_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_25 = _btb_293_bht_T_5 ? 2'h3 : _btb_293_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_26 = _btb_293_bht_T_3 ? 2'h3 : _btb_293_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_293_bht_T_27 = _btb_293_bht_T_1 ? 2'h1 : _btb_293_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9878 = btb_293_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6949
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9880 = btb_293_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_293_bht_T_27 : _GEN_8485; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_294_bht_T = btb_294_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_294_bht_T_1 = io_i_branch_resolve_pack_taken & btb_294_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_294_bht_T_2 = btb_294_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_294_bht_T_3 = io_i_branch_resolve_pack_taken & btb_294_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_294_bht_T_4 = btb_294_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_294_bht_T_5 = io_i_branch_resolve_pack_taken & btb_294_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_294_bht_T_6 = btb_294_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_294_bht_T_7 = io_i_branch_resolve_pack_taken & btb_294_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_294_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_294_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_294_bht_T_13 = _btb_0_bht_T_8 & _btb_294_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_294_bht_T_16 = _btb_0_bht_T_8 & _btb_294_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_294_bht_T_19 = _btb_0_bht_T_8 & _btb_294_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_294_bht_T_20 = _btb_294_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_21 = _btb_294_bht_T_16 ? 2'h0 : _btb_294_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_22 = _btb_294_bht_T_13 ? 2'h0 : _btb_294_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_23 = _btb_294_bht_T_10 ? 2'h0 : _btb_294_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_24 = _btb_294_bht_T_7 ? 2'h3 : _btb_294_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_25 = _btb_294_bht_T_5 ? 2'h3 : _btb_294_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_26 = _btb_294_bht_T_3 ? 2'h3 : _btb_294_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_294_bht_T_27 = _btb_294_bht_T_1 ? 2'h1 : _btb_294_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9882 = btb_294_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6950
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9884 = btb_294_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_294_bht_T_27 : _GEN_8486; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_295_bht_T = btb_295_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_295_bht_T_1 = io_i_branch_resolve_pack_taken & btb_295_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_295_bht_T_2 = btb_295_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_295_bht_T_3 = io_i_branch_resolve_pack_taken & btb_295_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_295_bht_T_4 = btb_295_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_295_bht_T_5 = io_i_branch_resolve_pack_taken & btb_295_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_295_bht_T_6 = btb_295_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_295_bht_T_7 = io_i_branch_resolve_pack_taken & btb_295_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_295_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_295_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_295_bht_T_13 = _btb_0_bht_T_8 & _btb_295_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_295_bht_T_16 = _btb_0_bht_T_8 & _btb_295_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_295_bht_T_19 = _btb_0_bht_T_8 & _btb_295_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_295_bht_T_20 = _btb_295_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_21 = _btb_295_bht_T_16 ? 2'h0 : _btb_295_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_22 = _btb_295_bht_T_13 ? 2'h0 : _btb_295_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_23 = _btb_295_bht_T_10 ? 2'h0 : _btb_295_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_24 = _btb_295_bht_T_7 ? 2'h3 : _btb_295_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_25 = _btb_295_bht_T_5 ? 2'h3 : _btb_295_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_26 = _btb_295_bht_T_3 ? 2'h3 : _btb_295_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_295_bht_T_27 = _btb_295_bht_T_1 ? 2'h1 : _btb_295_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9886 = btb_295_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6951
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9888 = btb_295_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_295_bht_T_27 : _GEN_8487; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_296_bht_T = btb_296_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_296_bht_T_1 = io_i_branch_resolve_pack_taken & btb_296_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_296_bht_T_2 = btb_296_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_296_bht_T_3 = io_i_branch_resolve_pack_taken & btb_296_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_296_bht_T_4 = btb_296_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_296_bht_T_5 = io_i_branch_resolve_pack_taken & btb_296_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_296_bht_T_6 = btb_296_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_296_bht_T_7 = io_i_branch_resolve_pack_taken & btb_296_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_296_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_296_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_296_bht_T_13 = _btb_0_bht_T_8 & _btb_296_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_296_bht_T_16 = _btb_0_bht_T_8 & _btb_296_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_296_bht_T_19 = _btb_0_bht_T_8 & _btb_296_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_296_bht_T_20 = _btb_296_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_21 = _btb_296_bht_T_16 ? 2'h0 : _btb_296_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_22 = _btb_296_bht_T_13 ? 2'h0 : _btb_296_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_23 = _btb_296_bht_T_10 ? 2'h0 : _btb_296_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_24 = _btb_296_bht_T_7 ? 2'h3 : _btb_296_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_25 = _btb_296_bht_T_5 ? 2'h3 : _btb_296_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_26 = _btb_296_bht_T_3 ? 2'h3 : _btb_296_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_296_bht_T_27 = _btb_296_bht_T_1 ? 2'h1 : _btb_296_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9890 = btb_296_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6952
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9892 = btb_296_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_296_bht_T_27 : _GEN_8488; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_297_bht_T = btb_297_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_297_bht_T_1 = io_i_branch_resolve_pack_taken & btb_297_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_297_bht_T_2 = btb_297_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_297_bht_T_3 = io_i_branch_resolve_pack_taken & btb_297_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_297_bht_T_4 = btb_297_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_297_bht_T_5 = io_i_branch_resolve_pack_taken & btb_297_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_297_bht_T_6 = btb_297_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_297_bht_T_7 = io_i_branch_resolve_pack_taken & btb_297_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_297_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_297_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_297_bht_T_13 = _btb_0_bht_T_8 & _btb_297_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_297_bht_T_16 = _btb_0_bht_T_8 & _btb_297_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_297_bht_T_19 = _btb_0_bht_T_8 & _btb_297_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_297_bht_T_20 = _btb_297_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_21 = _btb_297_bht_T_16 ? 2'h0 : _btb_297_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_22 = _btb_297_bht_T_13 ? 2'h0 : _btb_297_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_23 = _btb_297_bht_T_10 ? 2'h0 : _btb_297_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_24 = _btb_297_bht_T_7 ? 2'h3 : _btb_297_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_25 = _btb_297_bht_T_5 ? 2'h3 : _btb_297_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_26 = _btb_297_bht_T_3 ? 2'h3 : _btb_297_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_297_bht_T_27 = _btb_297_bht_T_1 ? 2'h1 : _btb_297_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9894 = btb_297_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6953
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9896 = btb_297_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_297_bht_T_27 : _GEN_8489; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_298_bht_T = btb_298_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_298_bht_T_1 = io_i_branch_resolve_pack_taken & btb_298_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_298_bht_T_2 = btb_298_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_298_bht_T_3 = io_i_branch_resolve_pack_taken & btb_298_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_298_bht_T_4 = btb_298_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_298_bht_T_5 = io_i_branch_resolve_pack_taken & btb_298_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_298_bht_T_6 = btb_298_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_298_bht_T_7 = io_i_branch_resolve_pack_taken & btb_298_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_298_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_298_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_298_bht_T_13 = _btb_0_bht_T_8 & _btb_298_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_298_bht_T_16 = _btb_0_bht_T_8 & _btb_298_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_298_bht_T_19 = _btb_0_bht_T_8 & _btb_298_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_298_bht_T_20 = _btb_298_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_21 = _btb_298_bht_T_16 ? 2'h0 : _btb_298_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_22 = _btb_298_bht_T_13 ? 2'h0 : _btb_298_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_23 = _btb_298_bht_T_10 ? 2'h0 : _btb_298_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_24 = _btb_298_bht_T_7 ? 2'h3 : _btb_298_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_25 = _btb_298_bht_T_5 ? 2'h3 : _btb_298_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_26 = _btb_298_bht_T_3 ? 2'h3 : _btb_298_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_298_bht_T_27 = _btb_298_bht_T_1 ? 2'h1 : _btb_298_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9898 = btb_298_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6954
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9900 = btb_298_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_298_bht_T_27 : _GEN_8490; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_299_bht_T = btb_299_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_299_bht_T_1 = io_i_branch_resolve_pack_taken & btb_299_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_299_bht_T_2 = btb_299_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_299_bht_T_3 = io_i_branch_resolve_pack_taken & btb_299_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_299_bht_T_4 = btb_299_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_299_bht_T_5 = io_i_branch_resolve_pack_taken & btb_299_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_299_bht_T_6 = btb_299_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_299_bht_T_7 = io_i_branch_resolve_pack_taken & btb_299_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_299_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_299_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_299_bht_T_13 = _btb_0_bht_T_8 & _btb_299_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_299_bht_T_16 = _btb_0_bht_T_8 & _btb_299_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_299_bht_T_19 = _btb_0_bht_T_8 & _btb_299_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_299_bht_T_20 = _btb_299_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_21 = _btb_299_bht_T_16 ? 2'h0 : _btb_299_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_22 = _btb_299_bht_T_13 ? 2'h0 : _btb_299_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_23 = _btb_299_bht_T_10 ? 2'h0 : _btb_299_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_24 = _btb_299_bht_T_7 ? 2'h3 : _btb_299_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_25 = _btb_299_bht_T_5 ? 2'h3 : _btb_299_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_26 = _btb_299_bht_T_3 ? 2'h3 : _btb_299_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_299_bht_T_27 = _btb_299_bht_T_1 ? 2'h1 : _btb_299_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9901 = btb_299_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_298_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_297_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_296_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_295_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_294_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_293_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_292_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_291_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_290_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_289_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_288_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_287_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_286_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_285_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9841)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9902 = btb_299_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6955
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9904 = btb_299_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_299_bht_T_27 : _GEN_8491; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_300_bht_T = btb_300_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_300_bht_T_1 = io_i_branch_resolve_pack_taken & btb_300_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_300_bht_T_2 = btb_300_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_300_bht_T_3 = io_i_branch_resolve_pack_taken & btb_300_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_300_bht_T_4 = btb_300_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_300_bht_T_5 = io_i_branch_resolve_pack_taken & btb_300_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_300_bht_T_6 = btb_300_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_300_bht_T_7 = io_i_branch_resolve_pack_taken & btb_300_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_300_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_300_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_300_bht_T_13 = _btb_0_bht_T_8 & _btb_300_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_300_bht_T_16 = _btb_0_bht_T_8 & _btb_300_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_300_bht_T_19 = _btb_0_bht_T_8 & _btb_300_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_300_bht_T_20 = _btb_300_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_21 = _btb_300_bht_T_16 ? 2'h0 : _btb_300_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_22 = _btb_300_bht_T_13 ? 2'h0 : _btb_300_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_23 = _btb_300_bht_T_10 ? 2'h0 : _btb_300_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_24 = _btb_300_bht_T_7 ? 2'h3 : _btb_300_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_25 = _btb_300_bht_T_5 ? 2'h3 : _btb_300_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_26 = _btb_300_bht_T_3 ? 2'h3 : _btb_300_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_300_bht_T_27 = _btb_300_bht_T_1 ? 2'h1 : _btb_300_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9906 = btb_300_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6956
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9908 = btb_300_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_300_bht_T_27 : _GEN_8492; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_301_bht_T = btb_301_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_301_bht_T_1 = io_i_branch_resolve_pack_taken & btb_301_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_301_bht_T_2 = btb_301_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_301_bht_T_3 = io_i_branch_resolve_pack_taken & btb_301_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_301_bht_T_4 = btb_301_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_301_bht_T_5 = io_i_branch_resolve_pack_taken & btb_301_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_301_bht_T_6 = btb_301_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_301_bht_T_7 = io_i_branch_resolve_pack_taken & btb_301_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_301_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_301_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_301_bht_T_13 = _btb_0_bht_T_8 & _btb_301_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_301_bht_T_16 = _btb_0_bht_T_8 & _btb_301_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_301_bht_T_19 = _btb_0_bht_T_8 & _btb_301_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_301_bht_T_20 = _btb_301_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_21 = _btb_301_bht_T_16 ? 2'h0 : _btb_301_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_22 = _btb_301_bht_T_13 ? 2'h0 : _btb_301_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_23 = _btb_301_bht_T_10 ? 2'h0 : _btb_301_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_24 = _btb_301_bht_T_7 ? 2'h3 : _btb_301_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_25 = _btb_301_bht_T_5 ? 2'h3 : _btb_301_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_26 = _btb_301_bht_T_3 ? 2'h3 : _btb_301_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_301_bht_T_27 = _btb_301_bht_T_1 ? 2'h1 : _btb_301_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9910 = btb_301_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6957
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9912 = btb_301_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_301_bht_T_27 : _GEN_8493; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_302_bht_T = btb_302_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_302_bht_T_1 = io_i_branch_resolve_pack_taken & btb_302_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_302_bht_T_2 = btb_302_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_302_bht_T_3 = io_i_branch_resolve_pack_taken & btb_302_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_302_bht_T_4 = btb_302_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_302_bht_T_5 = io_i_branch_resolve_pack_taken & btb_302_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_302_bht_T_6 = btb_302_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_302_bht_T_7 = io_i_branch_resolve_pack_taken & btb_302_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_302_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_302_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_302_bht_T_13 = _btb_0_bht_T_8 & _btb_302_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_302_bht_T_16 = _btb_0_bht_T_8 & _btb_302_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_302_bht_T_19 = _btb_0_bht_T_8 & _btb_302_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_302_bht_T_20 = _btb_302_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_21 = _btb_302_bht_T_16 ? 2'h0 : _btb_302_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_22 = _btb_302_bht_T_13 ? 2'h0 : _btb_302_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_23 = _btb_302_bht_T_10 ? 2'h0 : _btb_302_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_24 = _btb_302_bht_T_7 ? 2'h3 : _btb_302_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_25 = _btb_302_bht_T_5 ? 2'h3 : _btb_302_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_26 = _btb_302_bht_T_3 ? 2'h3 : _btb_302_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_302_bht_T_27 = _btb_302_bht_T_1 ? 2'h1 : _btb_302_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9914 = btb_302_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6958
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9916 = btb_302_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_302_bht_T_27 : _GEN_8494; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_303_bht_T = btb_303_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_303_bht_T_1 = io_i_branch_resolve_pack_taken & btb_303_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_303_bht_T_2 = btb_303_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_303_bht_T_3 = io_i_branch_resolve_pack_taken & btb_303_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_303_bht_T_4 = btb_303_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_303_bht_T_5 = io_i_branch_resolve_pack_taken & btb_303_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_303_bht_T_6 = btb_303_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_303_bht_T_7 = io_i_branch_resolve_pack_taken & btb_303_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_303_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_303_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_303_bht_T_13 = _btb_0_bht_T_8 & _btb_303_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_303_bht_T_16 = _btb_0_bht_T_8 & _btb_303_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_303_bht_T_19 = _btb_0_bht_T_8 & _btb_303_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_303_bht_T_20 = _btb_303_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_21 = _btb_303_bht_T_16 ? 2'h0 : _btb_303_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_22 = _btb_303_bht_T_13 ? 2'h0 : _btb_303_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_23 = _btb_303_bht_T_10 ? 2'h0 : _btb_303_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_24 = _btb_303_bht_T_7 ? 2'h3 : _btb_303_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_25 = _btb_303_bht_T_5 ? 2'h3 : _btb_303_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_26 = _btb_303_bht_T_3 ? 2'h3 : _btb_303_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_303_bht_T_27 = _btb_303_bht_T_1 ? 2'h1 : _btb_303_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9918 = btb_303_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6959
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9920 = btb_303_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_303_bht_T_27 : _GEN_8495; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_304_bht_T = btb_304_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_304_bht_T_1 = io_i_branch_resolve_pack_taken & btb_304_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_304_bht_T_2 = btb_304_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_304_bht_T_3 = io_i_branch_resolve_pack_taken & btb_304_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_304_bht_T_4 = btb_304_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_304_bht_T_5 = io_i_branch_resolve_pack_taken & btb_304_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_304_bht_T_6 = btb_304_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_304_bht_T_7 = io_i_branch_resolve_pack_taken & btb_304_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_304_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_304_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_304_bht_T_13 = _btb_0_bht_T_8 & _btb_304_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_304_bht_T_16 = _btb_0_bht_T_8 & _btb_304_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_304_bht_T_19 = _btb_0_bht_T_8 & _btb_304_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_304_bht_T_20 = _btb_304_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_21 = _btb_304_bht_T_16 ? 2'h0 : _btb_304_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_22 = _btb_304_bht_T_13 ? 2'h0 : _btb_304_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_23 = _btb_304_bht_T_10 ? 2'h0 : _btb_304_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_24 = _btb_304_bht_T_7 ? 2'h3 : _btb_304_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_25 = _btb_304_bht_T_5 ? 2'h3 : _btb_304_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_26 = _btb_304_bht_T_3 ? 2'h3 : _btb_304_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_304_bht_T_27 = _btb_304_bht_T_1 ? 2'h1 : _btb_304_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9922 = btb_304_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6960
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9924 = btb_304_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_304_bht_T_27 : _GEN_8496; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_305_bht_T = btb_305_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_305_bht_T_1 = io_i_branch_resolve_pack_taken & btb_305_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_305_bht_T_2 = btb_305_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_305_bht_T_3 = io_i_branch_resolve_pack_taken & btb_305_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_305_bht_T_4 = btb_305_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_305_bht_T_5 = io_i_branch_resolve_pack_taken & btb_305_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_305_bht_T_6 = btb_305_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_305_bht_T_7 = io_i_branch_resolve_pack_taken & btb_305_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_305_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_305_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_305_bht_T_13 = _btb_0_bht_T_8 & _btb_305_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_305_bht_T_16 = _btb_0_bht_T_8 & _btb_305_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_305_bht_T_19 = _btb_0_bht_T_8 & _btb_305_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_305_bht_T_20 = _btb_305_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_21 = _btb_305_bht_T_16 ? 2'h0 : _btb_305_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_22 = _btb_305_bht_T_13 ? 2'h0 : _btb_305_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_23 = _btb_305_bht_T_10 ? 2'h0 : _btb_305_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_24 = _btb_305_bht_T_7 ? 2'h3 : _btb_305_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_25 = _btb_305_bht_T_5 ? 2'h3 : _btb_305_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_26 = _btb_305_bht_T_3 ? 2'h3 : _btb_305_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_305_bht_T_27 = _btb_305_bht_T_1 ? 2'h1 : _btb_305_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9926 = btb_305_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6961
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9928 = btb_305_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_305_bht_T_27 : _GEN_8497; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_306_bht_T = btb_306_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_306_bht_T_1 = io_i_branch_resolve_pack_taken & btb_306_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_306_bht_T_2 = btb_306_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_306_bht_T_3 = io_i_branch_resolve_pack_taken & btb_306_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_306_bht_T_4 = btb_306_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_306_bht_T_5 = io_i_branch_resolve_pack_taken & btb_306_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_306_bht_T_6 = btb_306_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_306_bht_T_7 = io_i_branch_resolve_pack_taken & btb_306_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_306_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_306_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_306_bht_T_13 = _btb_0_bht_T_8 & _btb_306_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_306_bht_T_16 = _btb_0_bht_T_8 & _btb_306_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_306_bht_T_19 = _btb_0_bht_T_8 & _btb_306_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_306_bht_T_20 = _btb_306_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_21 = _btb_306_bht_T_16 ? 2'h0 : _btb_306_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_22 = _btb_306_bht_T_13 ? 2'h0 : _btb_306_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_23 = _btb_306_bht_T_10 ? 2'h0 : _btb_306_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_24 = _btb_306_bht_T_7 ? 2'h3 : _btb_306_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_25 = _btb_306_bht_T_5 ? 2'h3 : _btb_306_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_26 = _btb_306_bht_T_3 ? 2'h3 : _btb_306_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_306_bht_T_27 = _btb_306_bht_T_1 ? 2'h1 : _btb_306_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9930 = btb_306_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6962
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9932 = btb_306_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_306_bht_T_27 : _GEN_8498; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_307_bht_T = btb_307_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_307_bht_T_1 = io_i_branch_resolve_pack_taken & btb_307_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_307_bht_T_2 = btb_307_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_307_bht_T_3 = io_i_branch_resolve_pack_taken & btb_307_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_307_bht_T_4 = btb_307_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_307_bht_T_5 = io_i_branch_resolve_pack_taken & btb_307_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_307_bht_T_6 = btb_307_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_307_bht_T_7 = io_i_branch_resolve_pack_taken & btb_307_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_307_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_307_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_307_bht_T_13 = _btb_0_bht_T_8 & _btb_307_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_307_bht_T_16 = _btb_0_bht_T_8 & _btb_307_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_307_bht_T_19 = _btb_0_bht_T_8 & _btb_307_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_307_bht_T_20 = _btb_307_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_21 = _btb_307_bht_T_16 ? 2'h0 : _btb_307_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_22 = _btb_307_bht_T_13 ? 2'h0 : _btb_307_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_23 = _btb_307_bht_T_10 ? 2'h0 : _btb_307_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_24 = _btb_307_bht_T_7 ? 2'h3 : _btb_307_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_25 = _btb_307_bht_T_5 ? 2'h3 : _btb_307_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_26 = _btb_307_bht_T_3 ? 2'h3 : _btb_307_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_307_bht_T_27 = _btb_307_bht_T_1 ? 2'h1 : _btb_307_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9934 = btb_307_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6963
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9936 = btb_307_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_307_bht_T_27 : _GEN_8499; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_308_bht_T = btb_308_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_308_bht_T_1 = io_i_branch_resolve_pack_taken & btb_308_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_308_bht_T_2 = btb_308_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_308_bht_T_3 = io_i_branch_resolve_pack_taken & btb_308_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_308_bht_T_4 = btb_308_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_308_bht_T_5 = io_i_branch_resolve_pack_taken & btb_308_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_308_bht_T_6 = btb_308_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_308_bht_T_7 = io_i_branch_resolve_pack_taken & btb_308_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_308_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_308_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_308_bht_T_13 = _btb_0_bht_T_8 & _btb_308_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_308_bht_T_16 = _btb_0_bht_T_8 & _btb_308_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_308_bht_T_19 = _btb_0_bht_T_8 & _btb_308_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_308_bht_T_20 = _btb_308_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_21 = _btb_308_bht_T_16 ? 2'h0 : _btb_308_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_22 = _btb_308_bht_T_13 ? 2'h0 : _btb_308_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_23 = _btb_308_bht_T_10 ? 2'h0 : _btb_308_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_24 = _btb_308_bht_T_7 ? 2'h3 : _btb_308_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_25 = _btb_308_bht_T_5 ? 2'h3 : _btb_308_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_26 = _btb_308_bht_T_3 ? 2'h3 : _btb_308_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_308_bht_T_27 = _btb_308_bht_T_1 ? 2'h1 : _btb_308_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9938 = btb_308_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6964
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9940 = btb_308_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_308_bht_T_27 : _GEN_8500; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_309_bht_T = btb_309_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_309_bht_T_1 = io_i_branch_resolve_pack_taken & btb_309_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_309_bht_T_2 = btb_309_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_309_bht_T_3 = io_i_branch_resolve_pack_taken & btb_309_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_309_bht_T_4 = btb_309_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_309_bht_T_5 = io_i_branch_resolve_pack_taken & btb_309_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_309_bht_T_6 = btb_309_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_309_bht_T_7 = io_i_branch_resolve_pack_taken & btb_309_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_309_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_309_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_309_bht_T_13 = _btb_0_bht_T_8 & _btb_309_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_309_bht_T_16 = _btb_0_bht_T_8 & _btb_309_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_309_bht_T_19 = _btb_0_bht_T_8 & _btb_309_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_309_bht_T_20 = _btb_309_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_21 = _btb_309_bht_T_16 ? 2'h0 : _btb_309_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_22 = _btb_309_bht_T_13 ? 2'h0 : _btb_309_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_23 = _btb_309_bht_T_10 ? 2'h0 : _btb_309_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_24 = _btb_309_bht_T_7 ? 2'h3 : _btb_309_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_25 = _btb_309_bht_T_5 ? 2'h3 : _btb_309_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_26 = _btb_309_bht_T_3 ? 2'h3 : _btb_309_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_309_bht_T_27 = _btb_309_bht_T_1 ? 2'h1 : _btb_309_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9942 = btb_309_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6965
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9944 = btb_309_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_309_bht_T_27 : _GEN_8501; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_310_bht_T = btb_310_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_310_bht_T_1 = io_i_branch_resolve_pack_taken & btb_310_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_310_bht_T_2 = btb_310_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_310_bht_T_3 = io_i_branch_resolve_pack_taken & btb_310_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_310_bht_T_4 = btb_310_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_310_bht_T_5 = io_i_branch_resolve_pack_taken & btb_310_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_310_bht_T_6 = btb_310_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_310_bht_T_7 = io_i_branch_resolve_pack_taken & btb_310_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_310_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_310_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_310_bht_T_13 = _btb_0_bht_T_8 & _btb_310_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_310_bht_T_16 = _btb_0_bht_T_8 & _btb_310_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_310_bht_T_19 = _btb_0_bht_T_8 & _btb_310_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_310_bht_T_20 = _btb_310_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_21 = _btb_310_bht_T_16 ? 2'h0 : _btb_310_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_22 = _btb_310_bht_T_13 ? 2'h0 : _btb_310_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_23 = _btb_310_bht_T_10 ? 2'h0 : _btb_310_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_24 = _btb_310_bht_T_7 ? 2'h3 : _btb_310_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_25 = _btb_310_bht_T_5 ? 2'h3 : _btb_310_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_26 = _btb_310_bht_T_3 ? 2'h3 : _btb_310_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_310_bht_T_27 = _btb_310_bht_T_1 ? 2'h1 : _btb_310_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9946 = btb_310_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6966
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9948 = btb_310_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_310_bht_T_27 : _GEN_8502; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_311_bht_T = btb_311_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_311_bht_T_1 = io_i_branch_resolve_pack_taken & btb_311_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_311_bht_T_2 = btb_311_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_311_bht_T_3 = io_i_branch_resolve_pack_taken & btb_311_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_311_bht_T_4 = btb_311_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_311_bht_T_5 = io_i_branch_resolve_pack_taken & btb_311_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_311_bht_T_6 = btb_311_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_311_bht_T_7 = io_i_branch_resolve_pack_taken & btb_311_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_311_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_311_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_311_bht_T_13 = _btb_0_bht_T_8 & _btb_311_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_311_bht_T_16 = _btb_0_bht_T_8 & _btb_311_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_311_bht_T_19 = _btb_0_bht_T_8 & _btb_311_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_311_bht_T_20 = _btb_311_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_21 = _btb_311_bht_T_16 ? 2'h0 : _btb_311_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_22 = _btb_311_bht_T_13 ? 2'h0 : _btb_311_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_23 = _btb_311_bht_T_10 ? 2'h0 : _btb_311_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_24 = _btb_311_bht_T_7 ? 2'h3 : _btb_311_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_25 = _btb_311_bht_T_5 ? 2'h3 : _btb_311_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_26 = _btb_311_bht_T_3 ? 2'h3 : _btb_311_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_311_bht_T_27 = _btb_311_bht_T_1 ? 2'h1 : _btb_311_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9950 = btb_311_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6967
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9952 = btb_311_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_311_bht_T_27 : _GEN_8503; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_312_bht_T = btb_312_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_312_bht_T_1 = io_i_branch_resolve_pack_taken & btb_312_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_312_bht_T_2 = btb_312_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_312_bht_T_3 = io_i_branch_resolve_pack_taken & btb_312_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_312_bht_T_4 = btb_312_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_312_bht_T_5 = io_i_branch_resolve_pack_taken & btb_312_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_312_bht_T_6 = btb_312_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_312_bht_T_7 = io_i_branch_resolve_pack_taken & btb_312_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_312_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_312_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_312_bht_T_13 = _btb_0_bht_T_8 & _btb_312_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_312_bht_T_16 = _btb_0_bht_T_8 & _btb_312_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_312_bht_T_19 = _btb_0_bht_T_8 & _btb_312_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_312_bht_T_20 = _btb_312_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_21 = _btb_312_bht_T_16 ? 2'h0 : _btb_312_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_22 = _btb_312_bht_T_13 ? 2'h0 : _btb_312_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_23 = _btb_312_bht_T_10 ? 2'h0 : _btb_312_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_24 = _btb_312_bht_T_7 ? 2'h3 : _btb_312_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_25 = _btb_312_bht_T_5 ? 2'h3 : _btb_312_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_26 = _btb_312_bht_T_3 ? 2'h3 : _btb_312_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_312_bht_T_27 = _btb_312_bht_T_1 ? 2'h1 : _btb_312_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9954 = btb_312_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6968
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9956 = btb_312_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_312_bht_T_27 : _GEN_8504; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_313_bht_T = btb_313_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_313_bht_T_1 = io_i_branch_resolve_pack_taken & btb_313_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_313_bht_T_2 = btb_313_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_313_bht_T_3 = io_i_branch_resolve_pack_taken & btb_313_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_313_bht_T_4 = btb_313_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_313_bht_T_5 = io_i_branch_resolve_pack_taken & btb_313_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_313_bht_T_6 = btb_313_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_313_bht_T_7 = io_i_branch_resolve_pack_taken & btb_313_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_313_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_313_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_313_bht_T_13 = _btb_0_bht_T_8 & _btb_313_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_313_bht_T_16 = _btb_0_bht_T_8 & _btb_313_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_313_bht_T_19 = _btb_0_bht_T_8 & _btb_313_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_313_bht_T_20 = _btb_313_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_21 = _btb_313_bht_T_16 ? 2'h0 : _btb_313_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_22 = _btb_313_bht_T_13 ? 2'h0 : _btb_313_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_23 = _btb_313_bht_T_10 ? 2'h0 : _btb_313_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_24 = _btb_313_bht_T_7 ? 2'h3 : _btb_313_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_25 = _btb_313_bht_T_5 ? 2'h3 : _btb_313_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_26 = _btb_313_bht_T_3 ? 2'h3 : _btb_313_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_313_bht_T_27 = _btb_313_bht_T_1 ? 2'h1 : _btb_313_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9958 = btb_313_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6969
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9960 = btb_313_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_313_bht_T_27 : _GEN_8505; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_314_bht_T = btb_314_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_314_bht_T_1 = io_i_branch_resolve_pack_taken & btb_314_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_314_bht_T_2 = btb_314_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_314_bht_T_3 = io_i_branch_resolve_pack_taken & btb_314_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_314_bht_T_4 = btb_314_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_314_bht_T_5 = io_i_branch_resolve_pack_taken & btb_314_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_314_bht_T_6 = btb_314_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_314_bht_T_7 = io_i_branch_resolve_pack_taken & btb_314_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_314_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_314_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_314_bht_T_13 = _btb_0_bht_T_8 & _btb_314_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_314_bht_T_16 = _btb_0_bht_T_8 & _btb_314_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_314_bht_T_19 = _btb_0_bht_T_8 & _btb_314_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_314_bht_T_20 = _btb_314_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_21 = _btb_314_bht_T_16 ? 2'h0 : _btb_314_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_22 = _btb_314_bht_T_13 ? 2'h0 : _btb_314_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_23 = _btb_314_bht_T_10 ? 2'h0 : _btb_314_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_24 = _btb_314_bht_T_7 ? 2'h3 : _btb_314_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_25 = _btb_314_bht_T_5 ? 2'h3 : _btb_314_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_26 = _btb_314_bht_T_3 ? 2'h3 : _btb_314_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_314_bht_T_27 = _btb_314_bht_T_1 ? 2'h1 : _btb_314_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_9961 = btb_314_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_313_tag == io_i_branch_resolve_pack_pc[12:3]
     | (btb_312_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_311_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_310_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_309_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_308_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_307_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_306_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_305_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_304_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_303_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_302_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_301_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_300_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9901)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_9962 = btb_314_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6970
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9964 = btb_314_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_314_bht_T_27 : _GEN_8506; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_315_bht_T = btb_315_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_315_bht_T_1 = io_i_branch_resolve_pack_taken & btb_315_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_315_bht_T_2 = btb_315_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_315_bht_T_3 = io_i_branch_resolve_pack_taken & btb_315_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_315_bht_T_4 = btb_315_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_315_bht_T_5 = io_i_branch_resolve_pack_taken & btb_315_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_315_bht_T_6 = btb_315_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_315_bht_T_7 = io_i_branch_resolve_pack_taken & btb_315_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_315_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_315_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_315_bht_T_13 = _btb_0_bht_T_8 & _btb_315_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_315_bht_T_16 = _btb_0_bht_T_8 & _btb_315_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_315_bht_T_19 = _btb_0_bht_T_8 & _btb_315_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_315_bht_T_20 = _btb_315_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_21 = _btb_315_bht_T_16 ? 2'h0 : _btb_315_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_22 = _btb_315_bht_T_13 ? 2'h0 : _btb_315_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_23 = _btb_315_bht_T_10 ? 2'h0 : _btb_315_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_24 = _btb_315_bht_T_7 ? 2'h3 : _btb_315_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_25 = _btb_315_bht_T_5 ? 2'h3 : _btb_315_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_26 = _btb_315_bht_T_3 ? 2'h3 : _btb_315_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_315_bht_T_27 = _btb_315_bht_T_1 ? 2'h1 : _btb_315_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9966 = btb_315_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6971
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9968 = btb_315_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_315_bht_T_27 : _GEN_8507; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_316_bht_T = btb_316_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_316_bht_T_1 = io_i_branch_resolve_pack_taken & btb_316_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_316_bht_T_2 = btb_316_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_316_bht_T_3 = io_i_branch_resolve_pack_taken & btb_316_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_316_bht_T_4 = btb_316_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_316_bht_T_5 = io_i_branch_resolve_pack_taken & btb_316_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_316_bht_T_6 = btb_316_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_316_bht_T_7 = io_i_branch_resolve_pack_taken & btb_316_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_316_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_316_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_316_bht_T_13 = _btb_0_bht_T_8 & _btb_316_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_316_bht_T_16 = _btb_0_bht_T_8 & _btb_316_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_316_bht_T_19 = _btb_0_bht_T_8 & _btb_316_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_316_bht_T_20 = _btb_316_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_21 = _btb_316_bht_T_16 ? 2'h0 : _btb_316_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_22 = _btb_316_bht_T_13 ? 2'h0 : _btb_316_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_23 = _btb_316_bht_T_10 ? 2'h0 : _btb_316_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_24 = _btb_316_bht_T_7 ? 2'h3 : _btb_316_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_25 = _btb_316_bht_T_5 ? 2'h3 : _btb_316_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_26 = _btb_316_bht_T_3 ? 2'h3 : _btb_316_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_316_bht_T_27 = _btb_316_bht_T_1 ? 2'h1 : _btb_316_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9970 = btb_316_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6972
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9972 = btb_316_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_316_bht_T_27 : _GEN_8508; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_317_bht_T = btb_317_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_317_bht_T_1 = io_i_branch_resolve_pack_taken & btb_317_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_317_bht_T_2 = btb_317_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_317_bht_T_3 = io_i_branch_resolve_pack_taken & btb_317_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_317_bht_T_4 = btb_317_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_317_bht_T_5 = io_i_branch_resolve_pack_taken & btb_317_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_317_bht_T_6 = btb_317_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_317_bht_T_7 = io_i_branch_resolve_pack_taken & btb_317_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_317_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_317_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_317_bht_T_13 = _btb_0_bht_T_8 & _btb_317_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_317_bht_T_16 = _btb_0_bht_T_8 & _btb_317_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_317_bht_T_19 = _btb_0_bht_T_8 & _btb_317_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_317_bht_T_20 = _btb_317_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_21 = _btb_317_bht_T_16 ? 2'h0 : _btb_317_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_22 = _btb_317_bht_T_13 ? 2'h0 : _btb_317_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_23 = _btb_317_bht_T_10 ? 2'h0 : _btb_317_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_24 = _btb_317_bht_T_7 ? 2'h3 : _btb_317_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_25 = _btb_317_bht_T_5 ? 2'h3 : _btb_317_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_26 = _btb_317_bht_T_3 ? 2'h3 : _btb_317_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_317_bht_T_27 = _btb_317_bht_T_1 ? 2'h1 : _btb_317_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9974 = btb_317_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6973
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9976 = btb_317_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_317_bht_T_27 : _GEN_8509; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_318_bht_T = btb_318_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_318_bht_T_1 = io_i_branch_resolve_pack_taken & btb_318_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_318_bht_T_2 = btb_318_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_318_bht_T_3 = io_i_branch_resolve_pack_taken & btb_318_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_318_bht_T_4 = btb_318_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_318_bht_T_5 = io_i_branch_resolve_pack_taken & btb_318_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_318_bht_T_6 = btb_318_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_318_bht_T_7 = io_i_branch_resolve_pack_taken & btb_318_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_318_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_318_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_318_bht_T_13 = _btb_0_bht_T_8 & _btb_318_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_318_bht_T_16 = _btb_0_bht_T_8 & _btb_318_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_318_bht_T_19 = _btb_0_bht_T_8 & _btb_318_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_318_bht_T_20 = _btb_318_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_21 = _btb_318_bht_T_16 ? 2'h0 : _btb_318_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_22 = _btb_318_bht_T_13 ? 2'h0 : _btb_318_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_23 = _btb_318_bht_T_10 ? 2'h0 : _btb_318_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_24 = _btb_318_bht_T_7 ? 2'h3 : _btb_318_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_25 = _btb_318_bht_T_5 ? 2'h3 : _btb_318_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_26 = _btb_318_bht_T_3 ? 2'h3 : _btb_318_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_318_bht_T_27 = _btb_318_bht_T_1 ? 2'h1 : _btb_318_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9978 = btb_318_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6974
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9980 = btb_318_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_318_bht_T_27 : _GEN_8510; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_319_bht_T = btb_319_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_319_bht_T_1 = io_i_branch_resolve_pack_taken & btb_319_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_319_bht_T_2 = btb_319_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_319_bht_T_3 = io_i_branch_resolve_pack_taken & btb_319_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_319_bht_T_4 = btb_319_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_319_bht_T_5 = io_i_branch_resolve_pack_taken & btb_319_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_319_bht_T_6 = btb_319_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_319_bht_T_7 = io_i_branch_resolve_pack_taken & btb_319_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_319_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_319_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_319_bht_T_13 = _btb_0_bht_T_8 & _btb_319_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_319_bht_T_16 = _btb_0_bht_T_8 & _btb_319_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_319_bht_T_19 = _btb_0_bht_T_8 & _btb_319_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_319_bht_T_20 = _btb_319_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_21 = _btb_319_bht_T_16 ? 2'h0 : _btb_319_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_22 = _btb_319_bht_T_13 ? 2'h0 : _btb_319_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_23 = _btb_319_bht_T_10 ? 2'h0 : _btb_319_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_24 = _btb_319_bht_T_7 ? 2'h3 : _btb_319_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_25 = _btb_319_bht_T_5 ? 2'h3 : _btb_319_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_26 = _btb_319_bht_T_3 ? 2'h3 : _btb_319_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_319_bht_T_27 = _btb_319_bht_T_1 ? 2'h1 : _btb_319_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9982 = btb_319_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6975
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9984 = btb_319_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_319_bht_T_27 : _GEN_8511; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_320_bht_T = btb_320_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_320_bht_T_1 = io_i_branch_resolve_pack_taken & btb_320_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_320_bht_T_2 = btb_320_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_320_bht_T_3 = io_i_branch_resolve_pack_taken & btb_320_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_320_bht_T_4 = btb_320_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_320_bht_T_5 = io_i_branch_resolve_pack_taken & btb_320_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_320_bht_T_6 = btb_320_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_320_bht_T_7 = io_i_branch_resolve_pack_taken & btb_320_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_320_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_320_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_320_bht_T_13 = _btb_0_bht_T_8 & _btb_320_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_320_bht_T_16 = _btb_0_bht_T_8 & _btb_320_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_320_bht_T_19 = _btb_0_bht_T_8 & _btb_320_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_320_bht_T_20 = _btb_320_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_21 = _btb_320_bht_T_16 ? 2'h0 : _btb_320_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_22 = _btb_320_bht_T_13 ? 2'h0 : _btb_320_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_23 = _btb_320_bht_T_10 ? 2'h0 : _btb_320_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_24 = _btb_320_bht_T_7 ? 2'h3 : _btb_320_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_25 = _btb_320_bht_T_5 ? 2'h3 : _btb_320_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_26 = _btb_320_bht_T_3 ? 2'h3 : _btb_320_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_320_bht_T_27 = _btb_320_bht_T_1 ? 2'h1 : _btb_320_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9986 = btb_320_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6976
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9988 = btb_320_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_320_bht_T_27 : _GEN_8512; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_321_bht_T = btb_321_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_321_bht_T_1 = io_i_branch_resolve_pack_taken & btb_321_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_321_bht_T_2 = btb_321_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_321_bht_T_3 = io_i_branch_resolve_pack_taken & btb_321_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_321_bht_T_4 = btb_321_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_321_bht_T_5 = io_i_branch_resolve_pack_taken & btb_321_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_321_bht_T_6 = btb_321_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_321_bht_T_7 = io_i_branch_resolve_pack_taken & btb_321_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_321_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_321_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_321_bht_T_13 = _btb_0_bht_T_8 & _btb_321_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_321_bht_T_16 = _btb_0_bht_T_8 & _btb_321_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_321_bht_T_19 = _btb_0_bht_T_8 & _btb_321_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_321_bht_T_20 = _btb_321_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_21 = _btb_321_bht_T_16 ? 2'h0 : _btb_321_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_22 = _btb_321_bht_T_13 ? 2'h0 : _btb_321_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_23 = _btb_321_bht_T_10 ? 2'h0 : _btb_321_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_24 = _btb_321_bht_T_7 ? 2'h3 : _btb_321_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_25 = _btb_321_bht_T_5 ? 2'h3 : _btb_321_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_26 = _btb_321_bht_T_3 ? 2'h3 : _btb_321_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_321_bht_T_27 = _btb_321_bht_T_1 ? 2'h1 : _btb_321_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9990 = btb_321_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6977
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9992 = btb_321_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_321_bht_T_27 : _GEN_8513; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_322_bht_T = btb_322_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_322_bht_T_1 = io_i_branch_resolve_pack_taken & btb_322_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_322_bht_T_2 = btb_322_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_322_bht_T_3 = io_i_branch_resolve_pack_taken & btb_322_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_322_bht_T_4 = btb_322_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_322_bht_T_5 = io_i_branch_resolve_pack_taken & btb_322_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_322_bht_T_6 = btb_322_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_322_bht_T_7 = io_i_branch_resolve_pack_taken & btb_322_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_322_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_322_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_322_bht_T_13 = _btb_0_bht_T_8 & _btb_322_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_322_bht_T_16 = _btb_0_bht_T_8 & _btb_322_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_322_bht_T_19 = _btb_0_bht_T_8 & _btb_322_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_322_bht_T_20 = _btb_322_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_21 = _btb_322_bht_T_16 ? 2'h0 : _btb_322_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_22 = _btb_322_bht_T_13 ? 2'h0 : _btb_322_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_23 = _btb_322_bht_T_10 ? 2'h0 : _btb_322_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_24 = _btb_322_bht_T_7 ? 2'h3 : _btb_322_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_25 = _btb_322_bht_T_5 ? 2'h3 : _btb_322_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_26 = _btb_322_bht_T_3 ? 2'h3 : _btb_322_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_322_bht_T_27 = _btb_322_bht_T_1 ? 2'h1 : _btb_322_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9994 = btb_322_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6978
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_9996 = btb_322_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_322_bht_T_27 : _GEN_8514; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_323_bht_T = btb_323_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_323_bht_T_1 = io_i_branch_resolve_pack_taken & btb_323_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_323_bht_T_2 = btb_323_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_323_bht_T_3 = io_i_branch_resolve_pack_taken & btb_323_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_323_bht_T_4 = btb_323_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_323_bht_T_5 = io_i_branch_resolve_pack_taken & btb_323_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_323_bht_T_6 = btb_323_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_323_bht_T_7 = io_i_branch_resolve_pack_taken & btb_323_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_323_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_323_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_323_bht_T_13 = _btb_0_bht_T_8 & _btb_323_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_323_bht_T_16 = _btb_0_bht_T_8 & _btb_323_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_323_bht_T_19 = _btb_0_bht_T_8 & _btb_323_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_323_bht_T_20 = _btb_323_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_21 = _btb_323_bht_T_16 ? 2'h0 : _btb_323_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_22 = _btb_323_bht_T_13 ? 2'h0 : _btb_323_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_23 = _btb_323_bht_T_10 ? 2'h0 : _btb_323_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_24 = _btb_323_bht_T_7 ? 2'h3 : _btb_323_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_25 = _btb_323_bht_T_5 ? 2'h3 : _btb_323_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_26 = _btb_323_bht_T_3 ? 2'h3 : _btb_323_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_323_bht_T_27 = _btb_323_bht_T_1 ? 2'h1 : _btb_323_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_9998 = btb_323_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target : _GEN_6979
    ; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10000 = btb_323_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_323_bht_T_27 : _GEN_8515; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_324_bht_T = btb_324_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_324_bht_T_1 = io_i_branch_resolve_pack_taken & btb_324_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_324_bht_T_2 = btb_324_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_324_bht_T_3 = io_i_branch_resolve_pack_taken & btb_324_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_324_bht_T_4 = btb_324_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_324_bht_T_5 = io_i_branch_resolve_pack_taken & btb_324_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_324_bht_T_6 = btb_324_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_324_bht_T_7 = io_i_branch_resolve_pack_taken & btb_324_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_324_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_324_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_324_bht_T_13 = _btb_0_bht_T_8 & _btb_324_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_324_bht_T_16 = _btb_0_bht_T_8 & _btb_324_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_324_bht_T_19 = _btb_0_bht_T_8 & _btb_324_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_324_bht_T_20 = _btb_324_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_21 = _btb_324_bht_T_16 ? 2'h0 : _btb_324_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_22 = _btb_324_bht_T_13 ? 2'h0 : _btb_324_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_23 = _btb_324_bht_T_10 ? 2'h0 : _btb_324_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_24 = _btb_324_bht_T_7 ? 2'h3 : _btb_324_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_25 = _btb_324_bht_T_5 ? 2'h3 : _btb_324_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_26 = _btb_324_bht_T_3 ? 2'h3 : _btb_324_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_324_bht_T_27 = _btb_324_bht_T_1 ? 2'h1 : _btb_324_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10002 = btb_324_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6980; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10004 = btb_324_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_324_bht_T_27 : _GEN_8516; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_325_bht_T = btb_325_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_325_bht_T_1 = io_i_branch_resolve_pack_taken & btb_325_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_325_bht_T_2 = btb_325_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_325_bht_T_3 = io_i_branch_resolve_pack_taken & btb_325_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_325_bht_T_4 = btb_325_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_325_bht_T_5 = io_i_branch_resolve_pack_taken & btb_325_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_325_bht_T_6 = btb_325_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_325_bht_T_7 = io_i_branch_resolve_pack_taken & btb_325_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_325_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_325_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_325_bht_T_13 = _btb_0_bht_T_8 & _btb_325_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_325_bht_T_16 = _btb_0_bht_T_8 & _btb_325_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_325_bht_T_19 = _btb_0_bht_T_8 & _btb_325_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_325_bht_T_20 = _btb_325_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_21 = _btb_325_bht_T_16 ? 2'h0 : _btb_325_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_22 = _btb_325_bht_T_13 ? 2'h0 : _btb_325_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_23 = _btb_325_bht_T_10 ? 2'h0 : _btb_325_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_24 = _btb_325_bht_T_7 ? 2'h3 : _btb_325_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_25 = _btb_325_bht_T_5 ? 2'h3 : _btb_325_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_26 = _btb_325_bht_T_3 ? 2'h3 : _btb_325_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_325_bht_T_27 = _btb_325_bht_T_1 ? 2'h1 : _btb_325_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10006 = btb_325_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6981; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10008 = btb_325_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_325_bht_T_27 : _GEN_8517; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_326_bht_T = btb_326_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_326_bht_T_1 = io_i_branch_resolve_pack_taken & btb_326_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_326_bht_T_2 = btb_326_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_326_bht_T_3 = io_i_branch_resolve_pack_taken & btb_326_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_326_bht_T_4 = btb_326_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_326_bht_T_5 = io_i_branch_resolve_pack_taken & btb_326_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_326_bht_T_6 = btb_326_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_326_bht_T_7 = io_i_branch_resolve_pack_taken & btb_326_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_326_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_326_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_326_bht_T_13 = _btb_0_bht_T_8 & _btb_326_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_326_bht_T_16 = _btb_0_bht_T_8 & _btb_326_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_326_bht_T_19 = _btb_0_bht_T_8 & _btb_326_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_326_bht_T_20 = _btb_326_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_21 = _btb_326_bht_T_16 ? 2'h0 : _btb_326_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_22 = _btb_326_bht_T_13 ? 2'h0 : _btb_326_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_23 = _btb_326_bht_T_10 ? 2'h0 : _btb_326_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_24 = _btb_326_bht_T_7 ? 2'h3 : _btb_326_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_25 = _btb_326_bht_T_5 ? 2'h3 : _btb_326_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_26 = _btb_326_bht_T_3 ? 2'h3 : _btb_326_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_326_bht_T_27 = _btb_326_bht_T_1 ? 2'h1 : _btb_326_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10010 = btb_326_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6982; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10012 = btb_326_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_326_bht_T_27 : _GEN_8518; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_327_bht_T = btb_327_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_327_bht_T_1 = io_i_branch_resolve_pack_taken & btb_327_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_327_bht_T_2 = btb_327_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_327_bht_T_3 = io_i_branch_resolve_pack_taken & btb_327_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_327_bht_T_4 = btb_327_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_327_bht_T_5 = io_i_branch_resolve_pack_taken & btb_327_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_327_bht_T_6 = btb_327_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_327_bht_T_7 = io_i_branch_resolve_pack_taken & btb_327_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_327_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_327_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_327_bht_T_13 = _btb_0_bht_T_8 & _btb_327_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_327_bht_T_16 = _btb_0_bht_T_8 & _btb_327_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_327_bht_T_19 = _btb_0_bht_T_8 & _btb_327_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_327_bht_T_20 = _btb_327_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_21 = _btb_327_bht_T_16 ? 2'h0 : _btb_327_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_22 = _btb_327_bht_T_13 ? 2'h0 : _btb_327_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_23 = _btb_327_bht_T_10 ? 2'h0 : _btb_327_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_24 = _btb_327_bht_T_7 ? 2'h3 : _btb_327_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_25 = _btb_327_bht_T_5 ? 2'h3 : _btb_327_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_26 = _btb_327_bht_T_3 ? 2'h3 : _btb_327_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_327_bht_T_27 = _btb_327_bht_T_1 ? 2'h1 : _btb_327_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10014 = btb_327_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6983; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10016 = btb_327_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_327_bht_T_27 : _GEN_8519; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_328_bht_T = btb_328_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_328_bht_T_1 = io_i_branch_resolve_pack_taken & btb_328_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_328_bht_T_2 = btb_328_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_328_bht_T_3 = io_i_branch_resolve_pack_taken & btb_328_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_328_bht_T_4 = btb_328_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_328_bht_T_5 = io_i_branch_resolve_pack_taken & btb_328_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_328_bht_T_6 = btb_328_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_328_bht_T_7 = io_i_branch_resolve_pack_taken & btb_328_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_328_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_328_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_328_bht_T_13 = _btb_0_bht_T_8 & _btb_328_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_328_bht_T_16 = _btb_0_bht_T_8 & _btb_328_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_328_bht_T_19 = _btb_0_bht_T_8 & _btb_328_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_328_bht_T_20 = _btb_328_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_21 = _btb_328_bht_T_16 ? 2'h0 : _btb_328_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_22 = _btb_328_bht_T_13 ? 2'h0 : _btb_328_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_23 = _btb_328_bht_T_10 ? 2'h0 : _btb_328_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_24 = _btb_328_bht_T_7 ? 2'h3 : _btb_328_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_25 = _btb_328_bht_T_5 ? 2'h3 : _btb_328_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_26 = _btb_328_bht_T_3 ? 2'h3 : _btb_328_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_328_bht_T_27 = _btb_328_bht_T_1 ? 2'h1 : _btb_328_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10018 = btb_328_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6984; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10020 = btb_328_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_328_bht_T_27 : _GEN_8520; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_329_bht_T = btb_329_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_329_bht_T_1 = io_i_branch_resolve_pack_taken & btb_329_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_329_bht_T_2 = btb_329_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_329_bht_T_3 = io_i_branch_resolve_pack_taken & btb_329_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_329_bht_T_4 = btb_329_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_329_bht_T_5 = io_i_branch_resolve_pack_taken & btb_329_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_329_bht_T_6 = btb_329_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_329_bht_T_7 = io_i_branch_resolve_pack_taken & btb_329_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_329_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_329_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_329_bht_T_13 = _btb_0_bht_T_8 & _btb_329_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_329_bht_T_16 = _btb_0_bht_T_8 & _btb_329_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_329_bht_T_19 = _btb_0_bht_T_8 & _btb_329_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_329_bht_T_20 = _btb_329_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_21 = _btb_329_bht_T_16 ? 2'h0 : _btb_329_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_22 = _btb_329_bht_T_13 ? 2'h0 : _btb_329_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_23 = _btb_329_bht_T_10 ? 2'h0 : _btb_329_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_24 = _btb_329_bht_T_7 ? 2'h3 : _btb_329_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_25 = _btb_329_bht_T_5 ? 2'h3 : _btb_329_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_26 = _btb_329_bht_T_3 ? 2'h3 : _btb_329_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_329_bht_T_27 = _btb_329_bht_T_1 ? 2'h1 : _btb_329_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10021 = btb_329_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_328_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_327_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_326_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_325_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_324_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_323_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_322_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_321_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_320_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_319_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_318_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_317_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_316_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_315_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_9961)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10022 = btb_329_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6985; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10024 = btb_329_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_329_bht_T_27 : _GEN_8521; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_330_bht_T = btb_330_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_330_bht_T_1 = io_i_branch_resolve_pack_taken & btb_330_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_330_bht_T_2 = btb_330_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_330_bht_T_3 = io_i_branch_resolve_pack_taken & btb_330_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_330_bht_T_4 = btb_330_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_330_bht_T_5 = io_i_branch_resolve_pack_taken & btb_330_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_330_bht_T_6 = btb_330_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_330_bht_T_7 = io_i_branch_resolve_pack_taken & btb_330_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_330_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_330_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_330_bht_T_13 = _btb_0_bht_T_8 & _btb_330_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_330_bht_T_16 = _btb_0_bht_T_8 & _btb_330_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_330_bht_T_19 = _btb_0_bht_T_8 & _btb_330_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_330_bht_T_20 = _btb_330_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_21 = _btb_330_bht_T_16 ? 2'h0 : _btb_330_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_22 = _btb_330_bht_T_13 ? 2'h0 : _btb_330_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_23 = _btb_330_bht_T_10 ? 2'h0 : _btb_330_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_24 = _btb_330_bht_T_7 ? 2'h3 : _btb_330_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_25 = _btb_330_bht_T_5 ? 2'h3 : _btb_330_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_26 = _btb_330_bht_T_3 ? 2'h3 : _btb_330_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_330_bht_T_27 = _btb_330_bht_T_1 ? 2'h1 : _btb_330_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10026 = btb_330_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6986; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10028 = btb_330_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_330_bht_T_27 : _GEN_8522; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_331_bht_T = btb_331_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_331_bht_T_1 = io_i_branch_resolve_pack_taken & btb_331_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_331_bht_T_2 = btb_331_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_331_bht_T_3 = io_i_branch_resolve_pack_taken & btb_331_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_331_bht_T_4 = btb_331_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_331_bht_T_5 = io_i_branch_resolve_pack_taken & btb_331_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_331_bht_T_6 = btb_331_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_331_bht_T_7 = io_i_branch_resolve_pack_taken & btb_331_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_331_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_331_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_331_bht_T_13 = _btb_0_bht_T_8 & _btb_331_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_331_bht_T_16 = _btb_0_bht_T_8 & _btb_331_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_331_bht_T_19 = _btb_0_bht_T_8 & _btb_331_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_331_bht_T_20 = _btb_331_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_21 = _btb_331_bht_T_16 ? 2'h0 : _btb_331_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_22 = _btb_331_bht_T_13 ? 2'h0 : _btb_331_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_23 = _btb_331_bht_T_10 ? 2'h0 : _btb_331_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_24 = _btb_331_bht_T_7 ? 2'h3 : _btb_331_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_25 = _btb_331_bht_T_5 ? 2'h3 : _btb_331_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_26 = _btb_331_bht_T_3 ? 2'h3 : _btb_331_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_331_bht_T_27 = _btb_331_bht_T_1 ? 2'h1 : _btb_331_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10030 = btb_331_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6987; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10032 = btb_331_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_331_bht_T_27 : _GEN_8523; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_332_bht_T = btb_332_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_332_bht_T_1 = io_i_branch_resolve_pack_taken & btb_332_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_332_bht_T_2 = btb_332_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_332_bht_T_3 = io_i_branch_resolve_pack_taken & btb_332_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_332_bht_T_4 = btb_332_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_332_bht_T_5 = io_i_branch_resolve_pack_taken & btb_332_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_332_bht_T_6 = btb_332_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_332_bht_T_7 = io_i_branch_resolve_pack_taken & btb_332_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_332_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_332_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_332_bht_T_13 = _btb_0_bht_T_8 & _btb_332_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_332_bht_T_16 = _btb_0_bht_T_8 & _btb_332_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_332_bht_T_19 = _btb_0_bht_T_8 & _btb_332_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_332_bht_T_20 = _btb_332_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_21 = _btb_332_bht_T_16 ? 2'h0 : _btb_332_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_22 = _btb_332_bht_T_13 ? 2'h0 : _btb_332_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_23 = _btb_332_bht_T_10 ? 2'h0 : _btb_332_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_24 = _btb_332_bht_T_7 ? 2'h3 : _btb_332_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_25 = _btb_332_bht_T_5 ? 2'h3 : _btb_332_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_26 = _btb_332_bht_T_3 ? 2'h3 : _btb_332_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_332_bht_T_27 = _btb_332_bht_T_1 ? 2'h1 : _btb_332_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10034 = btb_332_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6988; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10036 = btb_332_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_332_bht_T_27 : _GEN_8524; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_333_bht_T = btb_333_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_333_bht_T_1 = io_i_branch_resolve_pack_taken & btb_333_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_333_bht_T_2 = btb_333_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_333_bht_T_3 = io_i_branch_resolve_pack_taken & btb_333_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_333_bht_T_4 = btb_333_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_333_bht_T_5 = io_i_branch_resolve_pack_taken & btb_333_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_333_bht_T_6 = btb_333_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_333_bht_T_7 = io_i_branch_resolve_pack_taken & btb_333_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_333_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_333_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_333_bht_T_13 = _btb_0_bht_T_8 & _btb_333_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_333_bht_T_16 = _btb_0_bht_T_8 & _btb_333_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_333_bht_T_19 = _btb_0_bht_T_8 & _btb_333_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_333_bht_T_20 = _btb_333_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_21 = _btb_333_bht_T_16 ? 2'h0 : _btb_333_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_22 = _btb_333_bht_T_13 ? 2'h0 : _btb_333_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_23 = _btb_333_bht_T_10 ? 2'h0 : _btb_333_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_24 = _btb_333_bht_T_7 ? 2'h3 : _btb_333_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_25 = _btb_333_bht_T_5 ? 2'h3 : _btb_333_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_26 = _btb_333_bht_T_3 ? 2'h3 : _btb_333_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_333_bht_T_27 = _btb_333_bht_T_1 ? 2'h1 : _btb_333_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10038 = btb_333_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6989; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10040 = btb_333_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_333_bht_T_27 : _GEN_8525; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_334_bht_T = btb_334_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_334_bht_T_1 = io_i_branch_resolve_pack_taken & btb_334_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_334_bht_T_2 = btb_334_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_334_bht_T_3 = io_i_branch_resolve_pack_taken & btb_334_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_334_bht_T_4 = btb_334_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_334_bht_T_5 = io_i_branch_resolve_pack_taken & btb_334_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_334_bht_T_6 = btb_334_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_334_bht_T_7 = io_i_branch_resolve_pack_taken & btb_334_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_334_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_334_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_334_bht_T_13 = _btb_0_bht_T_8 & _btb_334_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_334_bht_T_16 = _btb_0_bht_T_8 & _btb_334_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_334_bht_T_19 = _btb_0_bht_T_8 & _btb_334_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_334_bht_T_20 = _btb_334_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_21 = _btb_334_bht_T_16 ? 2'h0 : _btb_334_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_22 = _btb_334_bht_T_13 ? 2'h0 : _btb_334_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_23 = _btb_334_bht_T_10 ? 2'h0 : _btb_334_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_24 = _btb_334_bht_T_7 ? 2'h3 : _btb_334_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_25 = _btb_334_bht_T_5 ? 2'h3 : _btb_334_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_26 = _btb_334_bht_T_3 ? 2'h3 : _btb_334_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_334_bht_T_27 = _btb_334_bht_T_1 ? 2'h1 : _btb_334_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10042 = btb_334_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6990; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10044 = btb_334_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_334_bht_T_27 : _GEN_8526; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_335_bht_T = btb_335_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_335_bht_T_1 = io_i_branch_resolve_pack_taken & btb_335_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_335_bht_T_2 = btb_335_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_335_bht_T_3 = io_i_branch_resolve_pack_taken & btb_335_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_335_bht_T_4 = btb_335_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_335_bht_T_5 = io_i_branch_resolve_pack_taken & btb_335_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_335_bht_T_6 = btb_335_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_335_bht_T_7 = io_i_branch_resolve_pack_taken & btb_335_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_335_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_335_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_335_bht_T_13 = _btb_0_bht_T_8 & _btb_335_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_335_bht_T_16 = _btb_0_bht_T_8 & _btb_335_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_335_bht_T_19 = _btb_0_bht_T_8 & _btb_335_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_335_bht_T_20 = _btb_335_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_21 = _btb_335_bht_T_16 ? 2'h0 : _btb_335_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_22 = _btb_335_bht_T_13 ? 2'h0 : _btb_335_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_23 = _btb_335_bht_T_10 ? 2'h0 : _btb_335_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_24 = _btb_335_bht_T_7 ? 2'h3 : _btb_335_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_25 = _btb_335_bht_T_5 ? 2'h3 : _btb_335_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_26 = _btb_335_bht_T_3 ? 2'h3 : _btb_335_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_335_bht_T_27 = _btb_335_bht_T_1 ? 2'h1 : _btb_335_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10046 = btb_335_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6991; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10048 = btb_335_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_335_bht_T_27 : _GEN_8527; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_336_bht_T = btb_336_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_336_bht_T_1 = io_i_branch_resolve_pack_taken & btb_336_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_336_bht_T_2 = btb_336_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_336_bht_T_3 = io_i_branch_resolve_pack_taken & btb_336_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_336_bht_T_4 = btb_336_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_336_bht_T_5 = io_i_branch_resolve_pack_taken & btb_336_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_336_bht_T_6 = btb_336_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_336_bht_T_7 = io_i_branch_resolve_pack_taken & btb_336_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_336_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_336_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_336_bht_T_13 = _btb_0_bht_T_8 & _btb_336_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_336_bht_T_16 = _btb_0_bht_T_8 & _btb_336_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_336_bht_T_19 = _btb_0_bht_T_8 & _btb_336_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_336_bht_T_20 = _btb_336_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_21 = _btb_336_bht_T_16 ? 2'h0 : _btb_336_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_22 = _btb_336_bht_T_13 ? 2'h0 : _btb_336_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_23 = _btb_336_bht_T_10 ? 2'h0 : _btb_336_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_24 = _btb_336_bht_T_7 ? 2'h3 : _btb_336_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_25 = _btb_336_bht_T_5 ? 2'h3 : _btb_336_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_26 = _btb_336_bht_T_3 ? 2'h3 : _btb_336_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_336_bht_T_27 = _btb_336_bht_T_1 ? 2'h1 : _btb_336_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10050 = btb_336_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6992; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10052 = btb_336_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_336_bht_T_27 : _GEN_8528; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_337_bht_T = btb_337_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_337_bht_T_1 = io_i_branch_resolve_pack_taken & btb_337_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_337_bht_T_2 = btb_337_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_337_bht_T_3 = io_i_branch_resolve_pack_taken & btb_337_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_337_bht_T_4 = btb_337_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_337_bht_T_5 = io_i_branch_resolve_pack_taken & btb_337_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_337_bht_T_6 = btb_337_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_337_bht_T_7 = io_i_branch_resolve_pack_taken & btb_337_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_337_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_337_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_337_bht_T_13 = _btb_0_bht_T_8 & _btb_337_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_337_bht_T_16 = _btb_0_bht_T_8 & _btb_337_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_337_bht_T_19 = _btb_0_bht_T_8 & _btb_337_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_337_bht_T_20 = _btb_337_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_21 = _btb_337_bht_T_16 ? 2'h0 : _btb_337_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_22 = _btb_337_bht_T_13 ? 2'h0 : _btb_337_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_23 = _btb_337_bht_T_10 ? 2'h0 : _btb_337_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_24 = _btb_337_bht_T_7 ? 2'h3 : _btb_337_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_25 = _btb_337_bht_T_5 ? 2'h3 : _btb_337_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_26 = _btb_337_bht_T_3 ? 2'h3 : _btb_337_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_337_bht_T_27 = _btb_337_bht_T_1 ? 2'h1 : _btb_337_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10054 = btb_337_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6993; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10056 = btb_337_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_337_bht_T_27 : _GEN_8529; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_338_bht_T = btb_338_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_338_bht_T_1 = io_i_branch_resolve_pack_taken & btb_338_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_338_bht_T_2 = btb_338_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_338_bht_T_3 = io_i_branch_resolve_pack_taken & btb_338_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_338_bht_T_4 = btb_338_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_338_bht_T_5 = io_i_branch_resolve_pack_taken & btb_338_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_338_bht_T_6 = btb_338_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_338_bht_T_7 = io_i_branch_resolve_pack_taken & btb_338_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_338_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_338_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_338_bht_T_13 = _btb_0_bht_T_8 & _btb_338_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_338_bht_T_16 = _btb_0_bht_T_8 & _btb_338_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_338_bht_T_19 = _btb_0_bht_T_8 & _btb_338_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_338_bht_T_20 = _btb_338_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_21 = _btb_338_bht_T_16 ? 2'h0 : _btb_338_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_22 = _btb_338_bht_T_13 ? 2'h0 : _btb_338_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_23 = _btb_338_bht_T_10 ? 2'h0 : _btb_338_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_24 = _btb_338_bht_T_7 ? 2'h3 : _btb_338_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_25 = _btb_338_bht_T_5 ? 2'h3 : _btb_338_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_26 = _btb_338_bht_T_3 ? 2'h3 : _btb_338_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_338_bht_T_27 = _btb_338_bht_T_1 ? 2'h1 : _btb_338_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10058 = btb_338_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6994; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10060 = btb_338_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_338_bht_T_27 : _GEN_8530; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_339_bht_T = btb_339_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_339_bht_T_1 = io_i_branch_resolve_pack_taken & btb_339_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_339_bht_T_2 = btb_339_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_339_bht_T_3 = io_i_branch_resolve_pack_taken & btb_339_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_339_bht_T_4 = btb_339_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_339_bht_T_5 = io_i_branch_resolve_pack_taken & btb_339_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_339_bht_T_6 = btb_339_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_339_bht_T_7 = io_i_branch_resolve_pack_taken & btb_339_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_339_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_339_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_339_bht_T_13 = _btb_0_bht_T_8 & _btb_339_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_339_bht_T_16 = _btb_0_bht_T_8 & _btb_339_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_339_bht_T_19 = _btb_0_bht_T_8 & _btb_339_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_339_bht_T_20 = _btb_339_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_21 = _btb_339_bht_T_16 ? 2'h0 : _btb_339_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_22 = _btb_339_bht_T_13 ? 2'h0 : _btb_339_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_23 = _btb_339_bht_T_10 ? 2'h0 : _btb_339_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_24 = _btb_339_bht_T_7 ? 2'h3 : _btb_339_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_25 = _btb_339_bht_T_5 ? 2'h3 : _btb_339_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_26 = _btb_339_bht_T_3 ? 2'h3 : _btb_339_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_339_bht_T_27 = _btb_339_bht_T_1 ? 2'h1 : _btb_339_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10062 = btb_339_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6995; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10064 = btb_339_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_339_bht_T_27 : _GEN_8531; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_340_bht_T = btb_340_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_340_bht_T_1 = io_i_branch_resolve_pack_taken & btb_340_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_340_bht_T_2 = btb_340_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_340_bht_T_3 = io_i_branch_resolve_pack_taken & btb_340_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_340_bht_T_4 = btb_340_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_340_bht_T_5 = io_i_branch_resolve_pack_taken & btb_340_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_340_bht_T_6 = btb_340_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_340_bht_T_7 = io_i_branch_resolve_pack_taken & btb_340_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_340_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_340_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_340_bht_T_13 = _btb_0_bht_T_8 & _btb_340_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_340_bht_T_16 = _btb_0_bht_T_8 & _btb_340_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_340_bht_T_19 = _btb_0_bht_T_8 & _btb_340_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_340_bht_T_20 = _btb_340_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_21 = _btb_340_bht_T_16 ? 2'h0 : _btb_340_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_22 = _btb_340_bht_T_13 ? 2'h0 : _btb_340_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_23 = _btb_340_bht_T_10 ? 2'h0 : _btb_340_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_24 = _btb_340_bht_T_7 ? 2'h3 : _btb_340_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_25 = _btb_340_bht_T_5 ? 2'h3 : _btb_340_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_26 = _btb_340_bht_T_3 ? 2'h3 : _btb_340_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_340_bht_T_27 = _btb_340_bht_T_1 ? 2'h1 : _btb_340_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10066 = btb_340_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6996; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10068 = btb_340_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_340_bht_T_27 : _GEN_8532; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_341_bht_T = btb_341_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_341_bht_T_1 = io_i_branch_resolve_pack_taken & btb_341_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_341_bht_T_2 = btb_341_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_341_bht_T_3 = io_i_branch_resolve_pack_taken & btb_341_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_341_bht_T_4 = btb_341_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_341_bht_T_5 = io_i_branch_resolve_pack_taken & btb_341_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_341_bht_T_6 = btb_341_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_341_bht_T_7 = io_i_branch_resolve_pack_taken & btb_341_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_341_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_341_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_341_bht_T_13 = _btb_0_bht_T_8 & _btb_341_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_341_bht_T_16 = _btb_0_bht_T_8 & _btb_341_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_341_bht_T_19 = _btb_0_bht_T_8 & _btb_341_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_341_bht_T_20 = _btb_341_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_21 = _btb_341_bht_T_16 ? 2'h0 : _btb_341_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_22 = _btb_341_bht_T_13 ? 2'h0 : _btb_341_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_23 = _btb_341_bht_T_10 ? 2'h0 : _btb_341_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_24 = _btb_341_bht_T_7 ? 2'h3 : _btb_341_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_25 = _btb_341_bht_T_5 ? 2'h3 : _btb_341_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_26 = _btb_341_bht_T_3 ? 2'h3 : _btb_341_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_341_bht_T_27 = _btb_341_bht_T_1 ? 2'h1 : _btb_341_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10070 = btb_341_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6997; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10072 = btb_341_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_341_bht_T_27 : _GEN_8533; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_342_bht_T = btb_342_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_342_bht_T_1 = io_i_branch_resolve_pack_taken & btb_342_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_342_bht_T_2 = btb_342_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_342_bht_T_3 = io_i_branch_resolve_pack_taken & btb_342_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_342_bht_T_4 = btb_342_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_342_bht_T_5 = io_i_branch_resolve_pack_taken & btb_342_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_342_bht_T_6 = btb_342_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_342_bht_T_7 = io_i_branch_resolve_pack_taken & btb_342_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_342_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_342_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_342_bht_T_13 = _btb_0_bht_T_8 & _btb_342_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_342_bht_T_16 = _btb_0_bht_T_8 & _btb_342_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_342_bht_T_19 = _btb_0_bht_T_8 & _btb_342_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_342_bht_T_20 = _btb_342_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_21 = _btb_342_bht_T_16 ? 2'h0 : _btb_342_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_22 = _btb_342_bht_T_13 ? 2'h0 : _btb_342_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_23 = _btb_342_bht_T_10 ? 2'h0 : _btb_342_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_24 = _btb_342_bht_T_7 ? 2'h3 : _btb_342_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_25 = _btb_342_bht_T_5 ? 2'h3 : _btb_342_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_26 = _btb_342_bht_T_3 ? 2'h3 : _btb_342_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_342_bht_T_27 = _btb_342_bht_T_1 ? 2'h1 : _btb_342_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10074 = btb_342_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6998; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10076 = btb_342_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_342_bht_T_27 : _GEN_8534; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_343_bht_T = btb_343_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_343_bht_T_1 = io_i_branch_resolve_pack_taken & btb_343_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_343_bht_T_2 = btb_343_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_343_bht_T_3 = io_i_branch_resolve_pack_taken & btb_343_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_343_bht_T_4 = btb_343_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_343_bht_T_5 = io_i_branch_resolve_pack_taken & btb_343_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_343_bht_T_6 = btb_343_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_343_bht_T_7 = io_i_branch_resolve_pack_taken & btb_343_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_343_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_343_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_343_bht_T_13 = _btb_0_bht_T_8 & _btb_343_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_343_bht_T_16 = _btb_0_bht_T_8 & _btb_343_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_343_bht_T_19 = _btb_0_bht_T_8 & _btb_343_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_343_bht_T_20 = _btb_343_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_21 = _btb_343_bht_T_16 ? 2'h0 : _btb_343_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_22 = _btb_343_bht_T_13 ? 2'h0 : _btb_343_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_23 = _btb_343_bht_T_10 ? 2'h0 : _btb_343_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_24 = _btb_343_bht_T_7 ? 2'h3 : _btb_343_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_25 = _btb_343_bht_T_5 ? 2'h3 : _btb_343_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_26 = _btb_343_bht_T_3 ? 2'h3 : _btb_343_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_343_bht_T_27 = _btb_343_bht_T_1 ? 2'h1 : _btb_343_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10078 = btb_343_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_6999; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10080 = btb_343_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_343_bht_T_27 : _GEN_8535; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_344_bht_T = btb_344_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_344_bht_T_1 = io_i_branch_resolve_pack_taken & btb_344_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_344_bht_T_2 = btb_344_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_344_bht_T_3 = io_i_branch_resolve_pack_taken & btb_344_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_344_bht_T_4 = btb_344_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_344_bht_T_5 = io_i_branch_resolve_pack_taken & btb_344_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_344_bht_T_6 = btb_344_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_344_bht_T_7 = io_i_branch_resolve_pack_taken & btb_344_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_344_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_344_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_344_bht_T_13 = _btb_0_bht_T_8 & _btb_344_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_344_bht_T_16 = _btb_0_bht_T_8 & _btb_344_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_344_bht_T_19 = _btb_0_bht_T_8 & _btb_344_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_344_bht_T_20 = _btb_344_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_21 = _btb_344_bht_T_16 ? 2'h0 : _btb_344_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_22 = _btb_344_bht_T_13 ? 2'h0 : _btb_344_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_23 = _btb_344_bht_T_10 ? 2'h0 : _btb_344_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_24 = _btb_344_bht_T_7 ? 2'h3 : _btb_344_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_25 = _btb_344_bht_T_5 ? 2'h3 : _btb_344_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_26 = _btb_344_bht_T_3 ? 2'h3 : _btb_344_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_344_bht_T_27 = _btb_344_bht_T_1 ? 2'h1 : _btb_344_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10081 = btb_344_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_343_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_342_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_341_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_340_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_339_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_338_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_337_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_336_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_335_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_334_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_333_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_332_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_331_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_330_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10021)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10082 = btb_344_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7000; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10084 = btb_344_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_344_bht_T_27 : _GEN_8536; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_345_bht_T = btb_345_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_345_bht_T_1 = io_i_branch_resolve_pack_taken & btb_345_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_345_bht_T_2 = btb_345_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_345_bht_T_3 = io_i_branch_resolve_pack_taken & btb_345_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_345_bht_T_4 = btb_345_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_345_bht_T_5 = io_i_branch_resolve_pack_taken & btb_345_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_345_bht_T_6 = btb_345_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_345_bht_T_7 = io_i_branch_resolve_pack_taken & btb_345_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_345_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_345_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_345_bht_T_13 = _btb_0_bht_T_8 & _btb_345_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_345_bht_T_16 = _btb_0_bht_T_8 & _btb_345_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_345_bht_T_19 = _btb_0_bht_T_8 & _btb_345_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_345_bht_T_20 = _btb_345_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_21 = _btb_345_bht_T_16 ? 2'h0 : _btb_345_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_22 = _btb_345_bht_T_13 ? 2'h0 : _btb_345_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_23 = _btb_345_bht_T_10 ? 2'h0 : _btb_345_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_24 = _btb_345_bht_T_7 ? 2'h3 : _btb_345_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_25 = _btb_345_bht_T_5 ? 2'h3 : _btb_345_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_26 = _btb_345_bht_T_3 ? 2'h3 : _btb_345_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_345_bht_T_27 = _btb_345_bht_T_1 ? 2'h1 : _btb_345_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10086 = btb_345_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7001; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10088 = btb_345_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_345_bht_T_27 : _GEN_8537; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_346_bht_T = btb_346_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_346_bht_T_1 = io_i_branch_resolve_pack_taken & btb_346_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_346_bht_T_2 = btb_346_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_346_bht_T_3 = io_i_branch_resolve_pack_taken & btb_346_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_346_bht_T_4 = btb_346_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_346_bht_T_5 = io_i_branch_resolve_pack_taken & btb_346_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_346_bht_T_6 = btb_346_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_346_bht_T_7 = io_i_branch_resolve_pack_taken & btb_346_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_346_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_346_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_346_bht_T_13 = _btb_0_bht_T_8 & _btb_346_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_346_bht_T_16 = _btb_0_bht_T_8 & _btb_346_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_346_bht_T_19 = _btb_0_bht_T_8 & _btb_346_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_346_bht_T_20 = _btb_346_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_21 = _btb_346_bht_T_16 ? 2'h0 : _btb_346_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_22 = _btb_346_bht_T_13 ? 2'h0 : _btb_346_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_23 = _btb_346_bht_T_10 ? 2'h0 : _btb_346_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_24 = _btb_346_bht_T_7 ? 2'h3 : _btb_346_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_25 = _btb_346_bht_T_5 ? 2'h3 : _btb_346_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_26 = _btb_346_bht_T_3 ? 2'h3 : _btb_346_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_346_bht_T_27 = _btb_346_bht_T_1 ? 2'h1 : _btb_346_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10090 = btb_346_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7002; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10092 = btb_346_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_346_bht_T_27 : _GEN_8538; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_347_bht_T = btb_347_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_347_bht_T_1 = io_i_branch_resolve_pack_taken & btb_347_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_347_bht_T_2 = btb_347_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_347_bht_T_3 = io_i_branch_resolve_pack_taken & btb_347_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_347_bht_T_4 = btb_347_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_347_bht_T_5 = io_i_branch_resolve_pack_taken & btb_347_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_347_bht_T_6 = btb_347_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_347_bht_T_7 = io_i_branch_resolve_pack_taken & btb_347_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_347_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_347_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_347_bht_T_13 = _btb_0_bht_T_8 & _btb_347_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_347_bht_T_16 = _btb_0_bht_T_8 & _btb_347_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_347_bht_T_19 = _btb_0_bht_T_8 & _btb_347_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_347_bht_T_20 = _btb_347_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_21 = _btb_347_bht_T_16 ? 2'h0 : _btb_347_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_22 = _btb_347_bht_T_13 ? 2'h0 : _btb_347_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_23 = _btb_347_bht_T_10 ? 2'h0 : _btb_347_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_24 = _btb_347_bht_T_7 ? 2'h3 : _btb_347_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_25 = _btb_347_bht_T_5 ? 2'h3 : _btb_347_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_26 = _btb_347_bht_T_3 ? 2'h3 : _btb_347_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_347_bht_T_27 = _btb_347_bht_T_1 ? 2'h1 : _btb_347_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10094 = btb_347_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7003; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10096 = btb_347_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_347_bht_T_27 : _GEN_8539; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_348_bht_T = btb_348_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_348_bht_T_1 = io_i_branch_resolve_pack_taken & btb_348_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_348_bht_T_2 = btb_348_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_348_bht_T_3 = io_i_branch_resolve_pack_taken & btb_348_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_348_bht_T_4 = btb_348_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_348_bht_T_5 = io_i_branch_resolve_pack_taken & btb_348_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_348_bht_T_6 = btb_348_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_348_bht_T_7 = io_i_branch_resolve_pack_taken & btb_348_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_348_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_348_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_348_bht_T_13 = _btb_0_bht_T_8 & _btb_348_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_348_bht_T_16 = _btb_0_bht_T_8 & _btb_348_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_348_bht_T_19 = _btb_0_bht_T_8 & _btb_348_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_348_bht_T_20 = _btb_348_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_21 = _btb_348_bht_T_16 ? 2'h0 : _btb_348_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_22 = _btb_348_bht_T_13 ? 2'h0 : _btb_348_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_23 = _btb_348_bht_T_10 ? 2'h0 : _btb_348_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_24 = _btb_348_bht_T_7 ? 2'h3 : _btb_348_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_25 = _btb_348_bht_T_5 ? 2'h3 : _btb_348_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_26 = _btb_348_bht_T_3 ? 2'h3 : _btb_348_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_348_bht_T_27 = _btb_348_bht_T_1 ? 2'h1 : _btb_348_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10098 = btb_348_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7004; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10100 = btb_348_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_348_bht_T_27 : _GEN_8540; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_349_bht_T = btb_349_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_349_bht_T_1 = io_i_branch_resolve_pack_taken & btb_349_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_349_bht_T_2 = btb_349_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_349_bht_T_3 = io_i_branch_resolve_pack_taken & btb_349_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_349_bht_T_4 = btb_349_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_349_bht_T_5 = io_i_branch_resolve_pack_taken & btb_349_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_349_bht_T_6 = btb_349_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_349_bht_T_7 = io_i_branch_resolve_pack_taken & btb_349_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_349_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_349_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_349_bht_T_13 = _btb_0_bht_T_8 & _btb_349_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_349_bht_T_16 = _btb_0_bht_T_8 & _btb_349_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_349_bht_T_19 = _btb_0_bht_T_8 & _btb_349_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_349_bht_T_20 = _btb_349_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_21 = _btb_349_bht_T_16 ? 2'h0 : _btb_349_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_22 = _btb_349_bht_T_13 ? 2'h0 : _btb_349_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_23 = _btb_349_bht_T_10 ? 2'h0 : _btb_349_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_24 = _btb_349_bht_T_7 ? 2'h3 : _btb_349_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_25 = _btb_349_bht_T_5 ? 2'h3 : _btb_349_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_26 = _btb_349_bht_T_3 ? 2'h3 : _btb_349_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_349_bht_T_27 = _btb_349_bht_T_1 ? 2'h1 : _btb_349_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10102 = btb_349_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7005; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10104 = btb_349_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_349_bht_T_27 : _GEN_8541; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_350_bht_T = btb_350_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_350_bht_T_1 = io_i_branch_resolve_pack_taken & btb_350_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_350_bht_T_2 = btb_350_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_350_bht_T_3 = io_i_branch_resolve_pack_taken & btb_350_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_350_bht_T_4 = btb_350_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_350_bht_T_5 = io_i_branch_resolve_pack_taken & btb_350_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_350_bht_T_6 = btb_350_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_350_bht_T_7 = io_i_branch_resolve_pack_taken & btb_350_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_350_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_350_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_350_bht_T_13 = _btb_0_bht_T_8 & _btb_350_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_350_bht_T_16 = _btb_0_bht_T_8 & _btb_350_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_350_bht_T_19 = _btb_0_bht_T_8 & _btb_350_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_350_bht_T_20 = _btb_350_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_21 = _btb_350_bht_T_16 ? 2'h0 : _btb_350_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_22 = _btb_350_bht_T_13 ? 2'h0 : _btb_350_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_23 = _btb_350_bht_T_10 ? 2'h0 : _btb_350_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_24 = _btb_350_bht_T_7 ? 2'h3 : _btb_350_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_25 = _btb_350_bht_T_5 ? 2'h3 : _btb_350_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_26 = _btb_350_bht_T_3 ? 2'h3 : _btb_350_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_350_bht_T_27 = _btb_350_bht_T_1 ? 2'h1 : _btb_350_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10106 = btb_350_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7006; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10108 = btb_350_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_350_bht_T_27 : _GEN_8542; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_351_bht_T = btb_351_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_351_bht_T_1 = io_i_branch_resolve_pack_taken & btb_351_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_351_bht_T_2 = btb_351_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_351_bht_T_3 = io_i_branch_resolve_pack_taken & btb_351_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_351_bht_T_4 = btb_351_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_351_bht_T_5 = io_i_branch_resolve_pack_taken & btb_351_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_351_bht_T_6 = btb_351_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_351_bht_T_7 = io_i_branch_resolve_pack_taken & btb_351_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_351_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_351_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_351_bht_T_13 = _btb_0_bht_T_8 & _btb_351_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_351_bht_T_16 = _btb_0_bht_T_8 & _btb_351_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_351_bht_T_19 = _btb_0_bht_T_8 & _btb_351_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_351_bht_T_20 = _btb_351_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_21 = _btb_351_bht_T_16 ? 2'h0 : _btb_351_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_22 = _btb_351_bht_T_13 ? 2'h0 : _btb_351_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_23 = _btb_351_bht_T_10 ? 2'h0 : _btb_351_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_24 = _btb_351_bht_T_7 ? 2'h3 : _btb_351_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_25 = _btb_351_bht_T_5 ? 2'h3 : _btb_351_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_26 = _btb_351_bht_T_3 ? 2'h3 : _btb_351_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_351_bht_T_27 = _btb_351_bht_T_1 ? 2'h1 : _btb_351_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10110 = btb_351_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7007; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10112 = btb_351_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_351_bht_T_27 : _GEN_8543; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_352_bht_T = btb_352_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_352_bht_T_1 = io_i_branch_resolve_pack_taken & btb_352_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_352_bht_T_2 = btb_352_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_352_bht_T_3 = io_i_branch_resolve_pack_taken & btb_352_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_352_bht_T_4 = btb_352_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_352_bht_T_5 = io_i_branch_resolve_pack_taken & btb_352_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_352_bht_T_6 = btb_352_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_352_bht_T_7 = io_i_branch_resolve_pack_taken & btb_352_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_352_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_352_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_352_bht_T_13 = _btb_0_bht_T_8 & _btb_352_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_352_bht_T_16 = _btb_0_bht_T_8 & _btb_352_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_352_bht_T_19 = _btb_0_bht_T_8 & _btb_352_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_352_bht_T_20 = _btb_352_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_21 = _btb_352_bht_T_16 ? 2'h0 : _btb_352_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_22 = _btb_352_bht_T_13 ? 2'h0 : _btb_352_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_23 = _btb_352_bht_T_10 ? 2'h0 : _btb_352_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_24 = _btb_352_bht_T_7 ? 2'h3 : _btb_352_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_25 = _btb_352_bht_T_5 ? 2'h3 : _btb_352_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_26 = _btb_352_bht_T_3 ? 2'h3 : _btb_352_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_352_bht_T_27 = _btb_352_bht_T_1 ? 2'h1 : _btb_352_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10114 = btb_352_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7008; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10116 = btb_352_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_352_bht_T_27 : _GEN_8544; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_353_bht_T = btb_353_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_353_bht_T_1 = io_i_branch_resolve_pack_taken & btb_353_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_353_bht_T_2 = btb_353_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_353_bht_T_3 = io_i_branch_resolve_pack_taken & btb_353_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_353_bht_T_4 = btb_353_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_353_bht_T_5 = io_i_branch_resolve_pack_taken & btb_353_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_353_bht_T_6 = btb_353_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_353_bht_T_7 = io_i_branch_resolve_pack_taken & btb_353_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_353_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_353_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_353_bht_T_13 = _btb_0_bht_T_8 & _btb_353_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_353_bht_T_16 = _btb_0_bht_T_8 & _btb_353_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_353_bht_T_19 = _btb_0_bht_T_8 & _btb_353_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_353_bht_T_20 = _btb_353_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_21 = _btb_353_bht_T_16 ? 2'h0 : _btb_353_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_22 = _btb_353_bht_T_13 ? 2'h0 : _btb_353_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_23 = _btb_353_bht_T_10 ? 2'h0 : _btb_353_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_24 = _btb_353_bht_T_7 ? 2'h3 : _btb_353_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_25 = _btb_353_bht_T_5 ? 2'h3 : _btb_353_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_26 = _btb_353_bht_T_3 ? 2'h3 : _btb_353_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_353_bht_T_27 = _btb_353_bht_T_1 ? 2'h1 : _btb_353_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10118 = btb_353_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7009; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10120 = btb_353_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_353_bht_T_27 : _GEN_8545; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_354_bht_T = btb_354_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_354_bht_T_1 = io_i_branch_resolve_pack_taken & btb_354_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_354_bht_T_2 = btb_354_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_354_bht_T_3 = io_i_branch_resolve_pack_taken & btb_354_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_354_bht_T_4 = btb_354_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_354_bht_T_5 = io_i_branch_resolve_pack_taken & btb_354_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_354_bht_T_6 = btb_354_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_354_bht_T_7 = io_i_branch_resolve_pack_taken & btb_354_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_354_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_354_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_354_bht_T_13 = _btb_0_bht_T_8 & _btb_354_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_354_bht_T_16 = _btb_0_bht_T_8 & _btb_354_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_354_bht_T_19 = _btb_0_bht_T_8 & _btb_354_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_354_bht_T_20 = _btb_354_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_21 = _btb_354_bht_T_16 ? 2'h0 : _btb_354_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_22 = _btb_354_bht_T_13 ? 2'h0 : _btb_354_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_23 = _btb_354_bht_T_10 ? 2'h0 : _btb_354_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_24 = _btb_354_bht_T_7 ? 2'h3 : _btb_354_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_25 = _btb_354_bht_T_5 ? 2'h3 : _btb_354_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_26 = _btb_354_bht_T_3 ? 2'h3 : _btb_354_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_354_bht_T_27 = _btb_354_bht_T_1 ? 2'h1 : _btb_354_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10122 = btb_354_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7010; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10124 = btb_354_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_354_bht_T_27 : _GEN_8546; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_355_bht_T = btb_355_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_355_bht_T_1 = io_i_branch_resolve_pack_taken & btb_355_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_355_bht_T_2 = btb_355_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_355_bht_T_3 = io_i_branch_resolve_pack_taken & btb_355_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_355_bht_T_4 = btb_355_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_355_bht_T_5 = io_i_branch_resolve_pack_taken & btb_355_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_355_bht_T_6 = btb_355_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_355_bht_T_7 = io_i_branch_resolve_pack_taken & btb_355_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_355_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_355_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_355_bht_T_13 = _btb_0_bht_T_8 & _btb_355_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_355_bht_T_16 = _btb_0_bht_T_8 & _btb_355_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_355_bht_T_19 = _btb_0_bht_T_8 & _btb_355_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_355_bht_T_20 = _btb_355_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_21 = _btb_355_bht_T_16 ? 2'h0 : _btb_355_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_22 = _btb_355_bht_T_13 ? 2'h0 : _btb_355_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_23 = _btb_355_bht_T_10 ? 2'h0 : _btb_355_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_24 = _btb_355_bht_T_7 ? 2'h3 : _btb_355_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_25 = _btb_355_bht_T_5 ? 2'h3 : _btb_355_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_26 = _btb_355_bht_T_3 ? 2'h3 : _btb_355_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_355_bht_T_27 = _btb_355_bht_T_1 ? 2'h1 : _btb_355_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10126 = btb_355_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7011; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10128 = btb_355_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_355_bht_T_27 : _GEN_8547; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_356_bht_T = btb_356_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_356_bht_T_1 = io_i_branch_resolve_pack_taken & btb_356_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_356_bht_T_2 = btb_356_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_356_bht_T_3 = io_i_branch_resolve_pack_taken & btb_356_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_356_bht_T_4 = btb_356_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_356_bht_T_5 = io_i_branch_resolve_pack_taken & btb_356_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_356_bht_T_6 = btb_356_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_356_bht_T_7 = io_i_branch_resolve_pack_taken & btb_356_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_356_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_356_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_356_bht_T_13 = _btb_0_bht_T_8 & _btb_356_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_356_bht_T_16 = _btb_0_bht_T_8 & _btb_356_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_356_bht_T_19 = _btb_0_bht_T_8 & _btb_356_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_356_bht_T_20 = _btb_356_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_21 = _btb_356_bht_T_16 ? 2'h0 : _btb_356_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_22 = _btb_356_bht_T_13 ? 2'h0 : _btb_356_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_23 = _btb_356_bht_T_10 ? 2'h0 : _btb_356_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_24 = _btb_356_bht_T_7 ? 2'h3 : _btb_356_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_25 = _btb_356_bht_T_5 ? 2'h3 : _btb_356_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_26 = _btb_356_bht_T_3 ? 2'h3 : _btb_356_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_356_bht_T_27 = _btb_356_bht_T_1 ? 2'h1 : _btb_356_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10130 = btb_356_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7012; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10132 = btb_356_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_356_bht_T_27 : _GEN_8548; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_357_bht_T = btb_357_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_357_bht_T_1 = io_i_branch_resolve_pack_taken & btb_357_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_357_bht_T_2 = btb_357_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_357_bht_T_3 = io_i_branch_resolve_pack_taken & btb_357_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_357_bht_T_4 = btb_357_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_357_bht_T_5 = io_i_branch_resolve_pack_taken & btb_357_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_357_bht_T_6 = btb_357_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_357_bht_T_7 = io_i_branch_resolve_pack_taken & btb_357_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_357_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_357_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_357_bht_T_13 = _btb_0_bht_T_8 & _btb_357_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_357_bht_T_16 = _btb_0_bht_T_8 & _btb_357_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_357_bht_T_19 = _btb_0_bht_T_8 & _btb_357_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_357_bht_T_20 = _btb_357_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_21 = _btb_357_bht_T_16 ? 2'h0 : _btb_357_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_22 = _btb_357_bht_T_13 ? 2'h0 : _btb_357_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_23 = _btb_357_bht_T_10 ? 2'h0 : _btb_357_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_24 = _btb_357_bht_T_7 ? 2'h3 : _btb_357_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_25 = _btb_357_bht_T_5 ? 2'h3 : _btb_357_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_26 = _btb_357_bht_T_3 ? 2'h3 : _btb_357_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_357_bht_T_27 = _btb_357_bht_T_1 ? 2'h1 : _btb_357_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10134 = btb_357_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7013; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10136 = btb_357_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_357_bht_T_27 : _GEN_8549; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_358_bht_T = btb_358_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_358_bht_T_1 = io_i_branch_resolve_pack_taken & btb_358_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_358_bht_T_2 = btb_358_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_358_bht_T_3 = io_i_branch_resolve_pack_taken & btb_358_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_358_bht_T_4 = btb_358_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_358_bht_T_5 = io_i_branch_resolve_pack_taken & btb_358_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_358_bht_T_6 = btb_358_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_358_bht_T_7 = io_i_branch_resolve_pack_taken & btb_358_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_358_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_358_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_358_bht_T_13 = _btb_0_bht_T_8 & _btb_358_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_358_bht_T_16 = _btb_0_bht_T_8 & _btb_358_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_358_bht_T_19 = _btb_0_bht_T_8 & _btb_358_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_358_bht_T_20 = _btb_358_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_21 = _btb_358_bht_T_16 ? 2'h0 : _btb_358_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_22 = _btb_358_bht_T_13 ? 2'h0 : _btb_358_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_23 = _btb_358_bht_T_10 ? 2'h0 : _btb_358_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_24 = _btb_358_bht_T_7 ? 2'h3 : _btb_358_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_25 = _btb_358_bht_T_5 ? 2'h3 : _btb_358_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_26 = _btb_358_bht_T_3 ? 2'h3 : _btb_358_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_358_bht_T_27 = _btb_358_bht_T_1 ? 2'h1 : _btb_358_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10138 = btb_358_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7014; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10140 = btb_358_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_358_bht_T_27 : _GEN_8550; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_359_bht_T = btb_359_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_359_bht_T_1 = io_i_branch_resolve_pack_taken & btb_359_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_359_bht_T_2 = btb_359_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_359_bht_T_3 = io_i_branch_resolve_pack_taken & btb_359_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_359_bht_T_4 = btb_359_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_359_bht_T_5 = io_i_branch_resolve_pack_taken & btb_359_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_359_bht_T_6 = btb_359_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_359_bht_T_7 = io_i_branch_resolve_pack_taken & btb_359_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_359_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_359_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_359_bht_T_13 = _btb_0_bht_T_8 & _btb_359_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_359_bht_T_16 = _btb_0_bht_T_8 & _btb_359_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_359_bht_T_19 = _btb_0_bht_T_8 & _btb_359_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_359_bht_T_20 = _btb_359_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_21 = _btb_359_bht_T_16 ? 2'h0 : _btb_359_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_22 = _btb_359_bht_T_13 ? 2'h0 : _btb_359_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_23 = _btb_359_bht_T_10 ? 2'h0 : _btb_359_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_24 = _btb_359_bht_T_7 ? 2'h3 : _btb_359_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_25 = _btb_359_bht_T_5 ? 2'h3 : _btb_359_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_26 = _btb_359_bht_T_3 ? 2'h3 : _btb_359_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_359_bht_T_27 = _btb_359_bht_T_1 ? 2'h1 : _btb_359_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10141 = btb_359_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_358_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_357_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_356_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_355_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_354_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_353_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_352_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_351_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_350_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_349_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_348_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_347_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_346_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_345_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10081)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10142 = btb_359_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7015; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10144 = btb_359_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_359_bht_T_27 : _GEN_8551; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_360_bht_T = btb_360_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_360_bht_T_1 = io_i_branch_resolve_pack_taken & btb_360_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_360_bht_T_2 = btb_360_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_360_bht_T_3 = io_i_branch_resolve_pack_taken & btb_360_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_360_bht_T_4 = btb_360_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_360_bht_T_5 = io_i_branch_resolve_pack_taken & btb_360_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_360_bht_T_6 = btb_360_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_360_bht_T_7 = io_i_branch_resolve_pack_taken & btb_360_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_360_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_360_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_360_bht_T_13 = _btb_0_bht_T_8 & _btb_360_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_360_bht_T_16 = _btb_0_bht_T_8 & _btb_360_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_360_bht_T_19 = _btb_0_bht_T_8 & _btb_360_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_360_bht_T_20 = _btb_360_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_21 = _btb_360_bht_T_16 ? 2'h0 : _btb_360_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_22 = _btb_360_bht_T_13 ? 2'h0 : _btb_360_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_23 = _btb_360_bht_T_10 ? 2'h0 : _btb_360_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_24 = _btb_360_bht_T_7 ? 2'h3 : _btb_360_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_25 = _btb_360_bht_T_5 ? 2'h3 : _btb_360_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_26 = _btb_360_bht_T_3 ? 2'h3 : _btb_360_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_360_bht_T_27 = _btb_360_bht_T_1 ? 2'h1 : _btb_360_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10146 = btb_360_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7016; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10148 = btb_360_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_360_bht_T_27 : _GEN_8552; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_361_bht_T = btb_361_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_361_bht_T_1 = io_i_branch_resolve_pack_taken & btb_361_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_361_bht_T_2 = btb_361_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_361_bht_T_3 = io_i_branch_resolve_pack_taken & btb_361_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_361_bht_T_4 = btb_361_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_361_bht_T_5 = io_i_branch_resolve_pack_taken & btb_361_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_361_bht_T_6 = btb_361_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_361_bht_T_7 = io_i_branch_resolve_pack_taken & btb_361_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_361_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_361_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_361_bht_T_13 = _btb_0_bht_T_8 & _btb_361_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_361_bht_T_16 = _btb_0_bht_T_8 & _btb_361_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_361_bht_T_19 = _btb_0_bht_T_8 & _btb_361_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_361_bht_T_20 = _btb_361_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_21 = _btb_361_bht_T_16 ? 2'h0 : _btb_361_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_22 = _btb_361_bht_T_13 ? 2'h0 : _btb_361_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_23 = _btb_361_bht_T_10 ? 2'h0 : _btb_361_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_24 = _btb_361_bht_T_7 ? 2'h3 : _btb_361_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_25 = _btb_361_bht_T_5 ? 2'h3 : _btb_361_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_26 = _btb_361_bht_T_3 ? 2'h3 : _btb_361_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_361_bht_T_27 = _btb_361_bht_T_1 ? 2'h1 : _btb_361_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10150 = btb_361_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7017; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10152 = btb_361_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_361_bht_T_27 : _GEN_8553; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_362_bht_T = btb_362_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_362_bht_T_1 = io_i_branch_resolve_pack_taken & btb_362_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_362_bht_T_2 = btb_362_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_362_bht_T_3 = io_i_branch_resolve_pack_taken & btb_362_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_362_bht_T_4 = btb_362_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_362_bht_T_5 = io_i_branch_resolve_pack_taken & btb_362_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_362_bht_T_6 = btb_362_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_362_bht_T_7 = io_i_branch_resolve_pack_taken & btb_362_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_362_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_362_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_362_bht_T_13 = _btb_0_bht_T_8 & _btb_362_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_362_bht_T_16 = _btb_0_bht_T_8 & _btb_362_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_362_bht_T_19 = _btb_0_bht_T_8 & _btb_362_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_362_bht_T_20 = _btb_362_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_21 = _btb_362_bht_T_16 ? 2'h0 : _btb_362_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_22 = _btb_362_bht_T_13 ? 2'h0 : _btb_362_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_23 = _btb_362_bht_T_10 ? 2'h0 : _btb_362_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_24 = _btb_362_bht_T_7 ? 2'h3 : _btb_362_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_25 = _btb_362_bht_T_5 ? 2'h3 : _btb_362_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_26 = _btb_362_bht_T_3 ? 2'h3 : _btb_362_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_362_bht_T_27 = _btb_362_bht_T_1 ? 2'h1 : _btb_362_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10154 = btb_362_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7018; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10156 = btb_362_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_362_bht_T_27 : _GEN_8554; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_363_bht_T = btb_363_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_363_bht_T_1 = io_i_branch_resolve_pack_taken & btb_363_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_363_bht_T_2 = btb_363_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_363_bht_T_3 = io_i_branch_resolve_pack_taken & btb_363_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_363_bht_T_4 = btb_363_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_363_bht_T_5 = io_i_branch_resolve_pack_taken & btb_363_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_363_bht_T_6 = btb_363_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_363_bht_T_7 = io_i_branch_resolve_pack_taken & btb_363_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_363_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_363_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_363_bht_T_13 = _btb_0_bht_T_8 & _btb_363_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_363_bht_T_16 = _btb_0_bht_T_8 & _btb_363_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_363_bht_T_19 = _btb_0_bht_T_8 & _btb_363_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_363_bht_T_20 = _btb_363_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_21 = _btb_363_bht_T_16 ? 2'h0 : _btb_363_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_22 = _btb_363_bht_T_13 ? 2'h0 : _btb_363_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_23 = _btb_363_bht_T_10 ? 2'h0 : _btb_363_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_24 = _btb_363_bht_T_7 ? 2'h3 : _btb_363_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_25 = _btb_363_bht_T_5 ? 2'h3 : _btb_363_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_26 = _btb_363_bht_T_3 ? 2'h3 : _btb_363_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_363_bht_T_27 = _btb_363_bht_T_1 ? 2'h1 : _btb_363_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10158 = btb_363_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7019; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10160 = btb_363_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_363_bht_T_27 : _GEN_8555; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_364_bht_T = btb_364_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_364_bht_T_1 = io_i_branch_resolve_pack_taken & btb_364_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_364_bht_T_2 = btb_364_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_364_bht_T_3 = io_i_branch_resolve_pack_taken & btb_364_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_364_bht_T_4 = btb_364_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_364_bht_T_5 = io_i_branch_resolve_pack_taken & btb_364_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_364_bht_T_6 = btb_364_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_364_bht_T_7 = io_i_branch_resolve_pack_taken & btb_364_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_364_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_364_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_364_bht_T_13 = _btb_0_bht_T_8 & _btb_364_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_364_bht_T_16 = _btb_0_bht_T_8 & _btb_364_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_364_bht_T_19 = _btb_0_bht_T_8 & _btb_364_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_364_bht_T_20 = _btb_364_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_21 = _btb_364_bht_T_16 ? 2'h0 : _btb_364_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_22 = _btb_364_bht_T_13 ? 2'h0 : _btb_364_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_23 = _btb_364_bht_T_10 ? 2'h0 : _btb_364_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_24 = _btb_364_bht_T_7 ? 2'h3 : _btb_364_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_25 = _btb_364_bht_T_5 ? 2'h3 : _btb_364_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_26 = _btb_364_bht_T_3 ? 2'h3 : _btb_364_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_364_bht_T_27 = _btb_364_bht_T_1 ? 2'h1 : _btb_364_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10162 = btb_364_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7020; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10164 = btb_364_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_364_bht_T_27 : _GEN_8556; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_365_bht_T = btb_365_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_365_bht_T_1 = io_i_branch_resolve_pack_taken & btb_365_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_365_bht_T_2 = btb_365_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_365_bht_T_3 = io_i_branch_resolve_pack_taken & btb_365_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_365_bht_T_4 = btb_365_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_365_bht_T_5 = io_i_branch_resolve_pack_taken & btb_365_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_365_bht_T_6 = btb_365_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_365_bht_T_7 = io_i_branch_resolve_pack_taken & btb_365_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_365_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_365_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_365_bht_T_13 = _btb_0_bht_T_8 & _btb_365_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_365_bht_T_16 = _btb_0_bht_T_8 & _btb_365_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_365_bht_T_19 = _btb_0_bht_T_8 & _btb_365_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_365_bht_T_20 = _btb_365_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_21 = _btb_365_bht_T_16 ? 2'h0 : _btb_365_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_22 = _btb_365_bht_T_13 ? 2'h0 : _btb_365_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_23 = _btb_365_bht_T_10 ? 2'h0 : _btb_365_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_24 = _btb_365_bht_T_7 ? 2'h3 : _btb_365_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_25 = _btb_365_bht_T_5 ? 2'h3 : _btb_365_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_26 = _btb_365_bht_T_3 ? 2'h3 : _btb_365_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_365_bht_T_27 = _btb_365_bht_T_1 ? 2'h1 : _btb_365_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10166 = btb_365_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7021; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10168 = btb_365_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_365_bht_T_27 : _GEN_8557; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_366_bht_T = btb_366_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_366_bht_T_1 = io_i_branch_resolve_pack_taken & btb_366_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_366_bht_T_2 = btb_366_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_366_bht_T_3 = io_i_branch_resolve_pack_taken & btb_366_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_366_bht_T_4 = btb_366_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_366_bht_T_5 = io_i_branch_resolve_pack_taken & btb_366_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_366_bht_T_6 = btb_366_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_366_bht_T_7 = io_i_branch_resolve_pack_taken & btb_366_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_366_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_366_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_366_bht_T_13 = _btb_0_bht_T_8 & _btb_366_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_366_bht_T_16 = _btb_0_bht_T_8 & _btb_366_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_366_bht_T_19 = _btb_0_bht_T_8 & _btb_366_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_366_bht_T_20 = _btb_366_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_21 = _btb_366_bht_T_16 ? 2'h0 : _btb_366_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_22 = _btb_366_bht_T_13 ? 2'h0 : _btb_366_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_23 = _btb_366_bht_T_10 ? 2'h0 : _btb_366_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_24 = _btb_366_bht_T_7 ? 2'h3 : _btb_366_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_25 = _btb_366_bht_T_5 ? 2'h3 : _btb_366_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_26 = _btb_366_bht_T_3 ? 2'h3 : _btb_366_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_366_bht_T_27 = _btb_366_bht_T_1 ? 2'h1 : _btb_366_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10170 = btb_366_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7022; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10172 = btb_366_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_366_bht_T_27 : _GEN_8558; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_367_bht_T = btb_367_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_367_bht_T_1 = io_i_branch_resolve_pack_taken & btb_367_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_367_bht_T_2 = btb_367_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_367_bht_T_3 = io_i_branch_resolve_pack_taken & btb_367_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_367_bht_T_4 = btb_367_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_367_bht_T_5 = io_i_branch_resolve_pack_taken & btb_367_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_367_bht_T_6 = btb_367_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_367_bht_T_7 = io_i_branch_resolve_pack_taken & btb_367_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_367_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_367_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_367_bht_T_13 = _btb_0_bht_T_8 & _btb_367_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_367_bht_T_16 = _btb_0_bht_T_8 & _btb_367_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_367_bht_T_19 = _btb_0_bht_T_8 & _btb_367_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_367_bht_T_20 = _btb_367_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_21 = _btb_367_bht_T_16 ? 2'h0 : _btb_367_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_22 = _btb_367_bht_T_13 ? 2'h0 : _btb_367_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_23 = _btb_367_bht_T_10 ? 2'h0 : _btb_367_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_24 = _btb_367_bht_T_7 ? 2'h3 : _btb_367_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_25 = _btb_367_bht_T_5 ? 2'h3 : _btb_367_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_26 = _btb_367_bht_T_3 ? 2'h3 : _btb_367_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_367_bht_T_27 = _btb_367_bht_T_1 ? 2'h1 : _btb_367_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10174 = btb_367_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7023; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10176 = btb_367_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_367_bht_T_27 : _GEN_8559; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_368_bht_T = btb_368_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_368_bht_T_1 = io_i_branch_resolve_pack_taken & btb_368_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_368_bht_T_2 = btb_368_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_368_bht_T_3 = io_i_branch_resolve_pack_taken & btb_368_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_368_bht_T_4 = btb_368_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_368_bht_T_5 = io_i_branch_resolve_pack_taken & btb_368_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_368_bht_T_6 = btb_368_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_368_bht_T_7 = io_i_branch_resolve_pack_taken & btb_368_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_368_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_368_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_368_bht_T_13 = _btb_0_bht_T_8 & _btb_368_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_368_bht_T_16 = _btb_0_bht_T_8 & _btb_368_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_368_bht_T_19 = _btb_0_bht_T_8 & _btb_368_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_368_bht_T_20 = _btb_368_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_21 = _btb_368_bht_T_16 ? 2'h0 : _btb_368_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_22 = _btb_368_bht_T_13 ? 2'h0 : _btb_368_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_23 = _btb_368_bht_T_10 ? 2'h0 : _btb_368_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_24 = _btb_368_bht_T_7 ? 2'h3 : _btb_368_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_25 = _btb_368_bht_T_5 ? 2'h3 : _btb_368_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_26 = _btb_368_bht_T_3 ? 2'h3 : _btb_368_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_368_bht_T_27 = _btb_368_bht_T_1 ? 2'h1 : _btb_368_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10178 = btb_368_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7024; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10180 = btb_368_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_368_bht_T_27 : _GEN_8560; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_369_bht_T = btb_369_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_369_bht_T_1 = io_i_branch_resolve_pack_taken & btb_369_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_369_bht_T_2 = btb_369_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_369_bht_T_3 = io_i_branch_resolve_pack_taken & btb_369_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_369_bht_T_4 = btb_369_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_369_bht_T_5 = io_i_branch_resolve_pack_taken & btb_369_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_369_bht_T_6 = btb_369_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_369_bht_T_7 = io_i_branch_resolve_pack_taken & btb_369_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_369_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_369_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_369_bht_T_13 = _btb_0_bht_T_8 & _btb_369_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_369_bht_T_16 = _btb_0_bht_T_8 & _btb_369_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_369_bht_T_19 = _btb_0_bht_T_8 & _btb_369_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_369_bht_T_20 = _btb_369_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_21 = _btb_369_bht_T_16 ? 2'h0 : _btb_369_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_22 = _btb_369_bht_T_13 ? 2'h0 : _btb_369_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_23 = _btb_369_bht_T_10 ? 2'h0 : _btb_369_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_24 = _btb_369_bht_T_7 ? 2'h3 : _btb_369_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_25 = _btb_369_bht_T_5 ? 2'h3 : _btb_369_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_26 = _btb_369_bht_T_3 ? 2'h3 : _btb_369_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_369_bht_T_27 = _btb_369_bht_T_1 ? 2'h1 : _btb_369_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10182 = btb_369_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7025; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10184 = btb_369_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_369_bht_T_27 : _GEN_8561; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_370_bht_T = btb_370_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_370_bht_T_1 = io_i_branch_resolve_pack_taken & btb_370_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_370_bht_T_2 = btb_370_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_370_bht_T_3 = io_i_branch_resolve_pack_taken & btb_370_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_370_bht_T_4 = btb_370_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_370_bht_T_5 = io_i_branch_resolve_pack_taken & btb_370_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_370_bht_T_6 = btb_370_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_370_bht_T_7 = io_i_branch_resolve_pack_taken & btb_370_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_370_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_370_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_370_bht_T_13 = _btb_0_bht_T_8 & _btb_370_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_370_bht_T_16 = _btb_0_bht_T_8 & _btb_370_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_370_bht_T_19 = _btb_0_bht_T_8 & _btb_370_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_370_bht_T_20 = _btb_370_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_21 = _btb_370_bht_T_16 ? 2'h0 : _btb_370_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_22 = _btb_370_bht_T_13 ? 2'h0 : _btb_370_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_23 = _btb_370_bht_T_10 ? 2'h0 : _btb_370_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_24 = _btb_370_bht_T_7 ? 2'h3 : _btb_370_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_25 = _btb_370_bht_T_5 ? 2'h3 : _btb_370_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_26 = _btb_370_bht_T_3 ? 2'h3 : _btb_370_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_370_bht_T_27 = _btb_370_bht_T_1 ? 2'h1 : _btb_370_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10186 = btb_370_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7026; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10188 = btb_370_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_370_bht_T_27 : _GEN_8562; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_371_bht_T = btb_371_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_371_bht_T_1 = io_i_branch_resolve_pack_taken & btb_371_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_371_bht_T_2 = btb_371_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_371_bht_T_3 = io_i_branch_resolve_pack_taken & btb_371_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_371_bht_T_4 = btb_371_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_371_bht_T_5 = io_i_branch_resolve_pack_taken & btb_371_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_371_bht_T_6 = btb_371_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_371_bht_T_7 = io_i_branch_resolve_pack_taken & btb_371_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_371_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_371_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_371_bht_T_13 = _btb_0_bht_T_8 & _btb_371_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_371_bht_T_16 = _btb_0_bht_T_8 & _btb_371_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_371_bht_T_19 = _btb_0_bht_T_8 & _btb_371_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_371_bht_T_20 = _btb_371_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_21 = _btb_371_bht_T_16 ? 2'h0 : _btb_371_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_22 = _btb_371_bht_T_13 ? 2'h0 : _btb_371_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_23 = _btb_371_bht_T_10 ? 2'h0 : _btb_371_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_24 = _btb_371_bht_T_7 ? 2'h3 : _btb_371_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_25 = _btb_371_bht_T_5 ? 2'h3 : _btb_371_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_26 = _btb_371_bht_T_3 ? 2'h3 : _btb_371_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_371_bht_T_27 = _btb_371_bht_T_1 ? 2'h1 : _btb_371_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10190 = btb_371_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7027; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10192 = btb_371_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_371_bht_T_27 : _GEN_8563; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_372_bht_T = btb_372_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_372_bht_T_1 = io_i_branch_resolve_pack_taken & btb_372_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_372_bht_T_2 = btb_372_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_372_bht_T_3 = io_i_branch_resolve_pack_taken & btb_372_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_372_bht_T_4 = btb_372_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_372_bht_T_5 = io_i_branch_resolve_pack_taken & btb_372_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_372_bht_T_6 = btb_372_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_372_bht_T_7 = io_i_branch_resolve_pack_taken & btb_372_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_372_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_372_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_372_bht_T_13 = _btb_0_bht_T_8 & _btb_372_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_372_bht_T_16 = _btb_0_bht_T_8 & _btb_372_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_372_bht_T_19 = _btb_0_bht_T_8 & _btb_372_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_372_bht_T_20 = _btb_372_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_21 = _btb_372_bht_T_16 ? 2'h0 : _btb_372_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_22 = _btb_372_bht_T_13 ? 2'h0 : _btb_372_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_23 = _btb_372_bht_T_10 ? 2'h0 : _btb_372_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_24 = _btb_372_bht_T_7 ? 2'h3 : _btb_372_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_25 = _btb_372_bht_T_5 ? 2'h3 : _btb_372_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_26 = _btb_372_bht_T_3 ? 2'h3 : _btb_372_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_372_bht_T_27 = _btb_372_bht_T_1 ? 2'h1 : _btb_372_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10194 = btb_372_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7028; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10196 = btb_372_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_372_bht_T_27 : _GEN_8564; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_373_bht_T = btb_373_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_373_bht_T_1 = io_i_branch_resolve_pack_taken & btb_373_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_373_bht_T_2 = btb_373_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_373_bht_T_3 = io_i_branch_resolve_pack_taken & btb_373_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_373_bht_T_4 = btb_373_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_373_bht_T_5 = io_i_branch_resolve_pack_taken & btb_373_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_373_bht_T_6 = btb_373_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_373_bht_T_7 = io_i_branch_resolve_pack_taken & btb_373_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_373_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_373_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_373_bht_T_13 = _btb_0_bht_T_8 & _btb_373_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_373_bht_T_16 = _btb_0_bht_T_8 & _btb_373_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_373_bht_T_19 = _btb_0_bht_T_8 & _btb_373_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_373_bht_T_20 = _btb_373_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_21 = _btb_373_bht_T_16 ? 2'h0 : _btb_373_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_22 = _btb_373_bht_T_13 ? 2'h0 : _btb_373_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_23 = _btb_373_bht_T_10 ? 2'h0 : _btb_373_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_24 = _btb_373_bht_T_7 ? 2'h3 : _btb_373_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_25 = _btb_373_bht_T_5 ? 2'h3 : _btb_373_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_26 = _btb_373_bht_T_3 ? 2'h3 : _btb_373_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_373_bht_T_27 = _btb_373_bht_T_1 ? 2'h1 : _btb_373_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10198 = btb_373_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7029; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10200 = btb_373_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_373_bht_T_27 : _GEN_8565; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_374_bht_T = btb_374_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_374_bht_T_1 = io_i_branch_resolve_pack_taken & btb_374_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_374_bht_T_2 = btb_374_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_374_bht_T_3 = io_i_branch_resolve_pack_taken & btb_374_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_374_bht_T_4 = btb_374_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_374_bht_T_5 = io_i_branch_resolve_pack_taken & btb_374_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_374_bht_T_6 = btb_374_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_374_bht_T_7 = io_i_branch_resolve_pack_taken & btb_374_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_374_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_374_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_374_bht_T_13 = _btb_0_bht_T_8 & _btb_374_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_374_bht_T_16 = _btb_0_bht_T_8 & _btb_374_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_374_bht_T_19 = _btb_0_bht_T_8 & _btb_374_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_374_bht_T_20 = _btb_374_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_21 = _btb_374_bht_T_16 ? 2'h0 : _btb_374_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_22 = _btb_374_bht_T_13 ? 2'h0 : _btb_374_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_23 = _btb_374_bht_T_10 ? 2'h0 : _btb_374_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_24 = _btb_374_bht_T_7 ? 2'h3 : _btb_374_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_25 = _btb_374_bht_T_5 ? 2'h3 : _btb_374_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_26 = _btb_374_bht_T_3 ? 2'h3 : _btb_374_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_374_bht_T_27 = _btb_374_bht_T_1 ? 2'h1 : _btb_374_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10201 = btb_374_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_373_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_372_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_371_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_370_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_369_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_368_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_367_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_366_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_365_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_364_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_363_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_362_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_361_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_360_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10141)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10202 = btb_374_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7030; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10204 = btb_374_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_374_bht_T_27 : _GEN_8566; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_375_bht_T = btb_375_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_375_bht_T_1 = io_i_branch_resolve_pack_taken & btb_375_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_375_bht_T_2 = btb_375_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_375_bht_T_3 = io_i_branch_resolve_pack_taken & btb_375_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_375_bht_T_4 = btb_375_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_375_bht_T_5 = io_i_branch_resolve_pack_taken & btb_375_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_375_bht_T_6 = btb_375_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_375_bht_T_7 = io_i_branch_resolve_pack_taken & btb_375_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_375_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_375_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_375_bht_T_13 = _btb_0_bht_T_8 & _btb_375_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_375_bht_T_16 = _btb_0_bht_T_8 & _btb_375_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_375_bht_T_19 = _btb_0_bht_T_8 & _btb_375_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_375_bht_T_20 = _btb_375_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_21 = _btb_375_bht_T_16 ? 2'h0 : _btb_375_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_22 = _btb_375_bht_T_13 ? 2'h0 : _btb_375_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_23 = _btb_375_bht_T_10 ? 2'h0 : _btb_375_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_24 = _btb_375_bht_T_7 ? 2'h3 : _btb_375_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_25 = _btb_375_bht_T_5 ? 2'h3 : _btb_375_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_26 = _btb_375_bht_T_3 ? 2'h3 : _btb_375_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_375_bht_T_27 = _btb_375_bht_T_1 ? 2'h1 : _btb_375_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10206 = btb_375_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7031; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10208 = btb_375_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_375_bht_T_27 : _GEN_8567; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_376_bht_T = btb_376_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_376_bht_T_1 = io_i_branch_resolve_pack_taken & btb_376_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_376_bht_T_2 = btb_376_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_376_bht_T_3 = io_i_branch_resolve_pack_taken & btb_376_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_376_bht_T_4 = btb_376_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_376_bht_T_5 = io_i_branch_resolve_pack_taken & btb_376_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_376_bht_T_6 = btb_376_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_376_bht_T_7 = io_i_branch_resolve_pack_taken & btb_376_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_376_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_376_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_376_bht_T_13 = _btb_0_bht_T_8 & _btb_376_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_376_bht_T_16 = _btb_0_bht_T_8 & _btb_376_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_376_bht_T_19 = _btb_0_bht_T_8 & _btb_376_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_376_bht_T_20 = _btb_376_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_21 = _btb_376_bht_T_16 ? 2'h0 : _btb_376_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_22 = _btb_376_bht_T_13 ? 2'h0 : _btb_376_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_23 = _btb_376_bht_T_10 ? 2'h0 : _btb_376_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_24 = _btb_376_bht_T_7 ? 2'h3 : _btb_376_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_25 = _btb_376_bht_T_5 ? 2'h3 : _btb_376_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_26 = _btb_376_bht_T_3 ? 2'h3 : _btb_376_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_376_bht_T_27 = _btb_376_bht_T_1 ? 2'h1 : _btb_376_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10210 = btb_376_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7032; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10212 = btb_376_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_376_bht_T_27 : _GEN_8568; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_377_bht_T = btb_377_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_377_bht_T_1 = io_i_branch_resolve_pack_taken & btb_377_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_377_bht_T_2 = btb_377_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_377_bht_T_3 = io_i_branch_resolve_pack_taken & btb_377_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_377_bht_T_4 = btb_377_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_377_bht_T_5 = io_i_branch_resolve_pack_taken & btb_377_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_377_bht_T_6 = btb_377_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_377_bht_T_7 = io_i_branch_resolve_pack_taken & btb_377_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_377_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_377_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_377_bht_T_13 = _btb_0_bht_T_8 & _btb_377_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_377_bht_T_16 = _btb_0_bht_T_8 & _btb_377_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_377_bht_T_19 = _btb_0_bht_T_8 & _btb_377_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_377_bht_T_20 = _btb_377_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_21 = _btb_377_bht_T_16 ? 2'h0 : _btb_377_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_22 = _btb_377_bht_T_13 ? 2'h0 : _btb_377_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_23 = _btb_377_bht_T_10 ? 2'h0 : _btb_377_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_24 = _btb_377_bht_T_7 ? 2'h3 : _btb_377_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_25 = _btb_377_bht_T_5 ? 2'h3 : _btb_377_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_26 = _btb_377_bht_T_3 ? 2'h3 : _btb_377_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_377_bht_T_27 = _btb_377_bht_T_1 ? 2'h1 : _btb_377_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10214 = btb_377_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7033; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10216 = btb_377_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_377_bht_T_27 : _GEN_8569; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_378_bht_T = btb_378_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_378_bht_T_1 = io_i_branch_resolve_pack_taken & btb_378_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_378_bht_T_2 = btb_378_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_378_bht_T_3 = io_i_branch_resolve_pack_taken & btb_378_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_378_bht_T_4 = btb_378_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_378_bht_T_5 = io_i_branch_resolve_pack_taken & btb_378_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_378_bht_T_6 = btb_378_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_378_bht_T_7 = io_i_branch_resolve_pack_taken & btb_378_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_378_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_378_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_378_bht_T_13 = _btb_0_bht_T_8 & _btb_378_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_378_bht_T_16 = _btb_0_bht_T_8 & _btb_378_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_378_bht_T_19 = _btb_0_bht_T_8 & _btb_378_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_378_bht_T_20 = _btb_378_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_21 = _btb_378_bht_T_16 ? 2'h0 : _btb_378_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_22 = _btb_378_bht_T_13 ? 2'h0 : _btb_378_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_23 = _btb_378_bht_T_10 ? 2'h0 : _btb_378_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_24 = _btb_378_bht_T_7 ? 2'h3 : _btb_378_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_25 = _btb_378_bht_T_5 ? 2'h3 : _btb_378_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_26 = _btb_378_bht_T_3 ? 2'h3 : _btb_378_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_378_bht_T_27 = _btb_378_bht_T_1 ? 2'h1 : _btb_378_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10218 = btb_378_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7034; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10220 = btb_378_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_378_bht_T_27 : _GEN_8570; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_379_bht_T = btb_379_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_379_bht_T_1 = io_i_branch_resolve_pack_taken & btb_379_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_379_bht_T_2 = btb_379_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_379_bht_T_3 = io_i_branch_resolve_pack_taken & btb_379_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_379_bht_T_4 = btb_379_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_379_bht_T_5 = io_i_branch_resolve_pack_taken & btb_379_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_379_bht_T_6 = btb_379_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_379_bht_T_7 = io_i_branch_resolve_pack_taken & btb_379_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_379_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_379_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_379_bht_T_13 = _btb_0_bht_T_8 & _btb_379_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_379_bht_T_16 = _btb_0_bht_T_8 & _btb_379_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_379_bht_T_19 = _btb_0_bht_T_8 & _btb_379_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_379_bht_T_20 = _btb_379_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_21 = _btb_379_bht_T_16 ? 2'h0 : _btb_379_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_22 = _btb_379_bht_T_13 ? 2'h0 : _btb_379_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_23 = _btb_379_bht_T_10 ? 2'h0 : _btb_379_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_24 = _btb_379_bht_T_7 ? 2'h3 : _btb_379_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_25 = _btb_379_bht_T_5 ? 2'h3 : _btb_379_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_26 = _btb_379_bht_T_3 ? 2'h3 : _btb_379_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_379_bht_T_27 = _btb_379_bht_T_1 ? 2'h1 : _btb_379_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10222 = btb_379_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7035; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10224 = btb_379_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_379_bht_T_27 : _GEN_8571; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_380_bht_T = btb_380_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_380_bht_T_1 = io_i_branch_resolve_pack_taken & btb_380_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_380_bht_T_2 = btb_380_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_380_bht_T_3 = io_i_branch_resolve_pack_taken & btb_380_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_380_bht_T_4 = btb_380_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_380_bht_T_5 = io_i_branch_resolve_pack_taken & btb_380_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_380_bht_T_6 = btb_380_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_380_bht_T_7 = io_i_branch_resolve_pack_taken & btb_380_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_380_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_380_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_380_bht_T_13 = _btb_0_bht_T_8 & _btb_380_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_380_bht_T_16 = _btb_0_bht_T_8 & _btb_380_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_380_bht_T_19 = _btb_0_bht_T_8 & _btb_380_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_380_bht_T_20 = _btb_380_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_21 = _btb_380_bht_T_16 ? 2'h0 : _btb_380_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_22 = _btb_380_bht_T_13 ? 2'h0 : _btb_380_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_23 = _btb_380_bht_T_10 ? 2'h0 : _btb_380_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_24 = _btb_380_bht_T_7 ? 2'h3 : _btb_380_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_25 = _btb_380_bht_T_5 ? 2'h3 : _btb_380_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_26 = _btb_380_bht_T_3 ? 2'h3 : _btb_380_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_380_bht_T_27 = _btb_380_bht_T_1 ? 2'h1 : _btb_380_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10226 = btb_380_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7036; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10228 = btb_380_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_380_bht_T_27 : _GEN_8572; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_381_bht_T = btb_381_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_381_bht_T_1 = io_i_branch_resolve_pack_taken & btb_381_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_381_bht_T_2 = btb_381_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_381_bht_T_3 = io_i_branch_resolve_pack_taken & btb_381_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_381_bht_T_4 = btb_381_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_381_bht_T_5 = io_i_branch_resolve_pack_taken & btb_381_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_381_bht_T_6 = btb_381_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_381_bht_T_7 = io_i_branch_resolve_pack_taken & btb_381_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_381_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_381_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_381_bht_T_13 = _btb_0_bht_T_8 & _btb_381_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_381_bht_T_16 = _btb_0_bht_T_8 & _btb_381_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_381_bht_T_19 = _btb_0_bht_T_8 & _btb_381_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_381_bht_T_20 = _btb_381_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_21 = _btb_381_bht_T_16 ? 2'h0 : _btb_381_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_22 = _btb_381_bht_T_13 ? 2'h0 : _btb_381_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_23 = _btb_381_bht_T_10 ? 2'h0 : _btb_381_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_24 = _btb_381_bht_T_7 ? 2'h3 : _btb_381_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_25 = _btb_381_bht_T_5 ? 2'h3 : _btb_381_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_26 = _btb_381_bht_T_3 ? 2'h3 : _btb_381_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_381_bht_T_27 = _btb_381_bht_T_1 ? 2'h1 : _btb_381_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10230 = btb_381_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7037; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10232 = btb_381_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_381_bht_T_27 : _GEN_8573; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_382_bht_T = btb_382_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_382_bht_T_1 = io_i_branch_resolve_pack_taken & btb_382_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_382_bht_T_2 = btb_382_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_382_bht_T_3 = io_i_branch_resolve_pack_taken & btb_382_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_382_bht_T_4 = btb_382_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_382_bht_T_5 = io_i_branch_resolve_pack_taken & btb_382_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_382_bht_T_6 = btb_382_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_382_bht_T_7 = io_i_branch_resolve_pack_taken & btb_382_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_382_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_382_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_382_bht_T_13 = _btb_0_bht_T_8 & _btb_382_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_382_bht_T_16 = _btb_0_bht_T_8 & _btb_382_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_382_bht_T_19 = _btb_0_bht_T_8 & _btb_382_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_382_bht_T_20 = _btb_382_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_21 = _btb_382_bht_T_16 ? 2'h0 : _btb_382_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_22 = _btb_382_bht_T_13 ? 2'h0 : _btb_382_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_23 = _btb_382_bht_T_10 ? 2'h0 : _btb_382_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_24 = _btb_382_bht_T_7 ? 2'h3 : _btb_382_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_25 = _btb_382_bht_T_5 ? 2'h3 : _btb_382_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_26 = _btb_382_bht_T_3 ? 2'h3 : _btb_382_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_382_bht_T_27 = _btb_382_bht_T_1 ? 2'h1 : _btb_382_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10234 = btb_382_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7038; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10236 = btb_382_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_382_bht_T_27 : _GEN_8574; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_383_bht_T = btb_383_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_383_bht_T_1 = io_i_branch_resolve_pack_taken & btb_383_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_383_bht_T_2 = btb_383_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_383_bht_T_3 = io_i_branch_resolve_pack_taken & btb_383_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_383_bht_T_4 = btb_383_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_383_bht_T_5 = io_i_branch_resolve_pack_taken & btb_383_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_383_bht_T_6 = btb_383_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_383_bht_T_7 = io_i_branch_resolve_pack_taken & btb_383_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_383_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_383_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_383_bht_T_13 = _btb_0_bht_T_8 & _btb_383_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_383_bht_T_16 = _btb_0_bht_T_8 & _btb_383_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_383_bht_T_19 = _btb_0_bht_T_8 & _btb_383_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_383_bht_T_20 = _btb_383_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_21 = _btb_383_bht_T_16 ? 2'h0 : _btb_383_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_22 = _btb_383_bht_T_13 ? 2'h0 : _btb_383_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_23 = _btb_383_bht_T_10 ? 2'h0 : _btb_383_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_24 = _btb_383_bht_T_7 ? 2'h3 : _btb_383_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_25 = _btb_383_bht_T_5 ? 2'h3 : _btb_383_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_26 = _btb_383_bht_T_3 ? 2'h3 : _btb_383_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_383_bht_T_27 = _btb_383_bht_T_1 ? 2'h1 : _btb_383_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10238 = btb_383_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7039; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10240 = btb_383_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_383_bht_T_27 : _GEN_8575; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_384_bht_T = btb_384_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_384_bht_T_1 = io_i_branch_resolve_pack_taken & btb_384_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_384_bht_T_2 = btb_384_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_384_bht_T_3 = io_i_branch_resolve_pack_taken & btb_384_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_384_bht_T_4 = btb_384_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_384_bht_T_5 = io_i_branch_resolve_pack_taken & btb_384_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_384_bht_T_6 = btb_384_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_384_bht_T_7 = io_i_branch_resolve_pack_taken & btb_384_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_384_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_384_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_384_bht_T_13 = _btb_0_bht_T_8 & _btb_384_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_384_bht_T_16 = _btb_0_bht_T_8 & _btb_384_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_384_bht_T_19 = _btb_0_bht_T_8 & _btb_384_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_384_bht_T_20 = _btb_384_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_21 = _btb_384_bht_T_16 ? 2'h0 : _btb_384_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_22 = _btb_384_bht_T_13 ? 2'h0 : _btb_384_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_23 = _btb_384_bht_T_10 ? 2'h0 : _btb_384_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_24 = _btb_384_bht_T_7 ? 2'h3 : _btb_384_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_25 = _btb_384_bht_T_5 ? 2'h3 : _btb_384_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_26 = _btb_384_bht_T_3 ? 2'h3 : _btb_384_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_384_bht_T_27 = _btb_384_bht_T_1 ? 2'h1 : _btb_384_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10242 = btb_384_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7040; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10244 = btb_384_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_384_bht_T_27 : _GEN_8576; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_385_bht_T = btb_385_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_385_bht_T_1 = io_i_branch_resolve_pack_taken & btb_385_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_385_bht_T_2 = btb_385_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_385_bht_T_3 = io_i_branch_resolve_pack_taken & btb_385_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_385_bht_T_4 = btb_385_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_385_bht_T_5 = io_i_branch_resolve_pack_taken & btb_385_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_385_bht_T_6 = btb_385_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_385_bht_T_7 = io_i_branch_resolve_pack_taken & btb_385_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_385_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_385_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_385_bht_T_13 = _btb_0_bht_T_8 & _btb_385_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_385_bht_T_16 = _btb_0_bht_T_8 & _btb_385_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_385_bht_T_19 = _btb_0_bht_T_8 & _btb_385_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_385_bht_T_20 = _btb_385_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_21 = _btb_385_bht_T_16 ? 2'h0 : _btb_385_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_22 = _btb_385_bht_T_13 ? 2'h0 : _btb_385_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_23 = _btb_385_bht_T_10 ? 2'h0 : _btb_385_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_24 = _btb_385_bht_T_7 ? 2'h3 : _btb_385_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_25 = _btb_385_bht_T_5 ? 2'h3 : _btb_385_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_26 = _btb_385_bht_T_3 ? 2'h3 : _btb_385_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_385_bht_T_27 = _btb_385_bht_T_1 ? 2'h1 : _btb_385_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10246 = btb_385_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7041; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10248 = btb_385_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_385_bht_T_27 : _GEN_8577; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_386_bht_T = btb_386_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_386_bht_T_1 = io_i_branch_resolve_pack_taken & btb_386_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_386_bht_T_2 = btb_386_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_386_bht_T_3 = io_i_branch_resolve_pack_taken & btb_386_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_386_bht_T_4 = btb_386_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_386_bht_T_5 = io_i_branch_resolve_pack_taken & btb_386_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_386_bht_T_6 = btb_386_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_386_bht_T_7 = io_i_branch_resolve_pack_taken & btb_386_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_386_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_386_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_386_bht_T_13 = _btb_0_bht_T_8 & _btb_386_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_386_bht_T_16 = _btb_0_bht_T_8 & _btb_386_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_386_bht_T_19 = _btb_0_bht_T_8 & _btb_386_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_386_bht_T_20 = _btb_386_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_21 = _btb_386_bht_T_16 ? 2'h0 : _btb_386_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_22 = _btb_386_bht_T_13 ? 2'h0 : _btb_386_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_23 = _btb_386_bht_T_10 ? 2'h0 : _btb_386_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_24 = _btb_386_bht_T_7 ? 2'h3 : _btb_386_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_25 = _btb_386_bht_T_5 ? 2'h3 : _btb_386_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_26 = _btb_386_bht_T_3 ? 2'h3 : _btb_386_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_386_bht_T_27 = _btb_386_bht_T_1 ? 2'h1 : _btb_386_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10250 = btb_386_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7042; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10252 = btb_386_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_386_bht_T_27 : _GEN_8578; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_387_bht_T = btb_387_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_387_bht_T_1 = io_i_branch_resolve_pack_taken & btb_387_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_387_bht_T_2 = btb_387_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_387_bht_T_3 = io_i_branch_resolve_pack_taken & btb_387_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_387_bht_T_4 = btb_387_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_387_bht_T_5 = io_i_branch_resolve_pack_taken & btb_387_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_387_bht_T_6 = btb_387_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_387_bht_T_7 = io_i_branch_resolve_pack_taken & btb_387_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_387_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_387_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_387_bht_T_13 = _btb_0_bht_T_8 & _btb_387_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_387_bht_T_16 = _btb_0_bht_T_8 & _btb_387_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_387_bht_T_19 = _btb_0_bht_T_8 & _btb_387_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_387_bht_T_20 = _btb_387_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_21 = _btb_387_bht_T_16 ? 2'h0 : _btb_387_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_22 = _btb_387_bht_T_13 ? 2'h0 : _btb_387_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_23 = _btb_387_bht_T_10 ? 2'h0 : _btb_387_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_24 = _btb_387_bht_T_7 ? 2'h3 : _btb_387_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_25 = _btb_387_bht_T_5 ? 2'h3 : _btb_387_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_26 = _btb_387_bht_T_3 ? 2'h3 : _btb_387_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_387_bht_T_27 = _btb_387_bht_T_1 ? 2'h1 : _btb_387_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10254 = btb_387_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7043; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10256 = btb_387_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_387_bht_T_27 : _GEN_8579; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_388_bht_T = btb_388_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_388_bht_T_1 = io_i_branch_resolve_pack_taken & btb_388_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_388_bht_T_2 = btb_388_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_388_bht_T_3 = io_i_branch_resolve_pack_taken & btb_388_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_388_bht_T_4 = btb_388_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_388_bht_T_5 = io_i_branch_resolve_pack_taken & btb_388_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_388_bht_T_6 = btb_388_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_388_bht_T_7 = io_i_branch_resolve_pack_taken & btb_388_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_388_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_388_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_388_bht_T_13 = _btb_0_bht_T_8 & _btb_388_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_388_bht_T_16 = _btb_0_bht_T_8 & _btb_388_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_388_bht_T_19 = _btb_0_bht_T_8 & _btb_388_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_388_bht_T_20 = _btb_388_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_21 = _btb_388_bht_T_16 ? 2'h0 : _btb_388_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_22 = _btb_388_bht_T_13 ? 2'h0 : _btb_388_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_23 = _btb_388_bht_T_10 ? 2'h0 : _btb_388_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_24 = _btb_388_bht_T_7 ? 2'h3 : _btb_388_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_25 = _btb_388_bht_T_5 ? 2'h3 : _btb_388_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_26 = _btb_388_bht_T_3 ? 2'h3 : _btb_388_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_388_bht_T_27 = _btb_388_bht_T_1 ? 2'h1 : _btb_388_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10258 = btb_388_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7044; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10260 = btb_388_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_388_bht_T_27 : _GEN_8580; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_389_bht_T = btb_389_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_389_bht_T_1 = io_i_branch_resolve_pack_taken & btb_389_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_389_bht_T_2 = btb_389_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_389_bht_T_3 = io_i_branch_resolve_pack_taken & btb_389_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_389_bht_T_4 = btb_389_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_389_bht_T_5 = io_i_branch_resolve_pack_taken & btb_389_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_389_bht_T_6 = btb_389_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_389_bht_T_7 = io_i_branch_resolve_pack_taken & btb_389_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_389_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_389_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_389_bht_T_13 = _btb_0_bht_T_8 & _btb_389_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_389_bht_T_16 = _btb_0_bht_T_8 & _btb_389_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_389_bht_T_19 = _btb_0_bht_T_8 & _btb_389_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_389_bht_T_20 = _btb_389_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_21 = _btb_389_bht_T_16 ? 2'h0 : _btb_389_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_22 = _btb_389_bht_T_13 ? 2'h0 : _btb_389_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_23 = _btb_389_bht_T_10 ? 2'h0 : _btb_389_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_24 = _btb_389_bht_T_7 ? 2'h3 : _btb_389_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_25 = _btb_389_bht_T_5 ? 2'h3 : _btb_389_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_26 = _btb_389_bht_T_3 ? 2'h3 : _btb_389_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_389_bht_T_27 = _btb_389_bht_T_1 ? 2'h1 : _btb_389_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10261 = btb_389_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_388_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_387_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_386_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_385_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_384_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_383_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_382_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_381_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_380_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_379_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_378_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_377_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_376_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_375_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10201)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10262 = btb_389_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7045; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10264 = btb_389_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_389_bht_T_27 : _GEN_8581; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_390_bht_T = btb_390_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_390_bht_T_1 = io_i_branch_resolve_pack_taken & btb_390_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_390_bht_T_2 = btb_390_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_390_bht_T_3 = io_i_branch_resolve_pack_taken & btb_390_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_390_bht_T_4 = btb_390_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_390_bht_T_5 = io_i_branch_resolve_pack_taken & btb_390_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_390_bht_T_6 = btb_390_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_390_bht_T_7 = io_i_branch_resolve_pack_taken & btb_390_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_390_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_390_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_390_bht_T_13 = _btb_0_bht_T_8 & _btb_390_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_390_bht_T_16 = _btb_0_bht_T_8 & _btb_390_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_390_bht_T_19 = _btb_0_bht_T_8 & _btb_390_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_390_bht_T_20 = _btb_390_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_21 = _btb_390_bht_T_16 ? 2'h0 : _btb_390_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_22 = _btb_390_bht_T_13 ? 2'h0 : _btb_390_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_23 = _btb_390_bht_T_10 ? 2'h0 : _btb_390_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_24 = _btb_390_bht_T_7 ? 2'h3 : _btb_390_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_25 = _btb_390_bht_T_5 ? 2'h3 : _btb_390_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_26 = _btb_390_bht_T_3 ? 2'h3 : _btb_390_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_390_bht_T_27 = _btb_390_bht_T_1 ? 2'h1 : _btb_390_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10266 = btb_390_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7046; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10268 = btb_390_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_390_bht_T_27 : _GEN_8582; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_391_bht_T = btb_391_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_391_bht_T_1 = io_i_branch_resolve_pack_taken & btb_391_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_391_bht_T_2 = btb_391_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_391_bht_T_3 = io_i_branch_resolve_pack_taken & btb_391_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_391_bht_T_4 = btb_391_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_391_bht_T_5 = io_i_branch_resolve_pack_taken & btb_391_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_391_bht_T_6 = btb_391_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_391_bht_T_7 = io_i_branch_resolve_pack_taken & btb_391_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_391_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_391_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_391_bht_T_13 = _btb_0_bht_T_8 & _btb_391_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_391_bht_T_16 = _btb_0_bht_T_8 & _btb_391_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_391_bht_T_19 = _btb_0_bht_T_8 & _btb_391_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_391_bht_T_20 = _btb_391_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_21 = _btb_391_bht_T_16 ? 2'h0 : _btb_391_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_22 = _btb_391_bht_T_13 ? 2'h0 : _btb_391_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_23 = _btb_391_bht_T_10 ? 2'h0 : _btb_391_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_24 = _btb_391_bht_T_7 ? 2'h3 : _btb_391_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_25 = _btb_391_bht_T_5 ? 2'h3 : _btb_391_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_26 = _btb_391_bht_T_3 ? 2'h3 : _btb_391_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_391_bht_T_27 = _btb_391_bht_T_1 ? 2'h1 : _btb_391_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10270 = btb_391_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7047; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10272 = btb_391_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_391_bht_T_27 : _GEN_8583; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_392_bht_T = btb_392_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_392_bht_T_1 = io_i_branch_resolve_pack_taken & btb_392_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_392_bht_T_2 = btb_392_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_392_bht_T_3 = io_i_branch_resolve_pack_taken & btb_392_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_392_bht_T_4 = btb_392_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_392_bht_T_5 = io_i_branch_resolve_pack_taken & btb_392_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_392_bht_T_6 = btb_392_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_392_bht_T_7 = io_i_branch_resolve_pack_taken & btb_392_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_392_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_392_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_392_bht_T_13 = _btb_0_bht_T_8 & _btb_392_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_392_bht_T_16 = _btb_0_bht_T_8 & _btb_392_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_392_bht_T_19 = _btb_0_bht_T_8 & _btb_392_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_392_bht_T_20 = _btb_392_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_21 = _btb_392_bht_T_16 ? 2'h0 : _btb_392_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_22 = _btb_392_bht_T_13 ? 2'h0 : _btb_392_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_23 = _btb_392_bht_T_10 ? 2'h0 : _btb_392_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_24 = _btb_392_bht_T_7 ? 2'h3 : _btb_392_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_25 = _btb_392_bht_T_5 ? 2'h3 : _btb_392_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_26 = _btb_392_bht_T_3 ? 2'h3 : _btb_392_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_392_bht_T_27 = _btb_392_bht_T_1 ? 2'h1 : _btb_392_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10274 = btb_392_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7048; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10276 = btb_392_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_392_bht_T_27 : _GEN_8584; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_393_bht_T = btb_393_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_393_bht_T_1 = io_i_branch_resolve_pack_taken & btb_393_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_393_bht_T_2 = btb_393_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_393_bht_T_3 = io_i_branch_resolve_pack_taken & btb_393_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_393_bht_T_4 = btb_393_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_393_bht_T_5 = io_i_branch_resolve_pack_taken & btb_393_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_393_bht_T_6 = btb_393_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_393_bht_T_7 = io_i_branch_resolve_pack_taken & btb_393_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_393_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_393_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_393_bht_T_13 = _btb_0_bht_T_8 & _btb_393_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_393_bht_T_16 = _btb_0_bht_T_8 & _btb_393_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_393_bht_T_19 = _btb_0_bht_T_8 & _btb_393_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_393_bht_T_20 = _btb_393_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_21 = _btb_393_bht_T_16 ? 2'h0 : _btb_393_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_22 = _btb_393_bht_T_13 ? 2'h0 : _btb_393_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_23 = _btb_393_bht_T_10 ? 2'h0 : _btb_393_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_24 = _btb_393_bht_T_7 ? 2'h3 : _btb_393_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_25 = _btb_393_bht_T_5 ? 2'h3 : _btb_393_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_26 = _btb_393_bht_T_3 ? 2'h3 : _btb_393_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_393_bht_T_27 = _btb_393_bht_T_1 ? 2'h1 : _btb_393_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10278 = btb_393_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7049; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10280 = btb_393_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_393_bht_T_27 : _GEN_8585; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_394_bht_T = btb_394_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_394_bht_T_1 = io_i_branch_resolve_pack_taken & btb_394_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_394_bht_T_2 = btb_394_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_394_bht_T_3 = io_i_branch_resolve_pack_taken & btb_394_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_394_bht_T_4 = btb_394_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_394_bht_T_5 = io_i_branch_resolve_pack_taken & btb_394_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_394_bht_T_6 = btb_394_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_394_bht_T_7 = io_i_branch_resolve_pack_taken & btb_394_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_394_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_394_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_394_bht_T_13 = _btb_0_bht_T_8 & _btb_394_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_394_bht_T_16 = _btb_0_bht_T_8 & _btb_394_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_394_bht_T_19 = _btb_0_bht_T_8 & _btb_394_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_394_bht_T_20 = _btb_394_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_21 = _btb_394_bht_T_16 ? 2'h0 : _btb_394_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_22 = _btb_394_bht_T_13 ? 2'h0 : _btb_394_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_23 = _btb_394_bht_T_10 ? 2'h0 : _btb_394_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_24 = _btb_394_bht_T_7 ? 2'h3 : _btb_394_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_25 = _btb_394_bht_T_5 ? 2'h3 : _btb_394_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_26 = _btb_394_bht_T_3 ? 2'h3 : _btb_394_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_394_bht_T_27 = _btb_394_bht_T_1 ? 2'h1 : _btb_394_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10282 = btb_394_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7050; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10284 = btb_394_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_394_bht_T_27 : _GEN_8586; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_395_bht_T = btb_395_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_395_bht_T_1 = io_i_branch_resolve_pack_taken & btb_395_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_395_bht_T_2 = btb_395_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_395_bht_T_3 = io_i_branch_resolve_pack_taken & btb_395_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_395_bht_T_4 = btb_395_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_395_bht_T_5 = io_i_branch_resolve_pack_taken & btb_395_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_395_bht_T_6 = btb_395_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_395_bht_T_7 = io_i_branch_resolve_pack_taken & btb_395_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_395_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_395_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_395_bht_T_13 = _btb_0_bht_T_8 & _btb_395_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_395_bht_T_16 = _btb_0_bht_T_8 & _btb_395_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_395_bht_T_19 = _btb_0_bht_T_8 & _btb_395_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_395_bht_T_20 = _btb_395_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_21 = _btb_395_bht_T_16 ? 2'h0 : _btb_395_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_22 = _btb_395_bht_T_13 ? 2'h0 : _btb_395_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_23 = _btb_395_bht_T_10 ? 2'h0 : _btb_395_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_24 = _btb_395_bht_T_7 ? 2'h3 : _btb_395_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_25 = _btb_395_bht_T_5 ? 2'h3 : _btb_395_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_26 = _btb_395_bht_T_3 ? 2'h3 : _btb_395_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_395_bht_T_27 = _btb_395_bht_T_1 ? 2'h1 : _btb_395_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10286 = btb_395_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7051; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10288 = btb_395_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_395_bht_T_27 : _GEN_8587; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_396_bht_T = btb_396_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_396_bht_T_1 = io_i_branch_resolve_pack_taken & btb_396_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_396_bht_T_2 = btb_396_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_396_bht_T_3 = io_i_branch_resolve_pack_taken & btb_396_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_396_bht_T_4 = btb_396_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_396_bht_T_5 = io_i_branch_resolve_pack_taken & btb_396_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_396_bht_T_6 = btb_396_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_396_bht_T_7 = io_i_branch_resolve_pack_taken & btb_396_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_396_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_396_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_396_bht_T_13 = _btb_0_bht_T_8 & _btb_396_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_396_bht_T_16 = _btb_0_bht_T_8 & _btb_396_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_396_bht_T_19 = _btb_0_bht_T_8 & _btb_396_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_396_bht_T_20 = _btb_396_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_21 = _btb_396_bht_T_16 ? 2'h0 : _btb_396_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_22 = _btb_396_bht_T_13 ? 2'h0 : _btb_396_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_23 = _btb_396_bht_T_10 ? 2'h0 : _btb_396_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_24 = _btb_396_bht_T_7 ? 2'h3 : _btb_396_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_25 = _btb_396_bht_T_5 ? 2'h3 : _btb_396_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_26 = _btb_396_bht_T_3 ? 2'h3 : _btb_396_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_396_bht_T_27 = _btb_396_bht_T_1 ? 2'h1 : _btb_396_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10290 = btb_396_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7052; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10292 = btb_396_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_396_bht_T_27 : _GEN_8588; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_397_bht_T = btb_397_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_397_bht_T_1 = io_i_branch_resolve_pack_taken & btb_397_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_397_bht_T_2 = btb_397_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_397_bht_T_3 = io_i_branch_resolve_pack_taken & btb_397_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_397_bht_T_4 = btb_397_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_397_bht_T_5 = io_i_branch_resolve_pack_taken & btb_397_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_397_bht_T_6 = btb_397_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_397_bht_T_7 = io_i_branch_resolve_pack_taken & btb_397_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_397_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_397_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_397_bht_T_13 = _btb_0_bht_T_8 & _btb_397_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_397_bht_T_16 = _btb_0_bht_T_8 & _btb_397_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_397_bht_T_19 = _btb_0_bht_T_8 & _btb_397_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_397_bht_T_20 = _btb_397_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_21 = _btb_397_bht_T_16 ? 2'h0 : _btb_397_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_22 = _btb_397_bht_T_13 ? 2'h0 : _btb_397_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_23 = _btb_397_bht_T_10 ? 2'h0 : _btb_397_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_24 = _btb_397_bht_T_7 ? 2'h3 : _btb_397_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_25 = _btb_397_bht_T_5 ? 2'h3 : _btb_397_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_26 = _btb_397_bht_T_3 ? 2'h3 : _btb_397_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_397_bht_T_27 = _btb_397_bht_T_1 ? 2'h1 : _btb_397_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10294 = btb_397_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7053; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10296 = btb_397_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_397_bht_T_27 : _GEN_8589; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_398_bht_T = btb_398_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_398_bht_T_1 = io_i_branch_resolve_pack_taken & btb_398_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_398_bht_T_2 = btb_398_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_398_bht_T_3 = io_i_branch_resolve_pack_taken & btb_398_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_398_bht_T_4 = btb_398_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_398_bht_T_5 = io_i_branch_resolve_pack_taken & btb_398_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_398_bht_T_6 = btb_398_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_398_bht_T_7 = io_i_branch_resolve_pack_taken & btb_398_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_398_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_398_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_398_bht_T_13 = _btb_0_bht_T_8 & _btb_398_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_398_bht_T_16 = _btb_0_bht_T_8 & _btb_398_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_398_bht_T_19 = _btb_0_bht_T_8 & _btb_398_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_398_bht_T_20 = _btb_398_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_21 = _btb_398_bht_T_16 ? 2'h0 : _btb_398_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_22 = _btb_398_bht_T_13 ? 2'h0 : _btb_398_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_23 = _btb_398_bht_T_10 ? 2'h0 : _btb_398_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_24 = _btb_398_bht_T_7 ? 2'h3 : _btb_398_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_25 = _btb_398_bht_T_5 ? 2'h3 : _btb_398_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_26 = _btb_398_bht_T_3 ? 2'h3 : _btb_398_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_398_bht_T_27 = _btb_398_bht_T_1 ? 2'h1 : _btb_398_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10298 = btb_398_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7054; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10300 = btb_398_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_398_bht_T_27 : _GEN_8590; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_399_bht_T = btb_399_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_399_bht_T_1 = io_i_branch_resolve_pack_taken & btb_399_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_399_bht_T_2 = btb_399_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_399_bht_T_3 = io_i_branch_resolve_pack_taken & btb_399_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_399_bht_T_4 = btb_399_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_399_bht_T_5 = io_i_branch_resolve_pack_taken & btb_399_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_399_bht_T_6 = btb_399_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_399_bht_T_7 = io_i_branch_resolve_pack_taken & btb_399_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_399_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_399_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_399_bht_T_13 = _btb_0_bht_T_8 & _btb_399_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_399_bht_T_16 = _btb_0_bht_T_8 & _btb_399_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_399_bht_T_19 = _btb_0_bht_T_8 & _btb_399_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_399_bht_T_20 = _btb_399_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_21 = _btb_399_bht_T_16 ? 2'h0 : _btb_399_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_22 = _btb_399_bht_T_13 ? 2'h0 : _btb_399_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_23 = _btb_399_bht_T_10 ? 2'h0 : _btb_399_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_24 = _btb_399_bht_T_7 ? 2'h3 : _btb_399_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_25 = _btb_399_bht_T_5 ? 2'h3 : _btb_399_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_26 = _btb_399_bht_T_3 ? 2'h3 : _btb_399_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_399_bht_T_27 = _btb_399_bht_T_1 ? 2'h1 : _btb_399_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10302 = btb_399_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7055; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10304 = btb_399_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_399_bht_T_27 : _GEN_8591; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_400_bht_T = btb_400_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_400_bht_T_1 = io_i_branch_resolve_pack_taken & btb_400_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_400_bht_T_2 = btb_400_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_400_bht_T_3 = io_i_branch_resolve_pack_taken & btb_400_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_400_bht_T_4 = btb_400_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_400_bht_T_5 = io_i_branch_resolve_pack_taken & btb_400_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_400_bht_T_6 = btb_400_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_400_bht_T_7 = io_i_branch_resolve_pack_taken & btb_400_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_400_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_400_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_400_bht_T_13 = _btb_0_bht_T_8 & _btb_400_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_400_bht_T_16 = _btb_0_bht_T_8 & _btb_400_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_400_bht_T_19 = _btb_0_bht_T_8 & _btb_400_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_400_bht_T_20 = _btb_400_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_21 = _btb_400_bht_T_16 ? 2'h0 : _btb_400_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_22 = _btb_400_bht_T_13 ? 2'h0 : _btb_400_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_23 = _btb_400_bht_T_10 ? 2'h0 : _btb_400_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_24 = _btb_400_bht_T_7 ? 2'h3 : _btb_400_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_25 = _btb_400_bht_T_5 ? 2'h3 : _btb_400_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_26 = _btb_400_bht_T_3 ? 2'h3 : _btb_400_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_400_bht_T_27 = _btb_400_bht_T_1 ? 2'h1 : _btb_400_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10306 = btb_400_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7056; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10308 = btb_400_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_400_bht_T_27 : _GEN_8592; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_401_bht_T = btb_401_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_401_bht_T_1 = io_i_branch_resolve_pack_taken & btb_401_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_401_bht_T_2 = btb_401_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_401_bht_T_3 = io_i_branch_resolve_pack_taken & btb_401_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_401_bht_T_4 = btb_401_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_401_bht_T_5 = io_i_branch_resolve_pack_taken & btb_401_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_401_bht_T_6 = btb_401_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_401_bht_T_7 = io_i_branch_resolve_pack_taken & btb_401_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_401_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_401_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_401_bht_T_13 = _btb_0_bht_T_8 & _btb_401_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_401_bht_T_16 = _btb_0_bht_T_8 & _btb_401_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_401_bht_T_19 = _btb_0_bht_T_8 & _btb_401_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_401_bht_T_20 = _btb_401_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_21 = _btb_401_bht_T_16 ? 2'h0 : _btb_401_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_22 = _btb_401_bht_T_13 ? 2'h0 : _btb_401_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_23 = _btb_401_bht_T_10 ? 2'h0 : _btb_401_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_24 = _btb_401_bht_T_7 ? 2'h3 : _btb_401_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_25 = _btb_401_bht_T_5 ? 2'h3 : _btb_401_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_26 = _btb_401_bht_T_3 ? 2'h3 : _btb_401_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_401_bht_T_27 = _btb_401_bht_T_1 ? 2'h1 : _btb_401_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10310 = btb_401_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7057; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10312 = btb_401_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_401_bht_T_27 : _GEN_8593; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_402_bht_T = btb_402_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_402_bht_T_1 = io_i_branch_resolve_pack_taken & btb_402_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_402_bht_T_2 = btb_402_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_402_bht_T_3 = io_i_branch_resolve_pack_taken & btb_402_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_402_bht_T_4 = btb_402_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_402_bht_T_5 = io_i_branch_resolve_pack_taken & btb_402_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_402_bht_T_6 = btb_402_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_402_bht_T_7 = io_i_branch_resolve_pack_taken & btb_402_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_402_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_402_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_402_bht_T_13 = _btb_0_bht_T_8 & _btb_402_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_402_bht_T_16 = _btb_0_bht_T_8 & _btb_402_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_402_bht_T_19 = _btb_0_bht_T_8 & _btb_402_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_402_bht_T_20 = _btb_402_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_21 = _btb_402_bht_T_16 ? 2'h0 : _btb_402_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_22 = _btb_402_bht_T_13 ? 2'h0 : _btb_402_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_23 = _btb_402_bht_T_10 ? 2'h0 : _btb_402_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_24 = _btb_402_bht_T_7 ? 2'h3 : _btb_402_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_25 = _btb_402_bht_T_5 ? 2'h3 : _btb_402_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_26 = _btb_402_bht_T_3 ? 2'h3 : _btb_402_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_402_bht_T_27 = _btb_402_bht_T_1 ? 2'h1 : _btb_402_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10314 = btb_402_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7058; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10316 = btb_402_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_402_bht_T_27 : _GEN_8594; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_403_bht_T = btb_403_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_403_bht_T_1 = io_i_branch_resolve_pack_taken & btb_403_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_403_bht_T_2 = btb_403_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_403_bht_T_3 = io_i_branch_resolve_pack_taken & btb_403_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_403_bht_T_4 = btb_403_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_403_bht_T_5 = io_i_branch_resolve_pack_taken & btb_403_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_403_bht_T_6 = btb_403_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_403_bht_T_7 = io_i_branch_resolve_pack_taken & btb_403_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_403_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_403_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_403_bht_T_13 = _btb_0_bht_T_8 & _btb_403_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_403_bht_T_16 = _btb_0_bht_T_8 & _btb_403_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_403_bht_T_19 = _btb_0_bht_T_8 & _btb_403_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_403_bht_T_20 = _btb_403_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_21 = _btb_403_bht_T_16 ? 2'h0 : _btb_403_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_22 = _btb_403_bht_T_13 ? 2'h0 : _btb_403_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_23 = _btb_403_bht_T_10 ? 2'h0 : _btb_403_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_24 = _btb_403_bht_T_7 ? 2'h3 : _btb_403_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_25 = _btb_403_bht_T_5 ? 2'h3 : _btb_403_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_26 = _btb_403_bht_T_3 ? 2'h3 : _btb_403_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_403_bht_T_27 = _btb_403_bht_T_1 ? 2'h1 : _btb_403_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10318 = btb_403_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7059; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10320 = btb_403_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_403_bht_T_27 : _GEN_8595; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_404_bht_T = btb_404_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_404_bht_T_1 = io_i_branch_resolve_pack_taken & btb_404_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_404_bht_T_2 = btb_404_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_404_bht_T_3 = io_i_branch_resolve_pack_taken & btb_404_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_404_bht_T_4 = btb_404_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_404_bht_T_5 = io_i_branch_resolve_pack_taken & btb_404_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_404_bht_T_6 = btb_404_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_404_bht_T_7 = io_i_branch_resolve_pack_taken & btb_404_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_404_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_404_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_404_bht_T_13 = _btb_0_bht_T_8 & _btb_404_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_404_bht_T_16 = _btb_0_bht_T_8 & _btb_404_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_404_bht_T_19 = _btb_0_bht_T_8 & _btb_404_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_404_bht_T_20 = _btb_404_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_21 = _btb_404_bht_T_16 ? 2'h0 : _btb_404_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_22 = _btb_404_bht_T_13 ? 2'h0 : _btb_404_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_23 = _btb_404_bht_T_10 ? 2'h0 : _btb_404_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_24 = _btb_404_bht_T_7 ? 2'h3 : _btb_404_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_25 = _btb_404_bht_T_5 ? 2'h3 : _btb_404_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_26 = _btb_404_bht_T_3 ? 2'h3 : _btb_404_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_404_bht_T_27 = _btb_404_bht_T_1 ? 2'h1 : _btb_404_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10321 = btb_404_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_403_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_402_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_401_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_400_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_399_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_398_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_397_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_396_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_395_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_394_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_393_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_392_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_391_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_390_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10261)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10322 = btb_404_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7060; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10324 = btb_404_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_404_bht_T_27 : _GEN_8596; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_405_bht_T = btb_405_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_405_bht_T_1 = io_i_branch_resolve_pack_taken & btb_405_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_405_bht_T_2 = btb_405_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_405_bht_T_3 = io_i_branch_resolve_pack_taken & btb_405_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_405_bht_T_4 = btb_405_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_405_bht_T_5 = io_i_branch_resolve_pack_taken & btb_405_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_405_bht_T_6 = btb_405_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_405_bht_T_7 = io_i_branch_resolve_pack_taken & btb_405_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_405_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_405_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_405_bht_T_13 = _btb_0_bht_T_8 & _btb_405_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_405_bht_T_16 = _btb_0_bht_T_8 & _btb_405_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_405_bht_T_19 = _btb_0_bht_T_8 & _btb_405_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_405_bht_T_20 = _btb_405_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_21 = _btb_405_bht_T_16 ? 2'h0 : _btb_405_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_22 = _btb_405_bht_T_13 ? 2'h0 : _btb_405_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_23 = _btb_405_bht_T_10 ? 2'h0 : _btb_405_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_24 = _btb_405_bht_T_7 ? 2'h3 : _btb_405_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_25 = _btb_405_bht_T_5 ? 2'h3 : _btb_405_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_26 = _btb_405_bht_T_3 ? 2'h3 : _btb_405_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_405_bht_T_27 = _btb_405_bht_T_1 ? 2'h1 : _btb_405_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10326 = btb_405_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7061; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10328 = btb_405_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_405_bht_T_27 : _GEN_8597; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_406_bht_T = btb_406_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_406_bht_T_1 = io_i_branch_resolve_pack_taken & btb_406_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_406_bht_T_2 = btb_406_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_406_bht_T_3 = io_i_branch_resolve_pack_taken & btb_406_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_406_bht_T_4 = btb_406_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_406_bht_T_5 = io_i_branch_resolve_pack_taken & btb_406_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_406_bht_T_6 = btb_406_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_406_bht_T_7 = io_i_branch_resolve_pack_taken & btb_406_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_406_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_406_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_406_bht_T_13 = _btb_0_bht_T_8 & _btb_406_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_406_bht_T_16 = _btb_0_bht_T_8 & _btb_406_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_406_bht_T_19 = _btb_0_bht_T_8 & _btb_406_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_406_bht_T_20 = _btb_406_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_21 = _btb_406_bht_T_16 ? 2'h0 : _btb_406_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_22 = _btb_406_bht_T_13 ? 2'h0 : _btb_406_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_23 = _btb_406_bht_T_10 ? 2'h0 : _btb_406_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_24 = _btb_406_bht_T_7 ? 2'h3 : _btb_406_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_25 = _btb_406_bht_T_5 ? 2'h3 : _btb_406_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_26 = _btb_406_bht_T_3 ? 2'h3 : _btb_406_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_406_bht_T_27 = _btb_406_bht_T_1 ? 2'h1 : _btb_406_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10330 = btb_406_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7062; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10332 = btb_406_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_406_bht_T_27 : _GEN_8598; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_407_bht_T = btb_407_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_407_bht_T_1 = io_i_branch_resolve_pack_taken & btb_407_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_407_bht_T_2 = btb_407_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_407_bht_T_3 = io_i_branch_resolve_pack_taken & btb_407_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_407_bht_T_4 = btb_407_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_407_bht_T_5 = io_i_branch_resolve_pack_taken & btb_407_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_407_bht_T_6 = btb_407_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_407_bht_T_7 = io_i_branch_resolve_pack_taken & btb_407_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_407_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_407_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_407_bht_T_13 = _btb_0_bht_T_8 & _btb_407_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_407_bht_T_16 = _btb_0_bht_T_8 & _btb_407_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_407_bht_T_19 = _btb_0_bht_T_8 & _btb_407_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_407_bht_T_20 = _btb_407_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_21 = _btb_407_bht_T_16 ? 2'h0 : _btb_407_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_22 = _btb_407_bht_T_13 ? 2'h0 : _btb_407_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_23 = _btb_407_bht_T_10 ? 2'h0 : _btb_407_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_24 = _btb_407_bht_T_7 ? 2'h3 : _btb_407_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_25 = _btb_407_bht_T_5 ? 2'h3 : _btb_407_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_26 = _btb_407_bht_T_3 ? 2'h3 : _btb_407_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_407_bht_T_27 = _btb_407_bht_T_1 ? 2'h1 : _btb_407_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10334 = btb_407_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7063; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10336 = btb_407_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_407_bht_T_27 : _GEN_8599; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_408_bht_T = btb_408_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_408_bht_T_1 = io_i_branch_resolve_pack_taken & btb_408_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_408_bht_T_2 = btb_408_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_408_bht_T_3 = io_i_branch_resolve_pack_taken & btb_408_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_408_bht_T_4 = btb_408_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_408_bht_T_5 = io_i_branch_resolve_pack_taken & btb_408_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_408_bht_T_6 = btb_408_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_408_bht_T_7 = io_i_branch_resolve_pack_taken & btb_408_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_408_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_408_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_408_bht_T_13 = _btb_0_bht_T_8 & _btb_408_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_408_bht_T_16 = _btb_0_bht_T_8 & _btb_408_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_408_bht_T_19 = _btb_0_bht_T_8 & _btb_408_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_408_bht_T_20 = _btb_408_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_21 = _btb_408_bht_T_16 ? 2'h0 : _btb_408_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_22 = _btb_408_bht_T_13 ? 2'h0 : _btb_408_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_23 = _btb_408_bht_T_10 ? 2'h0 : _btb_408_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_24 = _btb_408_bht_T_7 ? 2'h3 : _btb_408_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_25 = _btb_408_bht_T_5 ? 2'h3 : _btb_408_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_26 = _btb_408_bht_T_3 ? 2'h3 : _btb_408_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_408_bht_T_27 = _btb_408_bht_T_1 ? 2'h1 : _btb_408_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10338 = btb_408_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7064; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10340 = btb_408_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_408_bht_T_27 : _GEN_8600; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_409_bht_T = btb_409_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_409_bht_T_1 = io_i_branch_resolve_pack_taken & btb_409_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_409_bht_T_2 = btb_409_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_409_bht_T_3 = io_i_branch_resolve_pack_taken & btb_409_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_409_bht_T_4 = btb_409_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_409_bht_T_5 = io_i_branch_resolve_pack_taken & btb_409_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_409_bht_T_6 = btb_409_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_409_bht_T_7 = io_i_branch_resolve_pack_taken & btb_409_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_409_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_409_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_409_bht_T_13 = _btb_0_bht_T_8 & _btb_409_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_409_bht_T_16 = _btb_0_bht_T_8 & _btb_409_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_409_bht_T_19 = _btb_0_bht_T_8 & _btb_409_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_409_bht_T_20 = _btb_409_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_21 = _btb_409_bht_T_16 ? 2'h0 : _btb_409_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_22 = _btb_409_bht_T_13 ? 2'h0 : _btb_409_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_23 = _btb_409_bht_T_10 ? 2'h0 : _btb_409_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_24 = _btb_409_bht_T_7 ? 2'h3 : _btb_409_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_25 = _btb_409_bht_T_5 ? 2'h3 : _btb_409_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_26 = _btb_409_bht_T_3 ? 2'h3 : _btb_409_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_409_bht_T_27 = _btb_409_bht_T_1 ? 2'h1 : _btb_409_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10342 = btb_409_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7065; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10344 = btb_409_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_409_bht_T_27 : _GEN_8601; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_410_bht_T = btb_410_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_410_bht_T_1 = io_i_branch_resolve_pack_taken & btb_410_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_410_bht_T_2 = btb_410_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_410_bht_T_3 = io_i_branch_resolve_pack_taken & btb_410_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_410_bht_T_4 = btb_410_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_410_bht_T_5 = io_i_branch_resolve_pack_taken & btb_410_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_410_bht_T_6 = btb_410_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_410_bht_T_7 = io_i_branch_resolve_pack_taken & btb_410_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_410_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_410_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_410_bht_T_13 = _btb_0_bht_T_8 & _btb_410_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_410_bht_T_16 = _btb_0_bht_T_8 & _btb_410_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_410_bht_T_19 = _btb_0_bht_T_8 & _btb_410_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_410_bht_T_20 = _btb_410_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_21 = _btb_410_bht_T_16 ? 2'h0 : _btb_410_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_22 = _btb_410_bht_T_13 ? 2'h0 : _btb_410_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_23 = _btb_410_bht_T_10 ? 2'h0 : _btb_410_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_24 = _btb_410_bht_T_7 ? 2'h3 : _btb_410_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_25 = _btb_410_bht_T_5 ? 2'h3 : _btb_410_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_26 = _btb_410_bht_T_3 ? 2'h3 : _btb_410_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_410_bht_T_27 = _btb_410_bht_T_1 ? 2'h1 : _btb_410_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10346 = btb_410_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7066; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10348 = btb_410_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_410_bht_T_27 : _GEN_8602; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_411_bht_T = btb_411_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_411_bht_T_1 = io_i_branch_resolve_pack_taken & btb_411_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_411_bht_T_2 = btb_411_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_411_bht_T_3 = io_i_branch_resolve_pack_taken & btb_411_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_411_bht_T_4 = btb_411_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_411_bht_T_5 = io_i_branch_resolve_pack_taken & btb_411_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_411_bht_T_6 = btb_411_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_411_bht_T_7 = io_i_branch_resolve_pack_taken & btb_411_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_411_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_411_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_411_bht_T_13 = _btb_0_bht_T_8 & _btb_411_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_411_bht_T_16 = _btb_0_bht_T_8 & _btb_411_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_411_bht_T_19 = _btb_0_bht_T_8 & _btb_411_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_411_bht_T_20 = _btb_411_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_21 = _btb_411_bht_T_16 ? 2'h0 : _btb_411_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_22 = _btb_411_bht_T_13 ? 2'h0 : _btb_411_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_23 = _btb_411_bht_T_10 ? 2'h0 : _btb_411_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_24 = _btb_411_bht_T_7 ? 2'h3 : _btb_411_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_25 = _btb_411_bht_T_5 ? 2'h3 : _btb_411_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_26 = _btb_411_bht_T_3 ? 2'h3 : _btb_411_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_411_bht_T_27 = _btb_411_bht_T_1 ? 2'h1 : _btb_411_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10350 = btb_411_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7067; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10352 = btb_411_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_411_bht_T_27 : _GEN_8603; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_412_bht_T = btb_412_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_412_bht_T_1 = io_i_branch_resolve_pack_taken & btb_412_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_412_bht_T_2 = btb_412_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_412_bht_T_3 = io_i_branch_resolve_pack_taken & btb_412_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_412_bht_T_4 = btb_412_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_412_bht_T_5 = io_i_branch_resolve_pack_taken & btb_412_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_412_bht_T_6 = btb_412_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_412_bht_T_7 = io_i_branch_resolve_pack_taken & btb_412_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_412_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_412_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_412_bht_T_13 = _btb_0_bht_T_8 & _btb_412_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_412_bht_T_16 = _btb_0_bht_T_8 & _btb_412_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_412_bht_T_19 = _btb_0_bht_T_8 & _btb_412_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_412_bht_T_20 = _btb_412_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_21 = _btb_412_bht_T_16 ? 2'h0 : _btb_412_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_22 = _btb_412_bht_T_13 ? 2'h0 : _btb_412_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_23 = _btb_412_bht_T_10 ? 2'h0 : _btb_412_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_24 = _btb_412_bht_T_7 ? 2'h3 : _btb_412_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_25 = _btb_412_bht_T_5 ? 2'h3 : _btb_412_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_26 = _btb_412_bht_T_3 ? 2'h3 : _btb_412_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_412_bht_T_27 = _btb_412_bht_T_1 ? 2'h1 : _btb_412_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10354 = btb_412_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7068; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10356 = btb_412_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_412_bht_T_27 : _GEN_8604; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_413_bht_T = btb_413_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_413_bht_T_1 = io_i_branch_resolve_pack_taken & btb_413_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_413_bht_T_2 = btb_413_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_413_bht_T_3 = io_i_branch_resolve_pack_taken & btb_413_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_413_bht_T_4 = btb_413_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_413_bht_T_5 = io_i_branch_resolve_pack_taken & btb_413_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_413_bht_T_6 = btb_413_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_413_bht_T_7 = io_i_branch_resolve_pack_taken & btb_413_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_413_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_413_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_413_bht_T_13 = _btb_0_bht_T_8 & _btb_413_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_413_bht_T_16 = _btb_0_bht_T_8 & _btb_413_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_413_bht_T_19 = _btb_0_bht_T_8 & _btb_413_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_413_bht_T_20 = _btb_413_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_21 = _btb_413_bht_T_16 ? 2'h0 : _btb_413_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_22 = _btb_413_bht_T_13 ? 2'h0 : _btb_413_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_23 = _btb_413_bht_T_10 ? 2'h0 : _btb_413_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_24 = _btb_413_bht_T_7 ? 2'h3 : _btb_413_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_25 = _btb_413_bht_T_5 ? 2'h3 : _btb_413_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_26 = _btb_413_bht_T_3 ? 2'h3 : _btb_413_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_413_bht_T_27 = _btb_413_bht_T_1 ? 2'h1 : _btb_413_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10358 = btb_413_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7069; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10360 = btb_413_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_413_bht_T_27 : _GEN_8605; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_414_bht_T = btb_414_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_414_bht_T_1 = io_i_branch_resolve_pack_taken & btb_414_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_414_bht_T_2 = btb_414_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_414_bht_T_3 = io_i_branch_resolve_pack_taken & btb_414_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_414_bht_T_4 = btb_414_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_414_bht_T_5 = io_i_branch_resolve_pack_taken & btb_414_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_414_bht_T_6 = btb_414_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_414_bht_T_7 = io_i_branch_resolve_pack_taken & btb_414_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_414_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_414_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_414_bht_T_13 = _btb_0_bht_T_8 & _btb_414_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_414_bht_T_16 = _btb_0_bht_T_8 & _btb_414_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_414_bht_T_19 = _btb_0_bht_T_8 & _btb_414_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_414_bht_T_20 = _btb_414_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_21 = _btb_414_bht_T_16 ? 2'h0 : _btb_414_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_22 = _btb_414_bht_T_13 ? 2'h0 : _btb_414_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_23 = _btb_414_bht_T_10 ? 2'h0 : _btb_414_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_24 = _btb_414_bht_T_7 ? 2'h3 : _btb_414_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_25 = _btb_414_bht_T_5 ? 2'h3 : _btb_414_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_26 = _btb_414_bht_T_3 ? 2'h3 : _btb_414_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_414_bht_T_27 = _btb_414_bht_T_1 ? 2'h1 : _btb_414_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10362 = btb_414_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7070; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10364 = btb_414_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_414_bht_T_27 : _GEN_8606; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_415_bht_T = btb_415_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_415_bht_T_1 = io_i_branch_resolve_pack_taken & btb_415_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_415_bht_T_2 = btb_415_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_415_bht_T_3 = io_i_branch_resolve_pack_taken & btb_415_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_415_bht_T_4 = btb_415_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_415_bht_T_5 = io_i_branch_resolve_pack_taken & btb_415_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_415_bht_T_6 = btb_415_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_415_bht_T_7 = io_i_branch_resolve_pack_taken & btb_415_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_415_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_415_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_415_bht_T_13 = _btb_0_bht_T_8 & _btb_415_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_415_bht_T_16 = _btb_0_bht_T_8 & _btb_415_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_415_bht_T_19 = _btb_0_bht_T_8 & _btb_415_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_415_bht_T_20 = _btb_415_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_21 = _btb_415_bht_T_16 ? 2'h0 : _btb_415_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_22 = _btb_415_bht_T_13 ? 2'h0 : _btb_415_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_23 = _btb_415_bht_T_10 ? 2'h0 : _btb_415_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_24 = _btb_415_bht_T_7 ? 2'h3 : _btb_415_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_25 = _btb_415_bht_T_5 ? 2'h3 : _btb_415_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_26 = _btb_415_bht_T_3 ? 2'h3 : _btb_415_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_415_bht_T_27 = _btb_415_bht_T_1 ? 2'h1 : _btb_415_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10366 = btb_415_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7071; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10368 = btb_415_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_415_bht_T_27 : _GEN_8607; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_416_bht_T = btb_416_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_416_bht_T_1 = io_i_branch_resolve_pack_taken & btb_416_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_416_bht_T_2 = btb_416_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_416_bht_T_3 = io_i_branch_resolve_pack_taken & btb_416_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_416_bht_T_4 = btb_416_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_416_bht_T_5 = io_i_branch_resolve_pack_taken & btb_416_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_416_bht_T_6 = btb_416_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_416_bht_T_7 = io_i_branch_resolve_pack_taken & btb_416_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_416_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_416_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_416_bht_T_13 = _btb_0_bht_T_8 & _btb_416_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_416_bht_T_16 = _btb_0_bht_T_8 & _btb_416_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_416_bht_T_19 = _btb_0_bht_T_8 & _btb_416_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_416_bht_T_20 = _btb_416_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_21 = _btb_416_bht_T_16 ? 2'h0 : _btb_416_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_22 = _btb_416_bht_T_13 ? 2'h0 : _btb_416_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_23 = _btb_416_bht_T_10 ? 2'h0 : _btb_416_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_24 = _btb_416_bht_T_7 ? 2'h3 : _btb_416_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_25 = _btb_416_bht_T_5 ? 2'h3 : _btb_416_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_26 = _btb_416_bht_T_3 ? 2'h3 : _btb_416_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_416_bht_T_27 = _btb_416_bht_T_1 ? 2'h1 : _btb_416_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10370 = btb_416_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7072; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10372 = btb_416_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_416_bht_T_27 : _GEN_8608; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_417_bht_T = btb_417_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_417_bht_T_1 = io_i_branch_resolve_pack_taken & btb_417_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_417_bht_T_2 = btb_417_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_417_bht_T_3 = io_i_branch_resolve_pack_taken & btb_417_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_417_bht_T_4 = btb_417_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_417_bht_T_5 = io_i_branch_resolve_pack_taken & btb_417_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_417_bht_T_6 = btb_417_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_417_bht_T_7 = io_i_branch_resolve_pack_taken & btb_417_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_417_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_417_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_417_bht_T_13 = _btb_0_bht_T_8 & _btb_417_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_417_bht_T_16 = _btb_0_bht_T_8 & _btb_417_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_417_bht_T_19 = _btb_0_bht_T_8 & _btb_417_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_417_bht_T_20 = _btb_417_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_21 = _btb_417_bht_T_16 ? 2'h0 : _btb_417_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_22 = _btb_417_bht_T_13 ? 2'h0 : _btb_417_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_23 = _btb_417_bht_T_10 ? 2'h0 : _btb_417_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_24 = _btb_417_bht_T_7 ? 2'h3 : _btb_417_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_25 = _btb_417_bht_T_5 ? 2'h3 : _btb_417_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_26 = _btb_417_bht_T_3 ? 2'h3 : _btb_417_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_417_bht_T_27 = _btb_417_bht_T_1 ? 2'h1 : _btb_417_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10374 = btb_417_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7073; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10376 = btb_417_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_417_bht_T_27 : _GEN_8609; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_418_bht_T = btb_418_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_418_bht_T_1 = io_i_branch_resolve_pack_taken & btb_418_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_418_bht_T_2 = btb_418_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_418_bht_T_3 = io_i_branch_resolve_pack_taken & btb_418_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_418_bht_T_4 = btb_418_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_418_bht_T_5 = io_i_branch_resolve_pack_taken & btb_418_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_418_bht_T_6 = btb_418_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_418_bht_T_7 = io_i_branch_resolve_pack_taken & btb_418_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_418_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_418_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_418_bht_T_13 = _btb_0_bht_T_8 & _btb_418_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_418_bht_T_16 = _btb_0_bht_T_8 & _btb_418_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_418_bht_T_19 = _btb_0_bht_T_8 & _btb_418_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_418_bht_T_20 = _btb_418_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_21 = _btb_418_bht_T_16 ? 2'h0 : _btb_418_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_22 = _btb_418_bht_T_13 ? 2'h0 : _btb_418_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_23 = _btb_418_bht_T_10 ? 2'h0 : _btb_418_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_24 = _btb_418_bht_T_7 ? 2'h3 : _btb_418_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_25 = _btb_418_bht_T_5 ? 2'h3 : _btb_418_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_26 = _btb_418_bht_T_3 ? 2'h3 : _btb_418_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_418_bht_T_27 = _btb_418_bht_T_1 ? 2'h1 : _btb_418_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10378 = btb_418_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7074; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10380 = btb_418_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_418_bht_T_27 : _GEN_8610; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_419_bht_T = btb_419_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_419_bht_T_1 = io_i_branch_resolve_pack_taken & btb_419_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_419_bht_T_2 = btb_419_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_419_bht_T_3 = io_i_branch_resolve_pack_taken & btb_419_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_419_bht_T_4 = btb_419_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_419_bht_T_5 = io_i_branch_resolve_pack_taken & btb_419_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_419_bht_T_6 = btb_419_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_419_bht_T_7 = io_i_branch_resolve_pack_taken & btb_419_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_419_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_419_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_419_bht_T_13 = _btb_0_bht_T_8 & _btb_419_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_419_bht_T_16 = _btb_0_bht_T_8 & _btb_419_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_419_bht_T_19 = _btb_0_bht_T_8 & _btb_419_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_419_bht_T_20 = _btb_419_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_21 = _btb_419_bht_T_16 ? 2'h0 : _btb_419_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_22 = _btb_419_bht_T_13 ? 2'h0 : _btb_419_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_23 = _btb_419_bht_T_10 ? 2'h0 : _btb_419_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_24 = _btb_419_bht_T_7 ? 2'h3 : _btb_419_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_25 = _btb_419_bht_T_5 ? 2'h3 : _btb_419_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_26 = _btb_419_bht_T_3 ? 2'h3 : _btb_419_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_419_bht_T_27 = _btb_419_bht_T_1 ? 2'h1 : _btb_419_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10381 = btb_419_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_418_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_417_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_416_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_415_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_414_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_413_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_412_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_411_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_410_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_409_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_408_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_407_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_406_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_405_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10321)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10382 = btb_419_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7075; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10384 = btb_419_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_419_bht_T_27 : _GEN_8611; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_420_bht_T = btb_420_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_420_bht_T_1 = io_i_branch_resolve_pack_taken & btb_420_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_420_bht_T_2 = btb_420_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_420_bht_T_3 = io_i_branch_resolve_pack_taken & btb_420_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_420_bht_T_4 = btb_420_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_420_bht_T_5 = io_i_branch_resolve_pack_taken & btb_420_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_420_bht_T_6 = btb_420_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_420_bht_T_7 = io_i_branch_resolve_pack_taken & btb_420_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_420_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_420_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_420_bht_T_13 = _btb_0_bht_T_8 & _btb_420_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_420_bht_T_16 = _btb_0_bht_T_8 & _btb_420_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_420_bht_T_19 = _btb_0_bht_T_8 & _btb_420_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_420_bht_T_20 = _btb_420_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_21 = _btb_420_bht_T_16 ? 2'h0 : _btb_420_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_22 = _btb_420_bht_T_13 ? 2'h0 : _btb_420_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_23 = _btb_420_bht_T_10 ? 2'h0 : _btb_420_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_24 = _btb_420_bht_T_7 ? 2'h3 : _btb_420_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_25 = _btb_420_bht_T_5 ? 2'h3 : _btb_420_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_26 = _btb_420_bht_T_3 ? 2'h3 : _btb_420_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_420_bht_T_27 = _btb_420_bht_T_1 ? 2'h1 : _btb_420_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10386 = btb_420_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7076; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10388 = btb_420_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_420_bht_T_27 : _GEN_8612; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_421_bht_T = btb_421_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_421_bht_T_1 = io_i_branch_resolve_pack_taken & btb_421_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_421_bht_T_2 = btb_421_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_421_bht_T_3 = io_i_branch_resolve_pack_taken & btb_421_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_421_bht_T_4 = btb_421_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_421_bht_T_5 = io_i_branch_resolve_pack_taken & btb_421_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_421_bht_T_6 = btb_421_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_421_bht_T_7 = io_i_branch_resolve_pack_taken & btb_421_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_421_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_421_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_421_bht_T_13 = _btb_0_bht_T_8 & _btb_421_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_421_bht_T_16 = _btb_0_bht_T_8 & _btb_421_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_421_bht_T_19 = _btb_0_bht_T_8 & _btb_421_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_421_bht_T_20 = _btb_421_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_21 = _btb_421_bht_T_16 ? 2'h0 : _btb_421_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_22 = _btb_421_bht_T_13 ? 2'h0 : _btb_421_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_23 = _btb_421_bht_T_10 ? 2'h0 : _btb_421_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_24 = _btb_421_bht_T_7 ? 2'h3 : _btb_421_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_25 = _btb_421_bht_T_5 ? 2'h3 : _btb_421_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_26 = _btb_421_bht_T_3 ? 2'h3 : _btb_421_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_421_bht_T_27 = _btb_421_bht_T_1 ? 2'h1 : _btb_421_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10390 = btb_421_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7077; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10392 = btb_421_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_421_bht_T_27 : _GEN_8613; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_422_bht_T = btb_422_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_422_bht_T_1 = io_i_branch_resolve_pack_taken & btb_422_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_422_bht_T_2 = btb_422_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_422_bht_T_3 = io_i_branch_resolve_pack_taken & btb_422_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_422_bht_T_4 = btb_422_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_422_bht_T_5 = io_i_branch_resolve_pack_taken & btb_422_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_422_bht_T_6 = btb_422_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_422_bht_T_7 = io_i_branch_resolve_pack_taken & btb_422_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_422_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_422_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_422_bht_T_13 = _btb_0_bht_T_8 & _btb_422_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_422_bht_T_16 = _btb_0_bht_T_8 & _btb_422_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_422_bht_T_19 = _btb_0_bht_T_8 & _btb_422_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_422_bht_T_20 = _btb_422_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_21 = _btb_422_bht_T_16 ? 2'h0 : _btb_422_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_22 = _btb_422_bht_T_13 ? 2'h0 : _btb_422_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_23 = _btb_422_bht_T_10 ? 2'h0 : _btb_422_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_24 = _btb_422_bht_T_7 ? 2'h3 : _btb_422_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_25 = _btb_422_bht_T_5 ? 2'h3 : _btb_422_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_26 = _btb_422_bht_T_3 ? 2'h3 : _btb_422_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_422_bht_T_27 = _btb_422_bht_T_1 ? 2'h1 : _btb_422_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10394 = btb_422_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7078; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10396 = btb_422_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_422_bht_T_27 : _GEN_8614; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_423_bht_T = btb_423_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_423_bht_T_1 = io_i_branch_resolve_pack_taken & btb_423_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_423_bht_T_2 = btb_423_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_423_bht_T_3 = io_i_branch_resolve_pack_taken & btb_423_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_423_bht_T_4 = btb_423_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_423_bht_T_5 = io_i_branch_resolve_pack_taken & btb_423_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_423_bht_T_6 = btb_423_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_423_bht_T_7 = io_i_branch_resolve_pack_taken & btb_423_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_423_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_423_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_423_bht_T_13 = _btb_0_bht_T_8 & _btb_423_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_423_bht_T_16 = _btb_0_bht_T_8 & _btb_423_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_423_bht_T_19 = _btb_0_bht_T_8 & _btb_423_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_423_bht_T_20 = _btb_423_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_21 = _btb_423_bht_T_16 ? 2'h0 : _btb_423_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_22 = _btb_423_bht_T_13 ? 2'h0 : _btb_423_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_23 = _btb_423_bht_T_10 ? 2'h0 : _btb_423_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_24 = _btb_423_bht_T_7 ? 2'h3 : _btb_423_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_25 = _btb_423_bht_T_5 ? 2'h3 : _btb_423_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_26 = _btb_423_bht_T_3 ? 2'h3 : _btb_423_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_423_bht_T_27 = _btb_423_bht_T_1 ? 2'h1 : _btb_423_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10398 = btb_423_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7079; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10400 = btb_423_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_423_bht_T_27 : _GEN_8615; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_424_bht_T = btb_424_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_424_bht_T_1 = io_i_branch_resolve_pack_taken & btb_424_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_424_bht_T_2 = btb_424_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_424_bht_T_3 = io_i_branch_resolve_pack_taken & btb_424_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_424_bht_T_4 = btb_424_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_424_bht_T_5 = io_i_branch_resolve_pack_taken & btb_424_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_424_bht_T_6 = btb_424_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_424_bht_T_7 = io_i_branch_resolve_pack_taken & btb_424_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_424_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_424_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_424_bht_T_13 = _btb_0_bht_T_8 & _btb_424_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_424_bht_T_16 = _btb_0_bht_T_8 & _btb_424_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_424_bht_T_19 = _btb_0_bht_T_8 & _btb_424_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_424_bht_T_20 = _btb_424_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_21 = _btb_424_bht_T_16 ? 2'h0 : _btb_424_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_22 = _btb_424_bht_T_13 ? 2'h0 : _btb_424_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_23 = _btb_424_bht_T_10 ? 2'h0 : _btb_424_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_24 = _btb_424_bht_T_7 ? 2'h3 : _btb_424_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_25 = _btb_424_bht_T_5 ? 2'h3 : _btb_424_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_26 = _btb_424_bht_T_3 ? 2'h3 : _btb_424_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_424_bht_T_27 = _btb_424_bht_T_1 ? 2'h1 : _btb_424_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10402 = btb_424_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7080; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10404 = btb_424_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_424_bht_T_27 : _GEN_8616; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_425_bht_T = btb_425_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_425_bht_T_1 = io_i_branch_resolve_pack_taken & btb_425_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_425_bht_T_2 = btb_425_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_425_bht_T_3 = io_i_branch_resolve_pack_taken & btb_425_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_425_bht_T_4 = btb_425_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_425_bht_T_5 = io_i_branch_resolve_pack_taken & btb_425_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_425_bht_T_6 = btb_425_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_425_bht_T_7 = io_i_branch_resolve_pack_taken & btb_425_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_425_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_425_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_425_bht_T_13 = _btb_0_bht_T_8 & _btb_425_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_425_bht_T_16 = _btb_0_bht_T_8 & _btb_425_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_425_bht_T_19 = _btb_0_bht_T_8 & _btb_425_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_425_bht_T_20 = _btb_425_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_21 = _btb_425_bht_T_16 ? 2'h0 : _btb_425_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_22 = _btb_425_bht_T_13 ? 2'h0 : _btb_425_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_23 = _btb_425_bht_T_10 ? 2'h0 : _btb_425_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_24 = _btb_425_bht_T_7 ? 2'h3 : _btb_425_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_25 = _btb_425_bht_T_5 ? 2'h3 : _btb_425_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_26 = _btb_425_bht_T_3 ? 2'h3 : _btb_425_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_425_bht_T_27 = _btb_425_bht_T_1 ? 2'h1 : _btb_425_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10406 = btb_425_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7081; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10408 = btb_425_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_425_bht_T_27 : _GEN_8617; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_426_bht_T = btb_426_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_426_bht_T_1 = io_i_branch_resolve_pack_taken & btb_426_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_426_bht_T_2 = btb_426_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_426_bht_T_3 = io_i_branch_resolve_pack_taken & btb_426_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_426_bht_T_4 = btb_426_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_426_bht_T_5 = io_i_branch_resolve_pack_taken & btb_426_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_426_bht_T_6 = btb_426_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_426_bht_T_7 = io_i_branch_resolve_pack_taken & btb_426_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_426_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_426_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_426_bht_T_13 = _btb_0_bht_T_8 & _btb_426_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_426_bht_T_16 = _btb_0_bht_T_8 & _btb_426_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_426_bht_T_19 = _btb_0_bht_T_8 & _btb_426_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_426_bht_T_20 = _btb_426_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_21 = _btb_426_bht_T_16 ? 2'h0 : _btb_426_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_22 = _btb_426_bht_T_13 ? 2'h0 : _btb_426_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_23 = _btb_426_bht_T_10 ? 2'h0 : _btb_426_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_24 = _btb_426_bht_T_7 ? 2'h3 : _btb_426_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_25 = _btb_426_bht_T_5 ? 2'h3 : _btb_426_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_26 = _btb_426_bht_T_3 ? 2'h3 : _btb_426_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_426_bht_T_27 = _btb_426_bht_T_1 ? 2'h1 : _btb_426_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10410 = btb_426_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7082; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10412 = btb_426_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_426_bht_T_27 : _GEN_8618; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_427_bht_T = btb_427_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_427_bht_T_1 = io_i_branch_resolve_pack_taken & btb_427_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_427_bht_T_2 = btb_427_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_427_bht_T_3 = io_i_branch_resolve_pack_taken & btb_427_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_427_bht_T_4 = btb_427_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_427_bht_T_5 = io_i_branch_resolve_pack_taken & btb_427_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_427_bht_T_6 = btb_427_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_427_bht_T_7 = io_i_branch_resolve_pack_taken & btb_427_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_427_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_427_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_427_bht_T_13 = _btb_0_bht_T_8 & _btb_427_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_427_bht_T_16 = _btb_0_bht_T_8 & _btb_427_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_427_bht_T_19 = _btb_0_bht_T_8 & _btb_427_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_427_bht_T_20 = _btb_427_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_21 = _btb_427_bht_T_16 ? 2'h0 : _btb_427_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_22 = _btb_427_bht_T_13 ? 2'h0 : _btb_427_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_23 = _btb_427_bht_T_10 ? 2'h0 : _btb_427_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_24 = _btb_427_bht_T_7 ? 2'h3 : _btb_427_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_25 = _btb_427_bht_T_5 ? 2'h3 : _btb_427_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_26 = _btb_427_bht_T_3 ? 2'h3 : _btb_427_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_427_bht_T_27 = _btb_427_bht_T_1 ? 2'h1 : _btb_427_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10414 = btb_427_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7083; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10416 = btb_427_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_427_bht_T_27 : _GEN_8619; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_428_bht_T = btb_428_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_428_bht_T_1 = io_i_branch_resolve_pack_taken & btb_428_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_428_bht_T_2 = btb_428_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_428_bht_T_3 = io_i_branch_resolve_pack_taken & btb_428_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_428_bht_T_4 = btb_428_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_428_bht_T_5 = io_i_branch_resolve_pack_taken & btb_428_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_428_bht_T_6 = btb_428_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_428_bht_T_7 = io_i_branch_resolve_pack_taken & btb_428_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_428_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_428_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_428_bht_T_13 = _btb_0_bht_T_8 & _btb_428_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_428_bht_T_16 = _btb_0_bht_T_8 & _btb_428_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_428_bht_T_19 = _btb_0_bht_T_8 & _btb_428_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_428_bht_T_20 = _btb_428_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_21 = _btb_428_bht_T_16 ? 2'h0 : _btb_428_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_22 = _btb_428_bht_T_13 ? 2'h0 : _btb_428_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_23 = _btb_428_bht_T_10 ? 2'h0 : _btb_428_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_24 = _btb_428_bht_T_7 ? 2'h3 : _btb_428_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_25 = _btb_428_bht_T_5 ? 2'h3 : _btb_428_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_26 = _btb_428_bht_T_3 ? 2'h3 : _btb_428_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_428_bht_T_27 = _btb_428_bht_T_1 ? 2'h1 : _btb_428_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10418 = btb_428_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7084; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10420 = btb_428_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_428_bht_T_27 : _GEN_8620; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_429_bht_T = btb_429_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_429_bht_T_1 = io_i_branch_resolve_pack_taken & btb_429_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_429_bht_T_2 = btb_429_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_429_bht_T_3 = io_i_branch_resolve_pack_taken & btb_429_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_429_bht_T_4 = btb_429_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_429_bht_T_5 = io_i_branch_resolve_pack_taken & btb_429_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_429_bht_T_6 = btb_429_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_429_bht_T_7 = io_i_branch_resolve_pack_taken & btb_429_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_429_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_429_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_429_bht_T_13 = _btb_0_bht_T_8 & _btb_429_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_429_bht_T_16 = _btb_0_bht_T_8 & _btb_429_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_429_bht_T_19 = _btb_0_bht_T_8 & _btb_429_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_429_bht_T_20 = _btb_429_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_21 = _btb_429_bht_T_16 ? 2'h0 : _btb_429_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_22 = _btb_429_bht_T_13 ? 2'h0 : _btb_429_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_23 = _btb_429_bht_T_10 ? 2'h0 : _btb_429_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_24 = _btb_429_bht_T_7 ? 2'h3 : _btb_429_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_25 = _btb_429_bht_T_5 ? 2'h3 : _btb_429_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_26 = _btb_429_bht_T_3 ? 2'h3 : _btb_429_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_429_bht_T_27 = _btb_429_bht_T_1 ? 2'h1 : _btb_429_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10422 = btb_429_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7085; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10424 = btb_429_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_429_bht_T_27 : _GEN_8621; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_430_bht_T = btb_430_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_430_bht_T_1 = io_i_branch_resolve_pack_taken & btb_430_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_430_bht_T_2 = btb_430_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_430_bht_T_3 = io_i_branch_resolve_pack_taken & btb_430_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_430_bht_T_4 = btb_430_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_430_bht_T_5 = io_i_branch_resolve_pack_taken & btb_430_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_430_bht_T_6 = btb_430_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_430_bht_T_7 = io_i_branch_resolve_pack_taken & btb_430_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_430_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_430_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_430_bht_T_13 = _btb_0_bht_T_8 & _btb_430_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_430_bht_T_16 = _btb_0_bht_T_8 & _btb_430_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_430_bht_T_19 = _btb_0_bht_T_8 & _btb_430_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_430_bht_T_20 = _btb_430_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_21 = _btb_430_bht_T_16 ? 2'h0 : _btb_430_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_22 = _btb_430_bht_T_13 ? 2'h0 : _btb_430_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_23 = _btb_430_bht_T_10 ? 2'h0 : _btb_430_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_24 = _btb_430_bht_T_7 ? 2'h3 : _btb_430_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_25 = _btb_430_bht_T_5 ? 2'h3 : _btb_430_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_26 = _btb_430_bht_T_3 ? 2'h3 : _btb_430_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_430_bht_T_27 = _btb_430_bht_T_1 ? 2'h1 : _btb_430_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10426 = btb_430_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7086; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10428 = btb_430_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_430_bht_T_27 : _GEN_8622; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_431_bht_T = btb_431_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_431_bht_T_1 = io_i_branch_resolve_pack_taken & btb_431_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_431_bht_T_2 = btb_431_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_431_bht_T_3 = io_i_branch_resolve_pack_taken & btb_431_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_431_bht_T_4 = btb_431_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_431_bht_T_5 = io_i_branch_resolve_pack_taken & btb_431_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_431_bht_T_6 = btb_431_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_431_bht_T_7 = io_i_branch_resolve_pack_taken & btb_431_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_431_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_431_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_431_bht_T_13 = _btb_0_bht_T_8 & _btb_431_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_431_bht_T_16 = _btb_0_bht_T_8 & _btb_431_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_431_bht_T_19 = _btb_0_bht_T_8 & _btb_431_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_431_bht_T_20 = _btb_431_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_21 = _btb_431_bht_T_16 ? 2'h0 : _btb_431_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_22 = _btb_431_bht_T_13 ? 2'h0 : _btb_431_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_23 = _btb_431_bht_T_10 ? 2'h0 : _btb_431_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_24 = _btb_431_bht_T_7 ? 2'h3 : _btb_431_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_25 = _btb_431_bht_T_5 ? 2'h3 : _btb_431_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_26 = _btb_431_bht_T_3 ? 2'h3 : _btb_431_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_431_bht_T_27 = _btb_431_bht_T_1 ? 2'h1 : _btb_431_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10430 = btb_431_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7087; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10432 = btb_431_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_431_bht_T_27 : _GEN_8623; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_432_bht_T = btb_432_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_432_bht_T_1 = io_i_branch_resolve_pack_taken & btb_432_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_432_bht_T_2 = btb_432_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_432_bht_T_3 = io_i_branch_resolve_pack_taken & btb_432_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_432_bht_T_4 = btb_432_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_432_bht_T_5 = io_i_branch_resolve_pack_taken & btb_432_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_432_bht_T_6 = btb_432_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_432_bht_T_7 = io_i_branch_resolve_pack_taken & btb_432_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_432_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_432_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_432_bht_T_13 = _btb_0_bht_T_8 & _btb_432_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_432_bht_T_16 = _btb_0_bht_T_8 & _btb_432_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_432_bht_T_19 = _btb_0_bht_T_8 & _btb_432_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_432_bht_T_20 = _btb_432_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_21 = _btb_432_bht_T_16 ? 2'h0 : _btb_432_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_22 = _btb_432_bht_T_13 ? 2'h0 : _btb_432_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_23 = _btb_432_bht_T_10 ? 2'h0 : _btb_432_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_24 = _btb_432_bht_T_7 ? 2'h3 : _btb_432_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_25 = _btb_432_bht_T_5 ? 2'h3 : _btb_432_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_26 = _btb_432_bht_T_3 ? 2'h3 : _btb_432_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_432_bht_T_27 = _btb_432_bht_T_1 ? 2'h1 : _btb_432_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10434 = btb_432_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7088; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10436 = btb_432_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_432_bht_T_27 : _GEN_8624; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_433_bht_T = btb_433_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_433_bht_T_1 = io_i_branch_resolve_pack_taken & btb_433_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_433_bht_T_2 = btb_433_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_433_bht_T_3 = io_i_branch_resolve_pack_taken & btb_433_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_433_bht_T_4 = btb_433_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_433_bht_T_5 = io_i_branch_resolve_pack_taken & btb_433_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_433_bht_T_6 = btb_433_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_433_bht_T_7 = io_i_branch_resolve_pack_taken & btb_433_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_433_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_433_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_433_bht_T_13 = _btb_0_bht_T_8 & _btb_433_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_433_bht_T_16 = _btb_0_bht_T_8 & _btb_433_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_433_bht_T_19 = _btb_0_bht_T_8 & _btb_433_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_433_bht_T_20 = _btb_433_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_21 = _btb_433_bht_T_16 ? 2'h0 : _btb_433_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_22 = _btb_433_bht_T_13 ? 2'h0 : _btb_433_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_23 = _btb_433_bht_T_10 ? 2'h0 : _btb_433_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_24 = _btb_433_bht_T_7 ? 2'h3 : _btb_433_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_25 = _btb_433_bht_T_5 ? 2'h3 : _btb_433_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_26 = _btb_433_bht_T_3 ? 2'h3 : _btb_433_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_433_bht_T_27 = _btb_433_bht_T_1 ? 2'h1 : _btb_433_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10438 = btb_433_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7089; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10440 = btb_433_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_433_bht_T_27 : _GEN_8625; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_434_bht_T = btb_434_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_434_bht_T_1 = io_i_branch_resolve_pack_taken & btb_434_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_434_bht_T_2 = btb_434_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_434_bht_T_3 = io_i_branch_resolve_pack_taken & btb_434_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_434_bht_T_4 = btb_434_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_434_bht_T_5 = io_i_branch_resolve_pack_taken & btb_434_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_434_bht_T_6 = btb_434_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_434_bht_T_7 = io_i_branch_resolve_pack_taken & btb_434_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_434_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_434_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_434_bht_T_13 = _btb_0_bht_T_8 & _btb_434_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_434_bht_T_16 = _btb_0_bht_T_8 & _btb_434_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_434_bht_T_19 = _btb_0_bht_T_8 & _btb_434_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_434_bht_T_20 = _btb_434_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_21 = _btb_434_bht_T_16 ? 2'h0 : _btb_434_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_22 = _btb_434_bht_T_13 ? 2'h0 : _btb_434_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_23 = _btb_434_bht_T_10 ? 2'h0 : _btb_434_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_24 = _btb_434_bht_T_7 ? 2'h3 : _btb_434_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_25 = _btb_434_bht_T_5 ? 2'h3 : _btb_434_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_26 = _btb_434_bht_T_3 ? 2'h3 : _btb_434_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_434_bht_T_27 = _btb_434_bht_T_1 ? 2'h1 : _btb_434_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10441 = btb_434_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_433_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_432_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_431_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_430_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_429_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_428_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_427_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_426_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_425_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_424_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_423_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_422_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_421_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_420_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10381)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10442 = btb_434_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7090; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10444 = btb_434_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_434_bht_T_27 : _GEN_8626; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_435_bht_T = btb_435_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_435_bht_T_1 = io_i_branch_resolve_pack_taken & btb_435_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_435_bht_T_2 = btb_435_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_435_bht_T_3 = io_i_branch_resolve_pack_taken & btb_435_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_435_bht_T_4 = btb_435_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_435_bht_T_5 = io_i_branch_resolve_pack_taken & btb_435_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_435_bht_T_6 = btb_435_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_435_bht_T_7 = io_i_branch_resolve_pack_taken & btb_435_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_435_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_435_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_435_bht_T_13 = _btb_0_bht_T_8 & _btb_435_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_435_bht_T_16 = _btb_0_bht_T_8 & _btb_435_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_435_bht_T_19 = _btb_0_bht_T_8 & _btb_435_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_435_bht_T_20 = _btb_435_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_21 = _btb_435_bht_T_16 ? 2'h0 : _btb_435_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_22 = _btb_435_bht_T_13 ? 2'h0 : _btb_435_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_23 = _btb_435_bht_T_10 ? 2'h0 : _btb_435_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_24 = _btb_435_bht_T_7 ? 2'h3 : _btb_435_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_25 = _btb_435_bht_T_5 ? 2'h3 : _btb_435_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_26 = _btb_435_bht_T_3 ? 2'h3 : _btb_435_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_435_bht_T_27 = _btb_435_bht_T_1 ? 2'h1 : _btb_435_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10446 = btb_435_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7091; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10448 = btb_435_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_435_bht_T_27 : _GEN_8627; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_436_bht_T = btb_436_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_436_bht_T_1 = io_i_branch_resolve_pack_taken & btb_436_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_436_bht_T_2 = btb_436_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_436_bht_T_3 = io_i_branch_resolve_pack_taken & btb_436_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_436_bht_T_4 = btb_436_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_436_bht_T_5 = io_i_branch_resolve_pack_taken & btb_436_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_436_bht_T_6 = btb_436_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_436_bht_T_7 = io_i_branch_resolve_pack_taken & btb_436_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_436_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_436_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_436_bht_T_13 = _btb_0_bht_T_8 & _btb_436_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_436_bht_T_16 = _btb_0_bht_T_8 & _btb_436_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_436_bht_T_19 = _btb_0_bht_T_8 & _btb_436_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_436_bht_T_20 = _btb_436_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_21 = _btb_436_bht_T_16 ? 2'h0 : _btb_436_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_22 = _btb_436_bht_T_13 ? 2'h0 : _btb_436_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_23 = _btb_436_bht_T_10 ? 2'h0 : _btb_436_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_24 = _btb_436_bht_T_7 ? 2'h3 : _btb_436_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_25 = _btb_436_bht_T_5 ? 2'h3 : _btb_436_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_26 = _btb_436_bht_T_3 ? 2'h3 : _btb_436_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_436_bht_T_27 = _btb_436_bht_T_1 ? 2'h1 : _btb_436_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10450 = btb_436_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7092; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10452 = btb_436_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_436_bht_T_27 : _GEN_8628; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_437_bht_T = btb_437_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_437_bht_T_1 = io_i_branch_resolve_pack_taken & btb_437_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_437_bht_T_2 = btb_437_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_437_bht_T_3 = io_i_branch_resolve_pack_taken & btb_437_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_437_bht_T_4 = btb_437_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_437_bht_T_5 = io_i_branch_resolve_pack_taken & btb_437_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_437_bht_T_6 = btb_437_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_437_bht_T_7 = io_i_branch_resolve_pack_taken & btb_437_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_437_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_437_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_437_bht_T_13 = _btb_0_bht_T_8 & _btb_437_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_437_bht_T_16 = _btb_0_bht_T_8 & _btb_437_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_437_bht_T_19 = _btb_0_bht_T_8 & _btb_437_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_437_bht_T_20 = _btb_437_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_21 = _btb_437_bht_T_16 ? 2'h0 : _btb_437_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_22 = _btb_437_bht_T_13 ? 2'h0 : _btb_437_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_23 = _btb_437_bht_T_10 ? 2'h0 : _btb_437_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_24 = _btb_437_bht_T_7 ? 2'h3 : _btb_437_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_25 = _btb_437_bht_T_5 ? 2'h3 : _btb_437_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_26 = _btb_437_bht_T_3 ? 2'h3 : _btb_437_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_437_bht_T_27 = _btb_437_bht_T_1 ? 2'h1 : _btb_437_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10454 = btb_437_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7093; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10456 = btb_437_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_437_bht_T_27 : _GEN_8629; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_438_bht_T = btb_438_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_438_bht_T_1 = io_i_branch_resolve_pack_taken & btb_438_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_438_bht_T_2 = btb_438_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_438_bht_T_3 = io_i_branch_resolve_pack_taken & btb_438_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_438_bht_T_4 = btb_438_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_438_bht_T_5 = io_i_branch_resolve_pack_taken & btb_438_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_438_bht_T_6 = btb_438_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_438_bht_T_7 = io_i_branch_resolve_pack_taken & btb_438_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_438_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_438_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_438_bht_T_13 = _btb_0_bht_T_8 & _btb_438_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_438_bht_T_16 = _btb_0_bht_T_8 & _btb_438_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_438_bht_T_19 = _btb_0_bht_T_8 & _btb_438_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_438_bht_T_20 = _btb_438_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_21 = _btb_438_bht_T_16 ? 2'h0 : _btb_438_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_22 = _btb_438_bht_T_13 ? 2'h0 : _btb_438_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_23 = _btb_438_bht_T_10 ? 2'h0 : _btb_438_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_24 = _btb_438_bht_T_7 ? 2'h3 : _btb_438_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_25 = _btb_438_bht_T_5 ? 2'h3 : _btb_438_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_26 = _btb_438_bht_T_3 ? 2'h3 : _btb_438_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_438_bht_T_27 = _btb_438_bht_T_1 ? 2'h1 : _btb_438_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10458 = btb_438_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7094; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10460 = btb_438_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_438_bht_T_27 : _GEN_8630; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_439_bht_T = btb_439_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_439_bht_T_1 = io_i_branch_resolve_pack_taken & btb_439_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_439_bht_T_2 = btb_439_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_439_bht_T_3 = io_i_branch_resolve_pack_taken & btb_439_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_439_bht_T_4 = btb_439_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_439_bht_T_5 = io_i_branch_resolve_pack_taken & btb_439_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_439_bht_T_6 = btb_439_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_439_bht_T_7 = io_i_branch_resolve_pack_taken & btb_439_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_439_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_439_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_439_bht_T_13 = _btb_0_bht_T_8 & _btb_439_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_439_bht_T_16 = _btb_0_bht_T_8 & _btb_439_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_439_bht_T_19 = _btb_0_bht_T_8 & _btb_439_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_439_bht_T_20 = _btb_439_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_21 = _btb_439_bht_T_16 ? 2'h0 : _btb_439_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_22 = _btb_439_bht_T_13 ? 2'h0 : _btb_439_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_23 = _btb_439_bht_T_10 ? 2'h0 : _btb_439_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_24 = _btb_439_bht_T_7 ? 2'h3 : _btb_439_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_25 = _btb_439_bht_T_5 ? 2'h3 : _btb_439_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_26 = _btb_439_bht_T_3 ? 2'h3 : _btb_439_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_439_bht_T_27 = _btb_439_bht_T_1 ? 2'h1 : _btb_439_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10462 = btb_439_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7095; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10464 = btb_439_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_439_bht_T_27 : _GEN_8631; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_440_bht_T = btb_440_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_440_bht_T_1 = io_i_branch_resolve_pack_taken & btb_440_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_440_bht_T_2 = btb_440_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_440_bht_T_3 = io_i_branch_resolve_pack_taken & btb_440_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_440_bht_T_4 = btb_440_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_440_bht_T_5 = io_i_branch_resolve_pack_taken & btb_440_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_440_bht_T_6 = btb_440_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_440_bht_T_7 = io_i_branch_resolve_pack_taken & btb_440_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_440_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_440_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_440_bht_T_13 = _btb_0_bht_T_8 & _btb_440_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_440_bht_T_16 = _btb_0_bht_T_8 & _btb_440_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_440_bht_T_19 = _btb_0_bht_T_8 & _btb_440_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_440_bht_T_20 = _btb_440_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_21 = _btb_440_bht_T_16 ? 2'h0 : _btb_440_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_22 = _btb_440_bht_T_13 ? 2'h0 : _btb_440_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_23 = _btb_440_bht_T_10 ? 2'h0 : _btb_440_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_24 = _btb_440_bht_T_7 ? 2'h3 : _btb_440_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_25 = _btb_440_bht_T_5 ? 2'h3 : _btb_440_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_26 = _btb_440_bht_T_3 ? 2'h3 : _btb_440_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_440_bht_T_27 = _btb_440_bht_T_1 ? 2'h1 : _btb_440_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10466 = btb_440_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7096; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10468 = btb_440_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_440_bht_T_27 : _GEN_8632; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_441_bht_T = btb_441_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_441_bht_T_1 = io_i_branch_resolve_pack_taken & btb_441_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_441_bht_T_2 = btb_441_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_441_bht_T_3 = io_i_branch_resolve_pack_taken & btb_441_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_441_bht_T_4 = btb_441_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_441_bht_T_5 = io_i_branch_resolve_pack_taken & btb_441_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_441_bht_T_6 = btb_441_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_441_bht_T_7 = io_i_branch_resolve_pack_taken & btb_441_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_441_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_441_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_441_bht_T_13 = _btb_0_bht_T_8 & _btb_441_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_441_bht_T_16 = _btb_0_bht_T_8 & _btb_441_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_441_bht_T_19 = _btb_0_bht_T_8 & _btb_441_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_441_bht_T_20 = _btb_441_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_21 = _btb_441_bht_T_16 ? 2'h0 : _btb_441_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_22 = _btb_441_bht_T_13 ? 2'h0 : _btb_441_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_23 = _btb_441_bht_T_10 ? 2'h0 : _btb_441_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_24 = _btb_441_bht_T_7 ? 2'h3 : _btb_441_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_25 = _btb_441_bht_T_5 ? 2'h3 : _btb_441_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_26 = _btb_441_bht_T_3 ? 2'h3 : _btb_441_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_441_bht_T_27 = _btb_441_bht_T_1 ? 2'h1 : _btb_441_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10470 = btb_441_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7097; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10472 = btb_441_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_441_bht_T_27 : _GEN_8633; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_442_bht_T = btb_442_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_442_bht_T_1 = io_i_branch_resolve_pack_taken & btb_442_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_442_bht_T_2 = btb_442_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_442_bht_T_3 = io_i_branch_resolve_pack_taken & btb_442_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_442_bht_T_4 = btb_442_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_442_bht_T_5 = io_i_branch_resolve_pack_taken & btb_442_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_442_bht_T_6 = btb_442_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_442_bht_T_7 = io_i_branch_resolve_pack_taken & btb_442_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_442_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_442_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_442_bht_T_13 = _btb_0_bht_T_8 & _btb_442_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_442_bht_T_16 = _btb_0_bht_T_8 & _btb_442_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_442_bht_T_19 = _btb_0_bht_T_8 & _btb_442_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_442_bht_T_20 = _btb_442_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_21 = _btb_442_bht_T_16 ? 2'h0 : _btb_442_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_22 = _btb_442_bht_T_13 ? 2'h0 : _btb_442_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_23 = _btb_442_bht_T_10 ? 2'h0 : _btb_442_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_24 = _btb_442_bht_T_7 ? 2'h3 : _btb_442_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_25 = _btb_442_bht_T_5 ? 2'h3 : _btb_442_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_26 = _btb_442_bht_T_3 ? 2'h3 : _btb_442_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_442_bht_T_27 = _btb_442_bht_T_1 ? 2'h1 : _btb_442_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10474 = btb_442_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7098; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10476 = btb_442_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_442_bht_T_27 : _GEN_8634; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_443_bht_T = btb_443_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_443_bht_T_1 = io_i_branch_resolve_pack_taken & btb_443_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_443_bht_T_2 = btb_443_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_443_bht_T_3 = io_i_branch_resolve_pack_taken & btb_443_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_443_bht_T_4 = btb_443_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_443_bht_T_5 = io_i_branch_resolve_pack_taken & btb_443_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_443_bht_T_6 = btb_443_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_443_bht_T_7 = io_i_branch_resolve_pack_taken & btb_443_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_443_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_443_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_443_bht_T_13 = _btb_0_bht_T_8 & _btb_443_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_443_bht_T_16 = _btb_0_bht_T_8 & _btb_443_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_443_bht_T_19 = _btb_0_bht_T_8 & _btb_443_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_443_bht_T_20 = _btb_443_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_21 = _btb_443_bht_T_16 ? 2'h0 : _btb_443_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_22 = _btb_443_bht_T_13 ? 2'h0 : _btb_443_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_23 = _btb_443_bht_T_10 ? 2'h0 : _btb_443_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_24 = _btb_443_bht_T_7 ? 2'h3 : _btb_443_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_25 = _btb_443_bht_T_5 ? 2'h3 : _btb_443_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_26 = _btb_443_bht_T_3 ? 2'h3 : _btb_443_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_443_bht_T_27 = _btb_443_bht_T_1 ? 2'h1 : _btb_443_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10478 = btb_443_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7099; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10480 = btb_443_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_443_bht_T_27 : _GEN_8635; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_444_bht_T = btb_444_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_444_bht_T_1 = io_i_branch_resolve_pack_taken & btb_444_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_444_bht_T_2 = btb_444_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_444_bht_T_3 = io_i_branch_resolve_pack_taken & btb_444_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_444_bht_T_4 = btb_444_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_444_bht_T_5 = io_i_branch_resolve_pack_taken & btb_444_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_444_bht_T_6 = btb_444_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_444_bht_T_7 = io_i_branch_resolve_pack_taken & btb_444_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_444_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_444_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_444_bht_T_13 = _btb_0_bht_T_8 & _btb_444_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_444_bht_T_16 = _btb_0_bht_T_8 & _btb_444_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_444_bht_T_19 = _btb_0_bht_T_8 & _btb_444_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_444_bht_T_20 = _btb_444_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_21 = _btb_444_bht_T_16 ? 2'h0 : _btb_444_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_22 = _btb_444_bht_T_13 ? 2'h0 : _btb_444_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_23 = _btb_444_bht_T_10 ? 2'h0 : _btb_444_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_24 = _btb_444_bht_T_7 ? 2'h3 : _btb_444_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_25 = _btb_444_bht_T_5 ? 2'h3 : _btb_444_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_26 = _btb_444_bht_T_3 ? 2'h3 : _btb_444_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_444_bht_T_27 = _btb_444_bht_T_1 ? 2'h1 : _btb_444_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10482 = btb_444_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7100; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10484 = btb_444_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_444_bht_T_27 : _GEN_8636; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_445_bht_T = btb_445_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_445_bht_T_1 = io_i_branch_resolve_pack_taken & btb_445_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_445_bht_T_2 = btb_445_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_445_bht_T_3 = io_i_branch_resolve_pack_taken & btb_445_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_445_bht_T_4 = btb_445_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_445_bht_T_5 = io_i_branch_resolve_pack_taken & btb_445_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_445_bht_T_6 = btb_445_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_445_bht_T_7 = io_i_branch_resolve_pack_taken & btb_445_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_445_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_445_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_445_bht_T_13 = _btb_0_bht_T_8 & _btb_445_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_445_bht_T_16 = _btb_0_bht_T_8 & _btb_445_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_445_bht_T_19 = _btb_0_bht_T_8 & _btb_445_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_445_bht_T_20 = _btb_445_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_21 = _btb_445_bht_T_16 ? 2'h0 : _btb_445_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_22 = _btb_445_bht_T_13 ? 2'h0 : _btb_445_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_23 = _btb_445_bht_T_10 ? 2'h0 : _btb_445_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_24 = _btb_445_bht_T_7 ? 2'h3 : _btb_445_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_25 = _btb_445_bht_T_5 ? 2'h3 : _btb_445_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_26 = _btb_445_bht_T_3 ? 2'h3 : _btb_445_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_445_bht_T_27 = _btb_445_bht_T_1 ? 2'h1 : _btb_445_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10486 = btb_445_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7101; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10488 = btb_445_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_445_bht_T_27 : _GEN_8637; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_446_bht_T = btb_446_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_446_bht_T_1 = io_i_branch_resolve_pack_taken & btb_446_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_446_bht_T_2 = btb_446_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_446_bht_T_3 = io_i_branch_resolve_pack_taken & btb_446_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_446_bht_T_4 = btb_446_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_446_bht_T_5 = io_i_branch_resolve_pack_taken & btb_446_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_446_bht_T_6 = btb_446_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_446_bht_T_7 = io_i_branch_resolve_pack_taken & btb_446_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_446_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_446_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_446_bht_T_13 = _btb_0_bht_T_8 & _btb_446_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_446_bht_T_16 = _btb_0_bht_T_8 & _btb_446_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_446_bht_T_19 = _btb_0_bht_T_8 & _btb_446_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_446_bht_T_20 = _btb_446_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_21 = _btb_446_bht_T_16 ? 2'h0 : _btb_446_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_22 = _btb_446_bht_T_13 ? 2'h0 : _btb_446_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_23 = _btb_446_bht_T_10 ? 2'h0 : _btb_446_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_24 = _btb_446_bht_T_7 ? 2'h3 : _btb_446_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_25 = _btb_446_bht_T_5 ? 2'h3 : _btb_446_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_26 = _btb_446_bht_T_3 ? 2'h3 : _btb_446_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_446_bht_T_27 = _btb_446_bht_T_1 ? 2'h1 : _btb_446_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10490 = btb_446_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7102; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10492 = btb_446_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_446_bht_T_27 : _GEN_8638; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_447_bht_T = btb_447_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_447_bht_T_1 = io_i_branch_resolve_pack_taken & btb_447_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_447_bht_T_2 = btb_447_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_447_bht_T_3 = io_i_branch_resolve_pack_taken & btb_447_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_447_bht_T_4 = btb_447_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_447_bht_T_5 = io_i_branch_resolve_pack_taken & btb_447_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_447_bht_T_6 = btb_447_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_447_bht_T_7 = io_i_branch_resolve_pack_taken & btb_447_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_447_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_447_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_447_bht_T_13 = _btb_0_bht_T_8 & _btb_447_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_447_bht_T_16 = _btb_0_bht_T_8 & _btb_447_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_447_bht_T_19 = _btb_0_bht_T_8 & _btb_447_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_447_bht_T_20 = _btb_447_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_21 = _btb_447_bht_T_16 ? 2'h0 : _btb_447_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_22 = _btb_447_bht_T_13 ? 2'h0 : _btb_447_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_23 = _btb_447_bht_T_10 ? 2'h0 : _btb_447_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_24 = _btb_447_bht_T_7 ? 2'h3 : _btb_447_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_25 = _btb_447_bht_T_5 ? 2'h3 : _btb_447_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_26 = _btb_447_bht_T_3 ? 2'h3 : _btb_447_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_447_bht_T_27 = _btb_447_bht_T_1 ? 2'h1 : _btb_447_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10494 = btb_447_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7103; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10496 = btb_447_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_447_bht_T_27 : _GEN_8639; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_448_bht_T = btb_448_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_448_bht_T_1 = io_i_branch_resolve_pack_taken & btb_448_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_448_bht_T_2 = btb_448_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_448_bht_T_3 = io_i_branch_resolve_pack_taken & btb_448_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_448_bht_T_4 = btb_448_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_448_bht_T_5 = io_i_branch_resolve_pack_taken & btb_448_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_448_bht_T_6 = btb_448_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_448_bht_T_7 = io_i_branch_resolve_pack_taken & btb_448_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_448_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_448_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_448_bht_T_13 = _btb_0_bht_T_8 & _btb_448_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_448_bht_T_16 = _btb_0_bht_T_8 & _btb_448_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_448_bht_T_19 = _btb_0_bht_T_8 & _btb_448_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_448_bht_T_20 = _btb_448_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_21 = _btb_448_bht_T_16 ? 2'h0 : _btb_448_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_22 = _btb_448_bht_T_13 ? 2'h0 : _btb_448_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_23 = _btb_448_bht_T_10 ? 2'h0 : _btb_448_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_24 = _btb_448_bht_T_7 ? 2'h3 : _btb_448_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_25 = _btb_448_bht_T_5 ? 2'h3 : _btb_448_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_26 = _btb_448_bht_T_3 ? 2'h3 : _btb_448_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_448_bht_T_27 = _btb_448_bht_T_1 ? 2'h1 : _btb_448_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10498 = btb_448_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7104; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10500 = btb_448_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_448_bht_T_27 : _GEN_8640; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_449_bht_T = btb_449_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_449_bht_T_1 = io_i_branch_resolve_pack_taken & btb_449_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_449_bht_T_2 = btb_449_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_449_bht_T_3 = io_i_branch_resolve_pack_taken & btb_449_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_449_bht_T_4 = btb_449_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_449_bht_T_5 = io_i_branch_resolve_pack_taken & btb_449_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_449_bht_T_6 = btb_449_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_449_bht_T_7 = io_i_branch_resolve_pack_taken & btb_449_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_449_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_449_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_449_bht_T_13 = _btb_0_bht_T_8 & _btb_449_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_449_bht_T_16 = _btb_0_bht_T_8 & _btb_449_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_449_bht_T_19 = _btb_0_bht_T_8 & _btb_449_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_449_bht_T_20 = _btb_449_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_21 = _btb_449_bht_T_16 ? 2'h0 : _btb_449_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_22 = _btb_449_bht_T_13 ? 2'h0 : _btb_449_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_23 = _btb_449_bht_T_10 ? 2'h0 : _btb_449_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_24 = _btb_449_bht_T_7 ? 2'h3 : _btb_449_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_25 = _btb_449_bht_T_5 ? 2'h3 : _btb_449_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_26 = _btb_449_bht_T_3 ? 2'h3 : _btb_449_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_449_bht_T_27 = _btb_449_bht_T_1 ? 2'h1 : _btb_449_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10501 = btb_449_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_448_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_447_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_446_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_445_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_444_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_443_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_442_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_441_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_440_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_439_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_438_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_437_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_436_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_435_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10441)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10502 = btb_449_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7105; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10504 = btb_449_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_449_bht_T_27 : _GEN_8641; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_450_bht_T = btb_450_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_450_bht_T_1 = io_i_branch_resolve_pack_taken & btb_450_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_450_bht_T_2 = btb_450_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_450_bht_T_3 = io_i_branch_resolve_pack_taken & btb_450_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_450_bht_T_4 = btb_450_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_450_bht_T_5 = io_i_branch_resolve_pack_taken & btb_450_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_450_bht_T_6 = btb_450_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_450_bht_T_7 = io_i_branch_resolve_pack_taken & btb_450_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_450_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_450_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_450_bht_T_13 = _btb_0_bht_T_8 & _btb_450_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_450_bht_T_16 = _btb_0_bht_T_8 & _btb_450_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_450_bht_T_19 = _btb_0_bht_T_8 & _btb_450_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_450_bht_T_20 = _btb_450_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_21 = _btb_450_bht_T_16 ? 2'h0 : _btb_450_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_22 = _btb_450_bht_T_13 ? 2'h0 : _btb_450_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_23 = _btb_450_bht_T_10 ? 2'h0 : _btb_450_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_24 = _btb_450_bht_T_7 ? 2'h3 : _btb_450_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_25 = _btb_450_bht_T_5 ? 2'h3 : _btb_450_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_26 = _btb_450_bht_T_3 ? 2'h3 : _btb_450_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_450_bht_T_27 = _btb_450_bht_T_1 ? 2'h1 : _btb_450_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10506 = btb_450_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7106; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10508 = btb_450_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_450_bht_T_27 : _GEN_8642; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_451_bht_T = btb_451_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_451_bht_T_1 = io_i_branch_resolve_pack_taken & btb_451_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_451_bht_T_2 = btb_451_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_451_bht_T_3 = io_i_branch_resolve_pack_taken & btb_451_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_451_bht_T_4 = btb_451_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_451_bht_T_5 = io_i_branch_resolve_pack_taken & btb_451_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_451_bht_T_6 = btb_451_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_451_bht_T_7 = io_i_branch_resolve_pack_taken & btb_451_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_451_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_451_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_451_bht_T_13 = _btb_0_bht_T_8 & _btb_451_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_451_bht_T_16 = _btb_0_bht_T_8 & _btb_451_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_451_bht_T_19 = _btb_0_bht_T_8 & _btb_451_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_451_bht_T_20 = _btb_451_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_21 = _btb_451_bht_T_16 ? 2'h0 : _btb_451_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_22 = _btb_451_bht_T_13 ? 2'h0 : _btb_451_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_23 = _btb_451_bht_T_10 ? 2'h0 : _btb_451_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_24 = _btb_451_bht_T_7 ? 2'h3 : _btb_451_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_25 = _btb_451_bht_T_5 ? 2'h3 : _btb_451_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_26 = _btb_451_bht_T_3 ? 2'h3 : _btb_451_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_451_bht_T_27 = _btb_451_bht_T_1 ? 2'h1 : _btb_451_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10510 = btb_451_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7107; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10512 = btb_451_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_451_bht_T_27 : _GEN_8643; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_452_bht_T = btb_452_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_452_bht_T_1 = io_i_branch_resolve_pack_taken & btb_452_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_452_bht_T_2 = btb_452_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_452_bht_T_3 = io_i_branch_resolve_pack_taken & btb_452_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_452_bht_T_4 = btb_452_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_452_bht_T_5 = io_i_branch_resolve_pack_taken & btb_452_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_452_bht_T_6 = btb_452_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_452_bht_T_7 = io_i_branch_resolve_pack_taken & btb_452_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_452_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_452_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_452_bht_T_13 = _btb_0_bht_T_8 & _btb_452_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_452_bht_T_16 = _btb_0_bht_T_8 & _btb_452_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_452_bht_T_19 = _btb_0_bht_T_8 & _btb_452_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_452_bht_T_20 = _btb_452_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_21 = _btb_452_bht_T_16 ? 2'h0 : _btb_452_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_22 = _btb_452_bht_T_13 ? 2'h0 : _btb_452_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_23 = _btb_452_bht_T_10 ? 2'h0 : _btb_452_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_24 = _btb_452_bht_T_7 ? 2'h3 : _btb_452_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_25 = _btb_452_bht_T_5 ? 2'h3 : _btb_452_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_26 = _btb_452_bht_T_3 ? 2'h3 : _btb_452_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_452_bht_T_27 = _btb_452_bht_T_1 ? 2'h1 : _btb_452_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10514 = btb_452_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7108; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10516 = btb_452_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_452_bht_T_27 : _GEN_8644; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_453_bht_T = btb_453_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_453_bht_T_1 = io_i_branch_resolve_pack_taken & btb_453_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_453_bht_T_2 = btb_453_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_453_bht_T_3 = io_i_branch_resolve_pack_taken & btb_453_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_453_bht_T_4 = btb_453_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_453_bht_T_5 = io_i_branch_resolve_pack_taken & btb_453_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_453_bht_T_6 = btb_453_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_453_bht_T_7 = io_i_branch_resolve_pack_taken & btb_453_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_453_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_453_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_453_bht_T_13 = _btb_0_bht_T_8 & _btb_453_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_453_bht_T_16 = _btb_0_bht_T_8 & _btb_453_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_453_bht_T_19 = _btb_0_bht_T_8 & _btb_453_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_453_bht_T_20 = _btb_453_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_21 = _btb_453_bht_T_16 ? 2'h0 : _btb_453_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_22 = _btb_453_bht_T_13 ? 2'h0 : _btb_453_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_23 = _btb_453_bht_T_10 ? 2'h0 : _btb_453_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_24 = _btb_453_bht_T_7 ? 2'h3 : _btb_453_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_25 = _btb_453_bht_T_5 ? 2'h3 : _btb_453_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_26 = _btb_453_bht_T_3 ? 2'h3 : _btb_453_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_453_bht_T_27 = _btb_453_bht_T_1 ? 2'h1 : _btb_453_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10518 = btb_453_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7109; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10520 = btb_453_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_453_bht_T_27 : _GEN_8645; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_454_bht_T = btb_454_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_454_bht_T_1 = io_i_branch_resolve_pack_taken & btb_454_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_454_bht_T_2 = btb_454_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_454_bht_T_3 = io_i_branch_resolve_pack_taken & btb_454_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_454_bht_T_4 = btb_454_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_454_bht_T_5 = io_i_branch_resolve_pack_taken & btb_454_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_454_bht_T_6 = btb_454_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_454_bht_T_7 = io_i_branch_resolve_pack_taken & btb_454_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_454_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_454_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_454_bht_T_13 = _btb_0_bht_T_8 & _btb_454_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_454_bht_T_16 = _btb_0_bht_T_8 & _btb_454_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_454_bht_T_19 = _btb_0_bht_T_8 & _btb_454_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_454_bht_T_20 = _btb_454_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_21 = _btb_454_bht_T_16 ? 2'h0 : _btb_454_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_22 = _btb_454_bht_T_13 ? 2'h0 : _btb_454_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_23 = _btb_454_bht_T_10 ? 2'h0 : _btb_454_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_24 = _btb_454_bht_T_7 ? 2'h3 : _btb_454_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_25 = _btb_454_bht_T_5 ? 2'h3 : _btb_454_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_26 = _btb_454_bht_T_3 ? 2'h3 : _btb_454_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_454_bht_T_27 = _btb_454_bht_T_1 ? 2'h1 : _btb_454_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10522 = btb_454_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7110; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10524 = btb_454_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_454_bht_T_27 : _GEN_8646; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_455_bht_T = btb_455_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_455_bht_T_1 = io_i_branch_resolve_pack_taken & btb_455_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_455_bht_T_2 = btb_455_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_455_bht_T_3 = io_i_branch_resolve_pack_taken & btb_455_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_455_bht_T_4 = btb_455_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_455_bht_T_5 = io_i_branch_resolve_pack_taken & btb_455_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_455_bht_T_6 = btb_455_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_455_bht_T_7 = io_i_branch_resolve_pack_taken & btb_455_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_455_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_455_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_455_bht_T_13 = _btb_0_bht_T_8 & _btb_455_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_455_bht_T_16 = _btb_0_bht_T_8 & _btb_455_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_455_bht_T_19 = _btb_0_bht_T_8 & _btb_455_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_455_bht_T_20 = _btb_455_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_21 = _btb_455_bht_T_16 ? 2'h0 : _btb_455_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_22 = _btb_455_bht_T_13 ? 2'h0 : _btb_455_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_23 = _btb_455_bht_T_10 ? 2'h0 : _btb_455_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_24 = _btb_455_bht_T_7 ? 2'h3 : _btb_455_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_25 = _btb_455_bht_T_5 ? 2'h3 : _btb_455_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_26 = _btb_455_bht_T_3 ? 2'h3 : _btb_455_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_455_bht_T_27 = _btb_455_bht_T_1 ? 2'h1 : _btb_455_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10526 = btb_455_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7111; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10528 = btb_455_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_455_bht_T_27 : _GEN_8647; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_456_bht_T = btb_456_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_456_bht_T_1 = io_i_branch_resolve_pack_taken & btb_456_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_456_bht_T_2 = btb_456_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_456_bht_T_3 = io_i_branch_resolve_pack_taken & btb_456_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_456_bht_T_4 = btb_456_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_456_bht_T_5 = io_i_branch_resolve_pack_taken & btb_456_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_456_bht_T_6 = btb_456_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_456_bht_T_7 = io_i_branch_resolve_pack_taken & btb_456_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_456_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_456_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_456_bht_T_13 = _btb_0_bht_T_8 & _btb_456_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_456_bht_T_16 = _btb_0_bht_T_8 & _btb_456_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_456_bht_T_19 = _btb_0_bht_T_8 & _btb_456_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_456_bht_T_20 = _btb_456_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_21 = _btb_456_bht_T_16 ? 2'h0 : _btb_456_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_22 = _btb_456_bht_T_13 ? 2'h0 : _btb_456_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_23 = _btb_456_bht_T_10 ? 2'h0 : _btb_456_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_24 = _btb_456_bht_T_7 ? 2'h3 : _btb_456_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_25 = _btb_456_bht_T_5 ? 2'h3 : _btb_456_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_26 = _btb_456_bht_T_3 ? 2'h3 : _btb_456_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_456_bht_T_27 = _btb_456_bht_T_1 ? 2'h1 : _btb_456_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10530 = btb_456_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7112; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10532 = btb_456_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_456_bht_T_27 : _GEN_8648; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_457_bht_T = btb_457_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_457_bht_T_1 = io_i_branch_resolve_pack_taken & btb_457_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_457_bht_T_2 = btb_457_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_457_bht_T_3 = io_i_branch_resolve_pack_taken & btb_457_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_457_bht_T_4 = btb_457_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_457_bht_T_5 = io_i_branch_resolve_pack_taken & btb_457_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_457_bht_T_6 = btb_457_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_457_bht_T_7 = io_i_branch_resolve_pack_taken & btb_457_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_457_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_457_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_457_bht_T_13 = _btb_0_bht_T_8 & _btb_457_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_457_bht_T_16 = _btb_0_bht_T_8 & _btb_457_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_457_bht_T_19 = _btb_0_bht_T_8 & _btb_457_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_457_bht_T_20 = _btb_457_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_21 = _btb_457_bht_T_16 ? 2'h0 : _btb_457_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_22 = _btb_457_bht_T_13 ? 2'h0 : _btb_457_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_23 = _btb_457_bht_T_10 ? 2'h0 : _btb_457_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_24 = _btb_457_bht_T_7 ? 2'h3 : _btb_457_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_25 = _btb_457_bht_T_5 ? 2'h3 : _btb_457_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_26 = _btb_457_bht_T_3 ? 2'h3 : _btb_457_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_457_bht_T_27 = _btb_457_bht_T_1 ? 2'h1 : _btb_457_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10534 = btb_457_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7113; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10536 = btb_457_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_457_bht_T_27 : _GEN_8649; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_458_bht_T = btb_458_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_458_bht_T_1 = io_i_branch_resolve_pack_taken & btb_458_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_458_bht_T_2 = btb_458_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_458_bht_T_3 = io_i_branch_resolve_pack_taken & btb_458_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_458_bht_T_4 = btb_458_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_458_bht_T_5 = io_i_branch_resolve_pack_taken & btb_458_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_458_bht_T_6 = btb_458_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_458_bht_T_7 = io_i_branch_resolve_pack_taken & btb_458_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_458_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_458_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_458_bht_T_13 = _btb_0_bht_T_8 & _btb_458_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_458_bht_T_16 = _btb_0_bht_T_8 & _btb_458_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_458_bht_T_19 = _btb_0_bht_T_8 & _btb_458_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_458_bht_T_20 = _btb_458_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_21 = _btb_458_bht_T_16 ? 2'h0 : _btb_458_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_22 = _btb_458_bht_T_13 ? 2'h0 : _btb_458_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_23 = _btb_458_bht_T_10 ? 2'h0 : _btb_458_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_24 = _btb_458_bht_T_7 ? 2'h3 : _btb_458_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_25 = _btb_458_bht_T_5 ? 2'h3 : _btb_458_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_26 = _btb_458_bht_T_3 ? 2'h3 : _btb_458_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_458_bht_T_27 = _btb_458_bht_T_1 ? 2'h1 : _btb_458_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10538 = btb_458_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7114; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10540 = btb_458_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_458_bht_T_27 : _GEN_8650; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_459_bht_T = btb_459_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_459_bht_T_1 = io_i_branch_resolve_pack_taken & btb_459_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_459_bht_T_2 = btb_459_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_459_bht_T_3 = io_i_branch_resolve_pack_taken & btb_459_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_459_bht_T_4 = btb_459_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_459_bht_T_5 = io_i_branch_resolve_pack_taken & btb_459_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_459_bht_T_6 = btb_459_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_459_bht_T_7 = io_i_branch_resolve_pack_taken & btb_459_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_459_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_459_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_459_bht_T_13 = _btb_0_bht_T_8 & _btb_459_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_459_bht_T_16 = _btb_0_bht_T_8 & _btb_459_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_459_bht_T_19 = _btb_0_bht_T_8 & _btb_459_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_459_bht_T_20 = _btb_459_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_21 = _btb_459_bht_T_16 ? 2'h0 : _btb_459_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_22 = _btb_459_bht_T_13 ? 2'h0 : _btb_459_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_23 = _btb_459_bht_T_10 ? 2'h0 : _btb_459_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_24 = _btb_459_bht_T_7 ? 2'h3 : _btb_459_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_25 = _btb_459_bht_T_5 ? 2'h3 : _btb_459_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_26 = _btb_459_bht_T_3 ? 2'h3 : _btb_459_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_459_bht_T_27 = _btb_459_bht_T_1 ? 2'h1 : _btb_459_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10542 = btb_459_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7115; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10544 = btb_459_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_459_bht_T_27 : _GEN_8651; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_460_bht_T = btb_460_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_460_bht_T_1 = io_i_branch_resolve_pack_taken & btb_460_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_460_bht_T_2 = btb_460_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_460_bht_T_3 = io_i_branch_resolve_pack_taken & btb_460_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_460_bht_T_4 = btb_460_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_460_bht_T_5 = io_i_branch_resolve_pack_taken & btb_460_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_460_bht_T_6 = btb_460_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_460_bht_T_7 = io_i_branch_resolve_pack_taken & btb_460_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_460_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_460_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_460_bht_T_13 = _btb_0_bht_T_8 & _btb_460_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_460_bht_T_16 = _btb_0_bht_T_8 & _btb_460_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_460_bht_T_19 = _btb_0_bht_T_8 & _btb_460_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_460_bht_T_20 = _btb_460_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_21 = _btb_460_bht_T_16 ? 2'h0 : _btb_460_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_22 = _btb_460_bht_T_13 ? 2'h0 : _btb_460_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_23 = _btb_460_bht_T_10 ? 2'h0 : _btb_460_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_24 = _btb_460_bht_T_7 ? 2'h3 : _btb_460_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_25 = _btb_460_bht_T_5 ? 2'h3 : _btb_460_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_26 = _btb_460_bht_T_3 ? 2'h3 : _btb_460_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_460_bht_T_27 = _btb_460_bht_T_1 ? 2'h1 : _btb_460_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10546 = btb_460_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7116; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10548 = btb_460_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_460_bht_T_27 : _GEN_8652; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_461_bht_T = btb_461_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_461_bht_T_1 = io_i_branch_resolve_pack_taken & btb_461_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_461_bht_T_2 = btb_461_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_461_bht_T_3 = io_i_branch_resolve_pack_taken & btb_461_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_461_bht_T_4 = btb_461_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_461_bht_T_5 = io_i_branch_resolve_pack_taken & btb_461_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_461_bht_T_6 = btb_461_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_461_bht_T_7 = io_i_branch_resolve_pack_taken & btb_461_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_461_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_461_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_461_bht_T_13 = _btb_0_bht_T_8 & _btb_461_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_461_bht_T_16 = _btb_0_bht_T_8 & _btb_461_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_461_bht_T_19 = _btb_0_bht_T_8 & _btb_461_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_461_bht_T_20 = _btb_461_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_21 = _btb_461_bht_T_16 ? 2'h0 : _btb_461_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_22 = _btb_461_bht_T_13 ? 2'h0 : _btb_461_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_23 = _btb_461_bht_T_10 ? 2'h0 : _btb_461_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_24 = _btb_461_bht_T_7 ? 2'h3 : _btb_461_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_25 = _btb_461_bht_T_5 ? 2'h3 : _btb_461_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_26 = _btb_461_bht_T_3 ? 2'h3 : _btb_461_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_461_bht_T_27 = _btb_461_bht_T_1 ? 2'h1 : _btb_461_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10550 = btb_461_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7117; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10552 = btb_461_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_461_bht_T_27 : _GEN_8653; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_462_bht_T = btb_462_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_462_bht_T_1 = io_i_branch_resolve_pack_taken & btb_462_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_462_bht_T_2 = btb_462_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_462_bht_T_3 = io_i_branch_resolve_pack_taken & btb_462_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_462_bht_T_4 = btb_462_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_462_bht_T_5 = io_i_branch_resolve_pack_taken & btb_462_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_462_bht_T_6 = btb_462_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_462_bht_T_7 = io_i_branch_resolve_pack_taken & btb_462_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_462_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_462_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_462_bht_T_13 = _btb_0_bht_T_8 & _btb_462_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_462_bht_T_16 = _btb_0_bht_T_8 & _btb_462_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_462_bht_T_19 = _btb_0_bht_T_8 & _btb_462_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_462_bht_T_20 = _btb_462_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_21 = _btb_462_bht_T_16 ? 2'h0 : _btb_462_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_22 = _btb_462_bht_T_13 ? 2'h0 : _btb_462_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_23 = _btb_462_bht_T_10 ? 2'h0 : _btb_462_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_24 = _btb_462_bht_T_7 ? 2'h3 : _btb_462_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_25 = _btb_462_bht_T_5 ? 2'h3 : _btb_462_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_26 = _btb_462_bht_T_3 ? 2'h3 : _btb_462_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_462_bht_T_27 = _btb_462_bht_T_1 ? 2'h1 : _btb_462_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10554 = btb_462_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7118; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10556 = btb_462_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_462_bht_T_27 : _GEN_8654; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_463_bht_T = btb_463_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_463_bht_T_1 = io_i_branch_resolve_pack_taken & btb_463_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_463_bht_T_2 = btb_463_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_463_bht_T_3 = io_i_branch_resolve_pack_taken & btb_463_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_463_bht_T_4 = btb_463_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_463_bht_T_5 = io_i_branch_resolve_pack_taken & btb_463_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_463_bht_T_6 = btb_463_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_463_bht_T_7 = io_i_branch_resolve_pack_taken & btb_463_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_463_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_463_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_463_bht_T_13 = _btb_0_bht_T_8 & _btb_463_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_463_bht_T_16 = _btb_0_bht_T_8 & _btb_463_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_463_bht_T_19 = _btb_0_bht_T_8 & _btb_463_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_463_bht_T_20 = _btb_463_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_21 = _btb_463_bht_T_16 ? 2'h0 : _btb_463_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_22 = _btb_463_bht_T_13 ? 2'h0 : _btb_463_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_23 = _btb_463_bht_T_10 ? 2'h0 : _btb_463_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_24 = _btb_463_bht_T_7 ? 2'h3 : _btb_463_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_25 = _btb_463_bht_T_5 ? 2'h3 : _btb_463_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_26 = _btb_463_bht_T_3 ? 2'h3 : _btb_463_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_463_bht_T_27 = _btb_463_bht_T_1 ? 2'h1 : _btb_463_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10558 = btb_463_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7119; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10560 = btb_463_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_463_bht_T_27 : _GEN_8655; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_464_bht_T = btb_464_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_464_bht_T_1 = io_i_branch_resolve_pack_taken & btb_464_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_464_bht_T_2 = btb_464_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_464_bht_T_3 = io_i_branch_resolve_pack_taken & btb_464_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_464_bht_T_4 = btb_464_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_464_bht_T_5 = io_i_branch_resolve_pack_taken & btb_464_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_464_bht_T_6 = btb_464_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_464_bht_T_7 = io_i_branch_resolve_pack_taken & btb_464_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_464_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_464_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_464_bht_T_13 = _btb_0_bht_T_8 & _btb_464_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_464_bht_T_16 = _btb_0_bht_T_8 & _btb_464_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_464_bht_T_19 = _btb_0_bht_T_8 & _btb_464_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_464_bht_T_20 = _btb_464_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_21 = _btb_464_bht_T_16 ? 2'h0 : _btb_464_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_22 = _btb_464_bht_T_13 ? 2'h0 : _btb_464_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_23 = _btb_464_bht_T_10 ? 2'h0 : _btb_464_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_24 = _btb_464_bht_T_7 ? 2'h3 : _btb_464_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_25 = _btb_464_bht_T_5 ? 2'h3 : _btb_464_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_26 = _btb_464_bht_T_3 ? 2'h3 : _btb_464_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_464_bht_T_27 = _btb_464_bht_T_1 ? 2'h1 : _btb_464_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10561 = btb_464_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_463_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_462_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_461_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_460_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_459_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_458_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_457_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_456_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_455_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_454_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_453_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_452_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_451_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_450_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10501)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10562 = btb_464_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7120; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10564 = btb_464_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_464_bht_T_27 : _GEN_8656; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_465_bht_T = btb_465_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_465_bht_T_1 = io_i_branch_resolve_pack_taken & btb_465_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_465_bht_T_2 = btb_465_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_465_bht_T_3 = io_i_branch_resolve_pack_taken & btb_465_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_465_bht_T_4 = btb_465_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_465_bht_T_5 = io_i_branch_resolve_pack_taken & btb_465_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_465_bht_T_6 = btb_465_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_465_bht_T_7 = io_i_branch_resolve_pack_taken & btb_465_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_465_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_465_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_465_bht_T_13 = _btb_0_bht_T_8 & _btb_465_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_465_bht_T_16 = _btb_0_bht_T_8 & _btb_465_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_465_bht_T_19 = _btb_0_bht_T_8 & _btb_465_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_465_bht_T_20 = _btb_465_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_21 = _btb_465_bht_T_16 ? 2'h0 : _btb_465_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_22 = _btb_465_bht_T_13 ? 2'h0 : _btb_465_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_23 = _btb_465_bht_T_10 ? 2'h0 : _btb_465_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_24 = _btb_465_bht_T_7 ? 2'h3 : _btb_465_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_25 = _btb_465_bht_T_5 ? 2'h3 : _btb_465_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_26 = _btb_465_bht_T_3 ? 2'h3 : _btb_465_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_465_bht_T_27 = _btb_465_bht_T_1 ? 2'h1 : _btb_465_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10566 = btb_465_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7121; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10568 = btb_465_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_465_bht_T_27 : _GEN_8657; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_466_bht_T = btb_466_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_466_bht_T_1 = io_i_branch_resolve_pack_taken & btb_466_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_466_bht_T_2 = btb_466_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_466_bht_T_3 = io_i_branch_resolve_pack_taken & btb_466_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_466_bht_T_4 = btb_466_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_466_bht_T_5 = io_i_branch_resolve_pack_taken & btb_466_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_466_bht_T_6 = btb_466_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_466_bht_T_7 = io_i_branch_resolve_pack_taken & btb_466_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_466_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_466_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_466_bht_T_13 = _btb_0_bht_T_8 & _btb_466_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_466_bht_T_16 = _btb_0_bht_T_8 & _btb_466_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_466_bht_T_19 = _btb_0_bht_T_8 & _btb_466_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_466_bht_T_20 = _btb_466_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_21 = _btb_466_bht_T_16 ? 2'h0 : _btb_466_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_22 = _btb_466_bht_T_13 ? 2'h0 : _btb_466_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_23 = _btb_466_bht_T_10 ? 2'h0 : _btb_466_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_24 = _btb_466_bht_T_7 ? 2'h3 : _btb_466_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_25 = _btb_466_bht_T_5 ? 2'h3 : _btb_466_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_26 = _btb_466_bht_T_3 ? 2'h3 : _btb_466_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_466_bht_T_27 = _btb_466_bht_T_1 ? 2'h1 : _btb_466_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10570 = btb_466_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7122; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10572 = btb_466_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_466_bht_T_27 : _GEN_8658; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_467_bht_T = btb_467_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_467_bht_T_1 = io_i_branch_resolve_pack_taken & btb_467_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_467_bht_T_2 = btb_467_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_467_bht_T_3 = io_i_branch_resolve_pack_taken & btb_467_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_467_bht_T_4 = btb_467_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_467_bht_T_5 = io_i_branch_resolve_pack_taken & btb_467_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_467_bht_T_6 = btb_467_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_467_bht_T_7 = io_i_branch_resolve_pack_taken & btb_467_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_467_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_467_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_467_bht_T_13 = _btb_0_bht_T_8 & _btb_467_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_467_bht_T_16 = _btb_0_bht_T_8 & _btb_467_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_467_bht_T_19 = _btb_0_bht_T_8 & _btb_467_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_467_bht_T_20 = _btb_467_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_21 = _btb_467_bht_T_16 ? 2'h0 : _btb_467_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_22 = _btb_467_bht_T_13 ? 2'h0 : _btb_467_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_23 = _btb_467_bht_T_10 ? 2'h0 : _btb_467_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_24 = _btb_467_bht_T_7 ? 2'h3 : _btb_467_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_25 = _btb_467_bht_T_5 ? 2'h3 : _btb_467_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_26 = _btb_467_bht_T_3 ? 2'h3 : _btb_467_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_467_bht_T_27 = _btb_467_bht_T_1 ? 2'h1 : _btb_467_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10574 = btb_467_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7123; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10576 = btb_467_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_467_bht_T_27 : _GEN_8659; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_468_bht_T = btb_468_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_468_bht_T_1 = io_i_branch_resolve_pack_taken & btb_468_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_468_bht_T_2 = btb_468_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_468_bht_T_3 = io_i_branch_resolve_pack_taken & btb_468_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_468_bht_T_4 = btb_468_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_468_bht_T_5 = io_i_branch_resolve_pack_taken & btb_468_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_468_bht_T_6 = btb_468_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_468_bht_T_7 = io_i_branch_resolve_pack_taken & btb_468_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_468_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_468_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_468_bht_T_13 = _btb_0_bht_T_8 & _btb_468_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_468_bht_T_16 = _btb_0_bht_T_8 & _btb_468_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_468_bht_T_19 = _btb_0_bht_T_8 & _btb_468_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_468_bht_T_20 = _btb_468_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_21 = _btb_468_bht_T_16 ? 2'h0 : _btb_468_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_22 = _btb_468_bht_T_13 ? 2'h0 : _btb_468_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_23 = _btb_468_bht_T_10 ? 2'h0 : _btb_468_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_24 = _btb_468_bht_T_7 ? 2'h3 : _btb_468_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_25 = _btb_468_bht_T_5 ? 2'h3 : _btb_468_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_26 = _btb_468_bht_T_3 ? 2'h3 : _btb_468_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_468_bht_T_27 = _btb_468_bht_T_1 ? 2'h1 : _btb_468_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10578 = btb_468_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7124; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10580 = btb_468_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_468_bht_T_27 : _GEN_8660; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_469_bht_T = btb_469_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_469_bht_T_1 = io_i_branch_resolve_pack_taken & btb_469_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_469_bht_T_2 = btb_469_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_469_bht_T_3 = io_i_branch_resolve_pack_taken & btb_469_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_469_bht_T_4 = btb_469_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_469_bht_T_5 = io_i_branch_resolve_pack_taken & btb_469_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_469_bht_T_6 = btb_469_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_469_bht_T_7 = io_i_branch_resolve_pack_taken & btb_469_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_469_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_469_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_469_bht_T_13 = _btb_0_bht_T_8 & _btb_469_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_469_bht_T_16 = _btb_0_bht_T_8 & _btb_469_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_469_bht_T_19 = _btb_0_bht_T_8 & _btb_469_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_469_bht_T_20 = _btb_469_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_21 = _btb_469_bht_T_16 ? 2'h0 : _btb_469_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_22 = _btb_469_bht_T_13 ? 2'h0 : _btb_469_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_23 = _btb_469_bht_T_10 ? 2'h0 : _btb_469_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_24 = _btb_469_bht_T_7 ? 2'h3 : _btb_469_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_25 = _btb_469_bht_T_5 ? 2'h3 : _btb_469_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_26 = _btb_469_bht_T_3 ? 2'h3 : _btb_469_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_469_bht_T_27 = _btb_469_bht_T_1 ? 2'h1 : _btb_469_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10582 = btb_469_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7125; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10584 = btb_469_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_469_bht_T_27 : _GEN_8661; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_470_bht_T = btb_470_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_470_bht_T_1 = io_i_branch_resolve_pack_taken & btb_470_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_470_bht_T_2 = btb_470_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_470_bht_T_3 = io_i_branch_resolve_pack_taken & btb_470_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_470_bht_T_4 = btb_470_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_470_bht_T_5 = io_i_branch_resolve_pack_taken & btb_470_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_470_bht_T_6 = btb_470_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_470_bht_T_7 = io_i_branch_resolve_pack_taken & btb_470_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_470_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_470_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_470_bht_T_13 = _btb_0_bht_T_8 & _btb_470_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_470_bht_T_16 = _btb_0_bht_T_8 & _btb_470_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_470_bht_T_19 = _btb_0_bht_T_8 & _btb_470_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_470_bht_T_20 = _btb_470_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_21 = _btb_470_bht_T_16 ? 2'h0 : _btb_470_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_22 = _btb_470_bht_T_13 ? 2'h0 : _btb_470_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_23 = _btb_470_bht_T_10 ? 2'h0 : _btb_470_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_24 = _btb_470_bht_T_7 ? 2'h3 : _btb_470_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_25 = _btb_470_bht_T_5 ? 2'h3 : _btb_470_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_26 = _btb_470_bht_T_3 ? 2'h3 : _btb_470_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_470_bht_T_27 = _btb_470_bht_T_1 ? 2'h1 : _btb_470_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10586 = btb_470_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7126; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10588 = btb_470_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_470_bht_T_27 : _GEN_8662; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_471_bht_T = btb_471_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_471_bht_T_1 = io_i_branch_resolve_pack_taken & btb_471_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_471_bht_T_2 = btb_471_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_471_bht_T_3 = io_i_branch_resolve_pack_taken & btb_471_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_471_bht_T_4 = btb_471_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_471_bht_T_5 = io_i_branch_resolve_pack_taken & btb_471_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_471_bht_T_6 = btb_471_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_471_bht_T_7 = io_i_branch_resolve_pack_taken & btb_471_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_471_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_471_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_471_bht_T_13 = _btb_0_bht_T_8 & _btb_471_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_471_bht_T_16 = _btb_0_bht_T_8 & _btb_471_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_471_bht_T_19 = _btb_0_bht_T_8 & _btb_471_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_471_bht_T_20 = _btb_471_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_21 = _btb_471_bht_T_16 ? 2'h0 : _btb_471_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_22 = _btb_471_bht_T_13 ? 2'h0 : _btb_471_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_23 = _btb_471_bht_T_10 ? 2'h0 : _btb_471_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_24 = _btb_471_bht_T_7 ? 2'h3 : _btb_471_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_25 = _btb_471_bht_T_5 ? 2'h3 : _btb_471_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_26 = _btb_471_bht_T_3 ? 2'h3 : _btb_471_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_471_bht_T_27 = _btb_471_bht_T_1 ? 2'h1 : _btb_471_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10590 = btb_471_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7127; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10592 = btb_471_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_471_bht_T_27 : _GEN_8663; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_472_bht_T = btb_472_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_472_bht_T_1 = io_i_branch_resolve_pack_taken & btb_472_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_472_bht_T_2 = btb_472_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_472_bht_T_3 = io_i_branch_resolve_pack_taken & btb_472_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_472_bht_T_4 = btb_472_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_472_bht_T_5 = io_i_branch_resolve_pack_taken & btb_472_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_472_bht_T_6 = btb_472_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_472_bht_T_7 = io_i_branch_resolve_pack_taken & btb_472_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_472_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_472_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_472_bht_T_13 = _btb_0_bht_T_8 & _btb_472_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_472_bht_T_16 = _btb_0_bht_T_8 & _btb_472_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_472_bht_T_19 = _btb_0_bht_T_8 & _btb_472_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_472_bht_T_20 = _btb_472_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_21 = _btb_472_bht_T_16 ? 2'h0 : _btb_472_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_22 = _btb_472_bht_T_13 ? 2'h0 : _btb_472_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_23 = _btb_472_bht_T_10 ? 2'h0 : _btb_472_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_24 = _btb_472_bht_T_7 ? 2'h3 : _btb_472_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_25 = _btb_472_bht_T_5 ? 2'h3 : _btb_472_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_26 = _btb_472_bht_T_3 ? 2'h3 : _btb_472_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_472_bht_T_27 = _btb_472_bht_T_1 ? 2'h1 : _btb_472_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10594 = btb_472_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7128; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10596 = btb_472_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_472_bht_T_27 : _GEN_8664; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_473_bht_T = btb_473_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_473_bht_T_1 = io_i_branch_resolve_pack_taken & btb_473_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_473_bht_T_2 = btb_473_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_473_bht_T_3 = io_i_branch_resolve_pack_taken & btb_473_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_473_bht_T_4 = btb_473_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_473_bht_T_5 = io_i_branch_resolve_pack_taken & btb_473_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_473_bht_T_6 = btb_473_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_473_bht_T_7 = io_i_branch_resolve_pack_taken & btb_473_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_473_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_473_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_473_bht_T_13 = _btb_0_bht_T_8 & _btb_473_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_473_bht_T_16 = _btb_0_bht_T_8 & _btb_473_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_473_bht_T_19 = _btb_0_bht_T_8 & _btb_473_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_473_bht_T_20 = _btb_473_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_21 = _btb_473_bht_T_16 ? 2'h0 : _btb_473_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_22 = _btb_473_bht_T_13 ? 2'h0 : _btb_473_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_23 = _btb_473_bht_T_10 ? 2'h0 : _btb_473_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_24 = _btb_473_bht_T_7 ? 2'h3 : _btb_473_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_25 = _btb_473_bht_T_5 ? 2'h3 : _btb_473_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_26 = _btb_473_bht_T_3 ? 2'h3 : _btb_473_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_473_bht_T_27 = _btb_473_bht_T_1 ? 2'h1 : _btb_473_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10598 = btb_473_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7129; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10600 = btb_473_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_473_bht_T_27 : _GEN_8665; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_474_bht_T = btb_474_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_474_bht_T_1 = io_i_branch_resolve_pack_taken & btb_474_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_474_bht_T_2 = btb_474_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_474_bht_T_3 = io_i_branch_resolve_pack_taken & btb_474_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_474_bht_T_4 = btb_474_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_474_bht_T_5 = io_i_branch_resolve_pack_taken & btb_474_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_474_bht_T_6 = btb_474_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_474_bht_T_7 = io_i_branch_resolve_pack_taken & btb_474_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_474_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_474_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_474_bht_T_13 = _btb_0_bht_T_8 & _btb_474_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_474_bht_T_16 = _btb_0_bht_T_8 & _btb_474_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_474_bht_T_19 = _btb_0_bht_T_8 & _btb_474_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_474_bht_T_20 = _btb_474_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_21 = _btb_474_bht_T_16 ? 2'h0 : _btb_474_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_22 = _btb_474_bht_T_13 ? 2'h0 : _btb_474_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_23 = _btb_474_bht_T_10 ? 2'h0 : _btb_474_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_24 = _btb_474_bht_T_7 ? 2'h3 : _btb_474_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_25 = _btb_474_bht_T_5 ? 2'h3 : _btb_474_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_26 = _btb_474_bht_T_3 ? 2'h3 : _btb_474_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_474_bht_T_27 = _btb_474_bht_T_1 ? 2'h1 : _btb_474_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10602 = btb_474_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7130; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10604 = btb_474_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_474_bht_T_27 : _GEN_8666; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_475_bht_T = btb_475_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_475_bht_T_1 = io_i_branch_resolve_pack_taken & btb_475_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_475_bht_T_2 = btb_475_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_475_bht_T_3 = io_i_branch_resolve_pack_taken & btb_475_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_475_bht_T_4 = btb_475_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_475_bht_T_5 = io_i_branch_resolve_pack_taken & btb_475_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_475_bht_T_6 = btb_475_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_475_bht_T_7 = io_i_branch_resolve_pack_taken & btb_475_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_475_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_475_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_475_bht_T_13 = _btb_0_bht_T_8 & _btb_475_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_475_bht_T_16 = _btb_0_bht_T_8 & _btb_475_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_475_bht_T_19 = _btb_0_bht_T_8 & _btb_475_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_475_bht_T_20 = _btb_475_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_21 = _btb_475_bht_T_16 ? 2'h0 : _btb_475_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_22 = _btb_475_bht_T_13 ? 2'h0 : _btb_475_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_23 = _btb_475_bht_T_10 ? 2'h0 : _btb_475_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_24 = _btb_475_bht_T_7 ? 2'h3 : _btb_475_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_25 = _btb_475_bht_T_5 ? 2'h3 : _btb_475_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_26 = _btb_475_bht_T_3 ? 2'h3 : _btb_475_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_475_bht_T_27 = _btb_475_bht_T_1 ? 2'h1 : _btb_475_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10606 = btb_475_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7131; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10608 = btb_475_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_475_bht_T_27 : _GEN_8667; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_476_bht_T = btb_476_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_476_bht_T_1 = io_i_branch_resolve_pack_taken & btb_476_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_476_bht_T_2 = btb_476_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_476_bht_T_3 = io_i_branch_resolve_pack_taken & btb_476_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_476_bht_T_4 = btb_476_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_476_bht_T_5 = io_i_branch_resolve_pack_taken & btb_476_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_476_bht_T_6 = btb_476_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_476_bht_T_7 = io_i_branch_resolve_pack_taken & btb_476_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_476_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_476_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_476_bht_T_13 = _btb_0_bht_T_8 & _btb_476_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_476_bht_T_16 = _btb_0_bht_T_8 & _btb_476_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_476_bht_T_19 = _btb_0_bht_T_8 & _btb_476_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_476_bht_T_20 = _btb_476_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_21 = _btb_476_bht_T_16 ? 2'h0 : _btb_476_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_22 = _btb_476_bht_T_13 ? 2'h0 : _btb_476_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_23 = _btb_476_bht_T_10 ? 2'h0 : _btb_476_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_24 = _btb_476_bht_T_7 ? 2'h3 : _btb_476_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_25 = _btb_476_bht_T_5 ? 2'h3 : _btb_476_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_26 = _btb_476_bht_T_3 ? 2'h3 : _btb_476_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_476_bht_T_27 = _btb_476_bht_T_1 ? 2'h1 : _btb_476_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10610 = btb_476_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7132; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10612 = btb_476_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_476_bht_T_27 : _GEN_8668; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_477_bht_T = btb_477_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_477_bht_T_1 = io_i_branch_resolve_pack_taken & btb_477_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_477_bht_T_2 = btb_477_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_477_bht_T_3 = io_i_branch_resolve_pack_taken & btb_477_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_477_bht_T_4 = btb_477_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_477_bht_T_5 = io_i_branch_resolve_pack_taken & btb_477_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_477_bht_T_6 = btb_477_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_477_bht_T_7 = io_i_branch_resolve_pack_taken & btb_477_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_477_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_477_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_477_bht_T_13 = _btb_0_bht_T_8 & _btb_477_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_477_bht_T_16 = _btb_0_bht_T_8 & _btb_477_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_477_bht_T_19 = _btb_0_bht_T_8 & _btb_477_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_477_bht_T_20 = _btb_477_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_21 = _btb_477_bht_T_16 ? 2'h0 : _btb_477_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_22 = _btb_477_bht_T_13 ? 2'h0 : _btb_477_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_23 = _btb_477_bht_T_10 ? 2'h0 : _btb_477_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_24 = _btb_477_bht_T_7 ? 2'h3 : _btb_477_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_25 = _btb_477_bht_T_5 ? 2'h3 : _btb_477_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_26 = _btb_477_bht_T_3 ? 2'h3 : _btb_477_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_477_bht_T_27 = _btb_477_bht_T_1 ? 2'h1 : _btb_477_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10614 = btb_477_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7133; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10616 = btb_477_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_477_bht_T_27 : _GEN_8669; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_478_bht_T = btb_478_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_478_bht_T_1 = io_i_branch_resolve_pack_taken & btb_478_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_478_bht_T_2 = btb_478_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_478_bht_T_3 = io_i_branch_resolve_pack_taken & btb_478_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_478_bht_T_4 = btb_478_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_478_bht_T_5 = io_i_branch_resolve_pack_taken & btb_478_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_478_bht_T_6 = btb_478_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_478_bht_T_7 = io_i_branch_resolve_pack_taken & btb_478_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_478_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_478_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_478_bht_T_13 = _btb_0_bht_T_8 & _btb_478_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_478_bht_T_16 = _btb_0_bht_T_8 & _btb_478_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_478_bht_T_19 = _btb_0_bht_T_8 & _btb_478_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_478_bht_T_20 = _btb_478_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_21 = _btb_478_bht_T_16 ? 2'h0 : _btb_478_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_22 = _btb_478_bht_T_13 ? 2'h0 : _btb_478_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_23 = _btb_478_bht_T_10 ? 2'h0 : _btb_478_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_24 = _btb_478_bht_T_7 ? 2'h3 : _btb_478_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_25 = _btb_478_bht_T_5 ? 2'h3 : _btb_478_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_26 = _btb_478_bht_T_3 ? 2'h3 : _btb_478_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_478_bht_T_27 = _btb_478_bht_T_1 ? 2'h1 : _btb_478_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10618 = btb_478_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7134; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10620 = btb_478_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_478_bht_T_27 : _GEN_8670; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_479_bht_T = btb_479_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_479_bht_T_1 = io_i_branch_resolve_pack_taken & btb_479_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_479_bht_T_2 = btb_479_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_479_bht_T_3 = io_i_branch_resolve_pack_taken & btb_479_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_479_bht_T_4 = btb_479_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_479_bht_T_5 = io_i_branch_resolve_pack_taken & btb_479_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_479_bht_T_6 = btb_479_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_479_bht_T_7 = io_i_branch_resolve_pack_taken & btb_479_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_479_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_479_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_479_bht_T_13 = _btb_0_bht_T_8 & _btb_479_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_479_bht_T_16 = _btb_0_bht_T_8 & _btb_479_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_479_bht_T_19 = _btb_0_bht_T_8 & _btb_479_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_479_bht_T_20 = _btb_479_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_21 = _btb_479_bht_T_16 ? 2'h0 : _btb_479_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_22 = _btb_479_bht_T_13 ? 2'h0 : _btb_479_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_23 = _btb_479_bht_T_10 ? 2'h0 : _btb_479_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_24 = _btb_479_bht_T_7 ? 2'h3 : _btb_479_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_25 = _btb_479_bht_T_5 ? 2'h3 : _btb_479_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_26 = _btb_479_bht_T_3 ? 2'h3 : _btb_479_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_479_bht_T_27 = _btb_479_bht_T_1 ? 2'h1 : _btb_479_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10621 = btb_479_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_478_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_477_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_476_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_475_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_474_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_473_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_472_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_471_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_470_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_469_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_468_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_467_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_466_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_465_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10561)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10622 = btb_479_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7135; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10624 = btb_479_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_479_bht_T_27 : _GEN_8671; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_480_bht_T = btb_480_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_480_bht_T_1 = io_i_branch_resolve_pack_taken & btb_480_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_480_bht_T_2 = btb_480_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_480_bht_T_3 = io_i_branch_resolve_pack_taken & btb_480_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_480_bht_T_4 = btb_480_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_480_bht_T_5 = io_i_branch_resolve_pack_taken & btb_480_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_480_bht_T_6 = btb_480_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_480_bht_T_7 = io_i_branch_resolve_pack_taken & btb_480_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_480_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_480_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_480_bht_T_13 = _btb_0_bht_T_8 & _btb_480_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_480_bht_T_16 = _btb_0_bht_T_8 & _btb_480_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_480_bht_T_19 = _btb_0_bht_T_8 & _btb_480_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_480_bht_T_20 = _btb_480_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_21 = _btb_480_bht_T_16 ? 2'h0 : _btb_480_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_22 = _btb_480_bht_T_13 ? 2'h0 : _btb_480_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_23 = _btb_480_bht_T_10 ? 2'h0 : _btb_480_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_24 = _btb_480_bht_T_7 ? 2'h3 : _btb_480_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_25 = _btb_480_bht_T_5 ? 2'h3 : _btb_480_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_26 = _btb_480_bht_T_3 ? 2'h3 : _btb_480_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_480_bht_T_27 = _btb_480_bht_T_1 ? 2'h1 : _btb_480_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10626 = btb_480_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7136; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10628 = btb_480_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_480_bht_T_27 : _GEN_8672; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_481_bht_T = btb_481_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_481_bht_T_1 = io_i_branch_resolve_pack_taken & btb_481_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_481_bht_T_2 = btb_481_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_481_bht_T_3 = io_i_branch_resolve_pack_taken & btb_481_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_481_bht_T_4 = btb_481_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_481_bht_T_5 = io_i_branch_resolve_pack_taken & btb_481_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_481_bht_T_6 = btb_481_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_481_bht_T_7 = io_i_branch_resolve_pack_taken & btb_481_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_481_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_481_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_481_bht_T_13 = _btb_0_bht_T_8 & _btb_481_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_481_bht_T_16 = _btb_0_bht_T_8 & _btb_481_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_481_bht_T_19 = _btb_0_bht_T_8 & _btb_481_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_481_bht_T_20 = _btb_481_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_21 = _btb_481_bht_T_16 ? 2'h0 : _btb_481_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_22 = _btb_481_bht_T_13 ? 2'h0 : _btb_481_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_23 = _btb_481_bht_T_10 ? 2'h0 : _btb_481_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_24 = _btb_481_bht_T_7 ? 2'h3 : _btb_481_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_25 = _btb_481_bht_T_5 ? 2'h3 : _btb_481_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_26 = _btb_481_bht_T_3 ? 2'h3 : _btb_481_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_481_bht_T_27 = _btb_481_bht_T_1 ? 2'h1 : _btb_481_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10630 = btb_481_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7137; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10632 = btb_481_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_481_bht_T_27 : _GEN_8673; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_482_bht_T = btb_482_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_482_bht_T_1 = io_i_branch_resolve_pack_taken & btb_482_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_482_bht_T_2 = btb_482_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_482_bht_T_3 = io_i_branch_resolve_pack_taken & btb_482_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_482_bht_T_4 = btb_482_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_482_bht_T_5 = io_i_branch_resolve_pack_taken & btb_482_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_482_bht_T_6 = btb_482_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_482_bht_T_7 = io_i_branch_resolve_pack_taken & btb_482_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_482_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_482_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_482_bht_T_13 = _btb_0_bht_T_8 & _btb_482_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_482_bht_T_16 = _btb_0_bht_T_8 & _btb_482_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_482_bht_T_19 = _btb_0_bht_T_8 & _btb_482_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_482_bht_T_20 = _btb_482_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_21 = _btb_482_bht_T_16 ? 2'h0 : _btb_482_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_22 = _btb_482_bht_T_13 ? 2'h0 : _btb_482_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_23 = _btb_482_bht_T_10 ? 2'h0 : _btb_482_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_24 = _btb_482_bht_T_7 ? 2'h3 : _btb_482_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_25 = _btb_482_bht_T_5 ? 2'h3 : _btb_482_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_26 = _btb_482_bht_T_3 ? 2'h3 : _btb_482_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_482_bht_T_27 = _btb_482_bht_T_1 ? 2'h1 : _btb_482_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10634 = btb_482_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7138; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10636 = btb_482_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_482_bht_T_27 : _GEN_8674; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_483_bht_T = btb_483_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_483_bht_T_1 = io_i_branch_resolve_pack_taken & btb_483_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_483_bht_T_2 = btb_483_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_483_bht_T_3 = io_i_branch_resolve_pack_taken & btb_483_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_483_bht_T_4 = btb_483_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_483_bht_T_5 = io_i_branch_resolve_pack_taken & btb_483_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_483_bht_T_6 = btb_483_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_483_bht_T_7 = io_i_branch_resolve_pack_taken & btb_483_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_483_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_483_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_483_bht_T_13 = _btb_0_bht_T_8 & _btb_483_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_483_bht_T_16 = _btb_0_bht_T_8 & _btb_483_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_483_bht_T_19 = _btb_0_bht_T_8 & _btb_483_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_483_bht_T_20 = _btb_483_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_21 = _btb_483_bht_T_16 ? 2'h0 : _btb_483_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_22 = _btb_483_bht_T_13 ? 2'h0 : _btb_483_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_23 = _btb_483_bht_T_10 ? 2'h0 : _btb_483_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_24 = _btb_483_bht_T_7 ? 2'h3 : _btb_483_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_25 = _btb_483_bht_T_5 ? 2'h3 : _btb_483_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_26 = _btb_483_bht_T_3 ? 2'h3 : _btb_483_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_483_bht_T_27 = _btb_483_bht_T_1 ? 2'h1 : _btb_483_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10638 = btb_483_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7139; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10640 = btb_483_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_483_bht_T_27 : _GEN_8675; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_484_bht_T = btb_484_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_484_bht_T_1 = io_i_branch_resolve_pack_taken & btb_484_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_484_bht_T_2 = btb_484_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_484_bht_T_3 = io_i_branch_resolve_pack_taken & btb_484_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_484_bht_T_4 = btb_484_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_484_bht_T_5 = io_i_branch_resolve_pack_taken & btb_484_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_484_bht_T_6 = btb_484_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_484_bht_T_7 = io_i_branch_resolve_pack_taken & btb_484_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_484_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_484_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_484_bht_T_13 = _btb_0_bht_T_8 & _btb_484_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_484_bht_T_16 = _btb_0_bht_T_8 & _btb_484_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_484_bht_T_19 = _btb_0_bht_T_8 & _btb_484_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_484_bht_T_20 = _btb_484_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_21 = _btb_484_bht_T_16 ? 2'h0 : _btb_484_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_22 = _btb_484_bht_T_13 ? 2'h0 : _btb_484_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_23 = _btb_484_bht_T_10 ? 2'h0 : _btb_484_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_24 = _btb_484_bht_T_7 ? 2'h3 : _btb_484_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_25 = _btb_484_bht_T_5 ? 2'h3 : _btb_484_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_26 = _btb_484_bht_T_3 ? 2'h3 : _btb_484_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_484_bht_T_27 = _btb_484_bht_T_1 ? 2'h1 : _btb_484_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10642 = btb_484_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7140; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10644 = btb_484_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_484_bht_T_27 : _GEN_8676; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_485_bht_T = btb_485_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_485_bht_T_1 = io_i_branch_resolve_pack_taken & btb_485_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_485_bht_T_2 = btb_485_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_485_bht_T_3 = io_i_branch_resolve_pack_taken & btb_485_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_485_bht_T_4 = btb_485_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_485_bht_T_5 = io_i_branch_resolve_pack_taken & btb_485_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_485_bht_T_6 = btb_485_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_485_bht_T_7 = io_i_branch_resolve_pack_taken & btb_485_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_485_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_485_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_485_bht_T_13 = _btb_0_bht_T_8 & _btb_485_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_485_bht_T_16 = _btb_0_bht_T_8 & _btb_485_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_485_bht_T_19 = _btb_0_bht_T_8 & _btb_485_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_485_bht_T_20 = _btb_485_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_21 = _btb_485_bht_T_16 ? 2'h0 : _btb_485_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_22 = _btb_485_bht_T_13 ? 2'h0 : _btb_485_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_23 = _btb_485_bht_T_10 ? 2'h0 : _btb_485_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_24 = _btb_485_bht_T_7 ? 2'h3 : _btb_485_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_25 = _btb_485_bht_T_5 ? 2'h3 : _btb_485_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_26 = _btb_485_bht_T_3 ? 2'h3 : _btb_485_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_485_bht_T_27 = _btb_485_bht_T_1 ? 2'h1 : _btb_485_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10646 = btb_485_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7141; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10648 = btb_485_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_485_bht_T_27 : _GEN_8677; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_486_bht_T = btb_486_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_486_bht_T_1 = io_i_branch_resolve_pack_taken & btb_486_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_486_bht_T_2 = btb_486_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_486_bht_T_3 = io_i_branch_resolve_pack_taken & btb_486_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_486_bht_T_4 = btb_486_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_486_bht_T_5 = io_i_branch_resolve_pack_taken & btb_486_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_486_bht_T_6 = btb_486_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_486_bht_T_7 = io_i_branch_resolve_pack_taken & btb_486_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_486_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_486_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_486_bht_T_13 = _btb_0_bht_T_8 & _btb_486_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_486_bht_T_16 = _btb_0_bht_T_8 & _btb_486_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_486_bht_T_19 = _btb_0_bht_T_8 & _btb_486_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_486_bht_T_20 = _btb_486_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_21 = _btb_486_bht_T_16 ? 2'h0 : _btb_486_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_22 = _btb_486_bht_T_13 ? 2'h0 : _btb_486_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_23 = _btb_486_bht_T_10 ? 2'h0 : _btb_486_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_24 = _btb_486_bht_T_7 ? 2'h3 : _btb_486_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_25 = _btb_486_bht_T_5 ? 2'h3 : _btb_486_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_26 = _btb_486_bht_T_3 ? 2'h3 : _btb_486_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_486_bht_T_27 = _btb_486_bht_T_1 ? 2'h1 : _btb_486_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10650 = btb_486_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7142; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10652 = btb_486_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_486_bht_T_27 : _GEN_8678; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_487_bht_T = btb_487_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_487_bht_T_1 = io_i_branch_resolve_pack_taken & btb_487_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_487_bht_T_2 = btb_487_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_487_bht_T_3 = io_i_branch_resolve_pack_taken & btb_487_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_487_bht_T_4 = btb_487_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_487_bht_T_5 = io_i_branch_resolve_pack_taken & btb_487_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_487_bht_T_6 = btb_487_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_487_bht_T_7 = io_i_branch_resolve_pack_taken & btb_487_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_487_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_487_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_487_bht_T_13 = _btb_0_bht_T_8 & _btb_487_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_487_bht_T_16 = _btb_0_bht_T_8 & _btb_487_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_487_bht_T_19 = _btb_0_bht_T_8 & _btb_487_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_487_bht_T_20 = _btb_487_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_21 = _btb_487_bht_T_16 ? 2'h0 : _btb_487_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_22 = _btb_487_bht_T_13 ? 2'h0 : _btb_487_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_23 = _btb_487_bht_T_10 ? 2'h0 : _btb_487_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_24 = _btb_487_bht_T_7 ? 2'h3 : _btb_487_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_25 = _btb_487_bht_T_5 ? 2'h3 : _btb_487_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_26 = _btb_487_bht_T_3 ? 2'h3 : _btb_487_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_487_bht_T_27 = _btb_487_bht_T_1 ? 2'h1 : _btb_487_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10654 = btb_487_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7143; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10656 = btb_487_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_487_bht_T_27 : _GEN_8679; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_488_bht_T = btb_488_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_488_bht_T_1 = io_i_branch_resolve_pack_taken & btb_488_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_488_bht_T_2 = btb_488_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_488_bht_T_3 = io_i_branch_resolve_pack_taken & btb_488_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_488_bht_T_4 = btb_488_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_488_bht_T_5 = io_i_branch_resolve_pack_taken & btb_488_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_488_bht_T_6 = btb_488_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_488_bht_T_7 = io_i_branch_resolve_pack_taken & btb_488_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_488_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_488_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_488_bht_T_13 = _btb_0_bht_T_8 & _btb_488_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_488_bht_T_16 = _btb_0_bht_T_8 & _btb_488_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_488_bht_T_19 = _btb_0_bht_T_8 & _btb_488_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_488_bht_T_20 = _btb_488_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_21 = _btb_488_bht_T_16 ? 2'h0 : _btb_488_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_22 = _btb_488_bht_T_13 ? 2'h0 : _btb_488_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_23 = _btb_488_bht_T_10 ? 2'h0 : _btb_488_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_24 = _btb_488_bht_T_7 ? 2'h3 : _btb_488_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_25 = _btb_488_bht_T_5 ? 2'h3 : _btb_488_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_26 = _btb_488_bht_T_3 ? 2'h3 : _btb_488_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_488_bht_T_27 = _btb_488_bht_T_1 ? 2'h1 : _btb_488_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10658 = btb_488_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7144; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10660 = btb_488_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_488_bht_T_27 : _GEN_8680; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_489_bht_T = btb_489_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_489_bht_T_1 = io_i_branch_resolve_pack_taken & btb_489_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_489_bht_T_2 = btb_489_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_489_bht_T_3 = io_i_branch_resolve_pack_taken & btb_489_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_489_bht_T_4 = btb_489_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_489_bht_T_5 = io_i_branch_resolve_pack_taken & btb_489_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_489_bht_T_6 = btb_489_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_489_bht_T_7 = io_i_branch_resolve_pack_taken & btb_489_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_489_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_489_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_489_bht_T_13 = _btb_0_bht_T_8 & _btb_489_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_489_bht_T_16 = _btb_0_bht_T_8 & _btb_489_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_489_bht_T_19 = _btb_0_bht_T_8 & _btb_489_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_489_bht_T_20 = _btb_489_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_21 = _btb_489_bht_T_16 ? 2'h0 : _btb_489_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_22 = _btb_489_bht_T_13 ? 2'h0 : _btb_489_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_23 = _btb_489_bht_T_10 ? 2'h0 : _btb_489_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_24 = _btb_489_bht_T_7 ? 2'h3 : _btb_489_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_25 = _btb_489_bht_T_5 ? 2'h3 : _btb_489_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_26 = _btb_489_bht_T_3 ? 2'h3 : _btb_489_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_489_bht_T_27 = _btb_489_bht_T_1 ? 2'h1 : _btb_489_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10662 = btb_489_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7145; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10664 = btb_489_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_489_bht_T_27 : _GEN_8681; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_490_bht_T = btb_490_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_490_bht_T_1 = io_i_branch_resolve_pack_taken & btb_490_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_490_bht_T_2 = btb_490_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_490_bht_T_3 = io_i_branch_resolve_pack_taken & btb_490_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_490_bht_T_4 = btb_490_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_490_bht_T_5 = io_i_branch_resolve_pack_taken & btb_490_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_490_bht_T_6 = btb_490_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_490_bht_T_7 = io_i_branch_resolve_pack_taken & btb_490_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_490_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_490_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_490_bht_T_13 = _btb_0_bht_T_8 & _btb_490_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_490_bht_T_16 = _btb_0_bht_T_8 & _btb_490_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_490_bht_T_19 = _btb_0_bht_T_8 & _btb_490_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_490_bht_T_20 = _btb_490_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_21 = _btb_490_bht_T_16 ? 2'h0 : _btb_490_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_22 = _btb_490_bht_T_13 ? 2'h0 : _btb_490_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_23 = _btb_490_bht_T_10 ? 2'h0 : _btb_490_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_24 = _btb_490_bht_T_7 ? 2'h3 : _btb_490_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_25 = _btb_490_bht_T_5 ? 2'h3 : _btb_490_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_26 = _btb_490_bht_T_3 ? 2'h3 : _btb_490_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_490_bht_T_27 = _btb_490_bht_T_1 ? 2'h1 : _btb_490_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10666 = btb_490_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7146; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10668 = btb_490_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_490_bht_T_27 : _GEN_8682; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_491_bht_T = btb_491_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_491_bht_T_1 = io_i_branch_resolve_pack_taken & btb_491_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_491_bht_T_2 = btb_491_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_491_bht_T_3 = io_i_branch_resolve_pack_taken & btb_491_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_491_bht_T_4 = btb_491_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_491_bht_T_5 = io_i_branch_resolve_pack_taken & btb_491_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_491_bht_T_6 = btb_491_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_491_bht_T_7 = io_i_branch_resolve_pack_taken & btb_491_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_491_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_491_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_491_bht_T_13 = _btb_0_bht_T_8 & _btb_491_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_491_bht_T_16 = _btb_0_bht_T_8 & _btb_491_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_491_bht_T_19 = _btb_0_bht_T_8 & _btb_491_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_491_bht_T_20 = _btb_491_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_21 = _btb_491_bht_T_16 ? 2'h0 : _btb_491_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_22 = _btb_491_bht_T_13 ? 2'h0 : _btb_491_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_23 = _btb_491_bht_T_10 ? 2'h0 : _btb_491_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_24 = _btb_491_bht_T_7 ? 2'h3 : _btb_491_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_25 = _btb_491_bht_T_5 ? 2'h3 : _btb_491_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_26 = _btb_491_bht_T_3 ? 2'h3 : _btb_491_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_491_bht_T_27 = _btb_491_bht_T_1 ? 2'h1 : _btb_491_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10670 = btb_491_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7147; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10672 = btb_491_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_491_bht_T_27 : _GEN_8683; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_492_bht_T = btb_492_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_492_bht_T_1 = io_i_branch_resolve_pack_taken & btb_492_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_492_bht_T_2 = btb_492_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_492_bht_T_3 = io_i_branch_resolve_pack_taken & btb_492_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_492_bht_T_4 = btb_492_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_492_bht_T_5 = io_i_branch_resolve_pack_taken & btb_492_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_492_bht_T_6 = btb_492_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_492_bht_T_7 = io_i_branch_resolve_pack_taken & btb_492_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_492_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_492_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_492_bht_T_13 = _btb_0_bht_T_8 & _btb_492_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_492_bht_T_16 = _btb_0_bht_T_8 & _btb_492_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_492_bht_T_19 = _btb_0_bht_T_8 & _btb_492_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_492_bht_T_20 = _btb_492_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_21 = _btb_492_bht_T_16 ? 2'h0 : _btb_492_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_22 = _btb_492_bht_T_13 ? 2'h0 : _btb_492_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_23 = _btb_492_bht_T_10 ? 2'h0 : _btb_492_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_24 = _btb_492_bht_T_7 ? 2'h3 : _btb_492_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_25 = _btb_492_bht_T_5 ? 2'h3 : _btb_492_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_26 = _btb_492_bht_T_3 ? 2'h3 : _btb_492_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_492_bht_T_27 = _btb_492_bht_T_1 ? 2'h1 : _btb_492_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10674 = btb_492_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7148; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10676 = btb_492_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_492_bht_T_27 : _GEN_8684; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_493_bht_T = btb_493_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_493_bht_T_1 = io_i_branch_resolve_pack_taken & btb_493_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_493_bht_T_2 = btb_493_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_493_bht_T_3 = io_i_branch_resolve_pack_taken & btb_493_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_493_bht_T_4 = btb_493_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_493_bht_T_5 = io_i_branch_resolve_pack_taken & btb_493_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_493_bht_T_6 = btb_493_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_493_bht_T_7 = io_i_branch_resolve_pack_taken & btb_493_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_493_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_493_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_493_bht_T_13 = _btb_0_bht_T_8 & _btb_493_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_493_bht_T_16 = _btb_0_bht_T_8 & _btb_493_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_493_bht_T_19 = _btb_0_bht_T_8 & _btb_493_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_493_bht_T_20 = _btb_493_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_21 = _btb_493_bht_T_16 ? 2'h0 : _btb_493_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_22 = _btb_493_bht_T_13 ? 2'h0 : _btb_493_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_23 = _btb_493_bht_T_10 ? 2'h0 : _btb_493_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_24 = _btb_493_bht_T_7 ? 2'h3 : _btb_493_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_25 = _btb_493_bht_T_5 ? 2'h3 : _btb_493_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_26 = _btb_493_bht_T_3 ? 2'h3 : _btb_493_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_493_bht_T_27 = _btb_493_bht_T_1 ? 2'h1 : _btb_493_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10678 = btb_493_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7149; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10680 = btb_493_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_493_bht_T_27 : _GEN_8685; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_494_bht_T = btb_494_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_494_bht_T_1 = io_i_branch_resolve_pack_taken & btb_494_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_494_bht_T_2 = btb_494_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_494_bht_T_3 = io_i_branch_resolve_pack_taken & btb_494_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_494_bht_T_4 = btb_494_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_494_bht_T_5 = io_i_branch_resolve_pack_taken & btb_494_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_494_bht_T_6 = btb_494_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_494_bht_T_7 = io_i_branch_resolve_pack_taken & btb_494_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_494_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_494_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_494_bht_T_13 = _btb_0_bht_T_8 & _btb_494_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_494_bht_T_16 = _btb_0_bht_T_8 & _btb_494_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_494_bht_T_19 = _btb_0_bht_T_8 & _btb_494_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_494_bht_T_20 = _btb_494_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_21 = _btb_494_bht_T_16 ? 2'h0 : _btb_494_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_22 = _btb_494_bht_T_13 ? 2'h0 : _btb_494_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_23 = _btb_494_bht_T_10 ? 2'h0 : _btb_494_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_24 = _btb_494_bht_T_7 ? 2'h3 : _btb_494_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_25 = _btb_494_bht_T_5 ? 2'h3 : _btb_494_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_26 = _btb_494_bht_T_3 ? 2'h3 : _btb_494_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_494_bht_T_27 = _btb_494_bht_T_1 ? 2'h1 : _btb_494_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10681 = btb_494_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_493_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_492_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_491_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_490_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_489_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_488_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_487_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_486_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_485_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_484_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_483_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_482_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_481_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_480_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10621)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10682 = btb_494_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7150; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10684 = btb_494_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_494_bht_T_27 : _GEN_8686; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_495_bht_T = btb_495_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_495_bht_T_1 = io_i_branch_resolve_pack_taken & btb_495_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_495_bht_T_2 = btb_495_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_495_bht_T_3 = io_i_branch_resolve_pack_taken & btb_495_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_495_bht_T_4 = btb_495_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_495_bht_T_5 = io_i_branch_resolve_pack_taken & btb_495_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_495_bht_T_6 = btb_495_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_495_bht_T_7 = io_i_branch_resolve_pack_taken & btb_495_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_495_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_495_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_495_bht_T_13 = _btb_0_bht_T_8 & _btb_495_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_495_bht_T_16 = _btb_0_bht_T_8 & _btb_495_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_495_bht_T_19 = _btb_0_bht_T_8 & _btb_495_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_495_bht_T_20 = _btb_495_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_21 = _btb_495_bht_T_16 ? 2'h0 : _btb_495_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_22 = _btb_495_bht_T_13 ? 2'h0 : _btb_495_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_23 = _btb_495_bht_T_10 ? 2'h0 : _btb_495_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_24 = _btb_495_bht_T_7 ? 2'h3 : _btb_495_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_25 = _btb_495_bht_T_5 ? 2'h3 : _btb_495_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_26 = _btb_495_bht_T_3 ? 2'h3 : _btb_495_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_495_bht_T_27 = _btb_495_bht_T_1 ? 2'h1 : _btb_495_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10686 = btb_495_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7151; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10688 = btb_495_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_495_bht_T_27 : _GEN_8687; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_496_bht_T = btb_496_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_496_bht_T_1 = io_i_branch_resolve_pack_taken & btb_496_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_496_bht_T_2 = btb_496_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_496_bht_T_3 = io_i_branch_resolve_pack_taken & btb_496_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_496_bht_T_4 = btb_496_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_496_bht_T_5 = io_i_branch_resolve_pack_taken & btb_496_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_496_bht_T_6 = btb_496_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_496_bht_T_7 = io_i_branch_resolve_pack_taken & btb_496_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_496_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_496_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_496_bht_T_13 = _btb_0_bht_T_8 & _btb_496_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_496_bht_T_16 = _btb_0_bht_T_8 & _btb_496_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_496_bht_T_19 = _btb_0_bht_T_8 & _btb_496_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_496_bht_T_20 = _btb_496_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_21 = _btb_496_bht_T_16 ? 2'h0 : _btb_496_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_22 = _btb_496_bht_T_13 ? 2'h0 : _btb_496_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_23 = _btb_496_bht_T_10 ? 2'h0 : _btb_496_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_24 = _btb_496_bht_T_7 ? 2'h3 : _btb_496_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_25 = _btb_496_bht_T_5 ? 2'h3 : _btb_496_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_26 = _btb_496_bht_T_3 ? 2'h3 : _btb_496_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_496_bht_T_27 = _btb_496_bht_T_1 ? 2'h1 : _btb_496_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10690 = btb_496_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7152; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10692 = btb_496_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_496_bht_T_27 : _GEN_8688; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_497_bht_T = btb_497_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_497_bht_T_1 = io_i_branch_resolve_pack_taken & btb_497_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_497_bht_T_2 = btb_497_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_497_bht_T_3 = io_i_branch_resolve_pack_taken & btb_497_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_497_bht_T_4 = btb_497_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_497_bht_T_5 = io_i_branch_resolve_pack_taken & btb_497_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_497_bht_T_6 = btb_497_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_497_bht_T_7 = io_i_branch_resolve_pack_taken & btb_497_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_497_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_497_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_497_bht_T_13 = _btb_0_bht_T_8 & _btb_497_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_497_bht_T_16 = _btb_0_bht_T_8 & _btb_497_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_497_bht_T_19 = _btb_0_bht_T_8 & _btb_497_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_497_bht_T_20 = _btb_497_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_21 = _btb_497_bht_T_16 ? 2'h0 : _btb_497_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_22 = _btb_497_bht_T_13 ? 2'h0 : _btb_497_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_23 = _btb_497_bht_T_10 ? 2'h0 : _btb_497_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_24 = _btb_497_bht_T_7 ? 2'h3 : _btb_497_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_25 = _btb_497_bht_T_5 ? 2'h3 : _btb_497_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_26 = _btb_497_bht_T_3 ? 2'h3 : _btb_497_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_497_bht_T_27 = _btb_497_bht_T_1 ? 2'h1 : _btb_497_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10694 = btb_497_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7153; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10696 = btb_497_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_497_bht_T_27 : _GEN_8689; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_498_bht_T = btb_498_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_498_bht_T_1 = io_i_branch_resolve_pack_taken & btb_498_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_498_bht_T_2 = btb_498_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_498_bht_T_3 = io_i_branch_resolve_pack_taken & btb_498_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_498_bht_T_4 = btb_498_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_498_bht_T_5 = io_i_branch_resolve_pack_taken & btb_498_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_498_bht_T_6 = btb_498_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_498_bht_T_7 = io_i_branch_resolve_pack_taken & btb_498_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_498_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_498_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_498_bht_T_13 = _btb_0_bht_T_8 & _btb_498_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_498_bht_T_16 = _btb_0_bht_T_8 & _btb_498_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_498_bht_T_19 = _btb_0_bht_T_8 & _btb_498_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_498_bht_T_20 = _btb_498_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_21 = _btb_498_bht_T_16 ? 2'h0 : _btb_498_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_22 = _btb_498_bht_T_13 ? 2'h0 : _btb_498_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_23 = _btb_498_bht_T_10 ? 2'h0 : _btb_498_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_24 = _btb_498_bht_T_7 ? 2'h3 : _btb_498_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_25 = _btb_498_bht_T_5 ? 2'h3 : _btb_498_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_26 = _btb_498_bht_T_3 ? 2'h3 : _btb_498_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_498_bht_T_27 = _btb_498_bht_T_1 ? 2'h1 : _btb_498_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10698 = btb_498_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7154; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10700 = btb_498_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_498_bht_T_27 : _GEN_8690; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_499_bht_T = btb_499_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_499_bht_T_1 = io_i_branch_resolve_pack_taken & btb_499_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_499_bht_T_2 = btb_499_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_499_bht_T_3 = io_i_branch_resolve_pack_taken & btb_499_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_499_bht_T_4 = btb_499_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_499_bht_T_5 = io_i_branch_resolve_pack_taken & btb_499_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_499_bht_T_6 = btb_499_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_499_bht_T_7 = io_i_branch_resolve_pack_taken & btb_499_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_499_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_499_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_499_bht_T_13 = _btb_0_bht_T_8 & _btb_499_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_499_bht_T_16 = _btb_0_bht_T_8 & _btb_499_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_499_bht_T_19 = _btb_0_bht_T_8 & _btb_499_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_499_bht_T_20 = _btb_499_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_21 = _btb_499_bht_T_16 ? 2'h0 : _btb_499_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_22 = _btb_499_bht_T_13 ? 2'h0 : _btb_499_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_23 = _btb_499_bht_T_10 ? 2'h0 : _btb_499_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_24 = _btb_499_bht_T_7 ? 2'h3 : _btb_499_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_25 = _btb_499_bht_T_5 ? 2'h3 : _btb_499_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_26 = _btb_499_bht_T_3 ? 2'h3 : _btb_499_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_499_bht_T_27 = _btb_499_bht_T_1 ? 2'h1 : _btb_499_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10702 = btb_499_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7155; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10704 = btb_499_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_499_bht_T_27 : _GEN_8691; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_500_bht_T = btb_500_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_500_bht_T_1 = io_i_branch_resolve_pack_taken & btb_500_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_500_bht_T_2 = btb_500_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_500_bht_T_3 = io_i_branch_resolve_pack_taken & btb_500_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_500_bht_T_4 = btb_500_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_500_bht_T_5 = io_i_branch_resolve_pack_taken & btb_500_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_500_bht_T_6 = btb_500_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_500_bht_T_7 = io_i_branch_resolve_pack_taken & btb_500_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_500_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_500_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_500_bht_T_13 = _btb_0_bht_T_8 & _btb_500_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_500_bht_T_16 = _btb_0_bht_T_8 & _btb_500_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_500_bht_T_19 = _btb_0_bht_T_8 & _btb_500_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_500_bht_T_20 = _btb_500_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_21 = _btb_500_bht_T_16 ? 2'h0 : _btb_500_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_22 = _btb_500_bht_T_13 ? 2'h0 : _btb_500_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_23 = _btb_500_bht_T_10 ? 2'h0 : _btb_500_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_24 = _btb_500_bht_T_7 ? 2'h3 : _btb_500_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_25 = _btb_500_bht_T_5 ? 2'h3 : _btb_500_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_26 = _btb_500_bht_T_3 ? 2'h3 : _btb_500_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_500_bht_T_27 = _btb_500_bht_T_1 ? 2'h1 : _btb_500_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10706 = btb_500_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7156; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10708 = btb_500_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_500_bht_T_27 : _GEN_8692; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_501_bht_T = btb_501_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_501_bht_T_1 = io_i_branch_resolve_pack_taken & btb_501_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_501_bht_T_2 = btb_501_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_501_bht_T_3 = io_i_branch_resolve_pack_taken & btb_501_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_501_bht_T_4 = btb_501_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_501_bht_T_5 = io_i_branch_resolve_pack_taken & btb_501_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_501_bht_T_6 = btb_501_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_501_bht_T_7 = io_i_branch_resolve_pack_taken & btb_501_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_501_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_501_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_501_bht_T_13 = _btb_0_bht_T_8 & _btb_501_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_501_bht_T_16 = _btb_0_bht_T_8 & _btb_501_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_501_bht_T_19 = _btb_0_bht_T_8 & _btb_501_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_501_bht_T_20 = _btb_501_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_21 = _btb_501_bht_T_16 ? 2'h0 : _btb_501_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_22 = _btb_501_bht_T_13 ? 2'h0 : _btb_501_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_23 = _btb_501_bht_T_10 ? 2'h0 : _btb_501_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_24 = _btb_501_bht_T_7 ? 2'h3 : _btb_501_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_25 = _btb_501_bht_T_5 ? 2'h3 : _btb_501_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_26 = _btb_501_bht_T_3 ? 2'h3 : _btb_501_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_501_bht_T_27 = _btb_501_bht_T_1 ? 2'h1 : _btb_501_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10710 = btb_501_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7157; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10712 = btb_501_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_501_bht_T_27 : _GEN_8693; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_502_bht_T = btb_502_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_502_bht_T_1 = io_i_branch_resolve_pack_taken & btb_502_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_502_bht_T_2 = btb_502_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_502_bht_T_3 = io_i_branch_resolve_pack_taken & btb_502_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_502_bht_T_4 = btb_502_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_502_bht_T_5 = io_i_branch_resolve_pack_taken & btb_502_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_502_bht_T_6 = btb_502_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_502_bht_T_7 = io_i_branch_resolve_pack_taken & btb_502_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_502_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_502_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_502_bht_T_13 = _btb_0_bht_T_8 & _btb_502_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_502_bht_T_16 = _btb_0_bht_T_8 & _btb_502_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_502_bht_T_19 = _btb_0_bht_T_8 & _btb_502_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_502_bht_T_20 = _btb_502_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_21 = _btb_502_bht_T_16 ? 2'h0 : _btb_502_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_22 = _btb_502_bht_T_13 ? 2'h0 : _btb_502_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_23 = _btb_502_bht_T_10 ? 2'h0 : _btb_502_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_24 = _btb_502_bht_T_7 ? 2'h3 : _btb_502_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_25 = _btb_502_bht_T_5 ? 2'h3 : _btb_502_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_26 = _btb_502_bht_T_3 ? 2'h3 : _btb_502_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_502_bht_T_27 = _btb_502_bht_T_1 ? 2'h1 : _btb_502_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10714 = btb_502_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7158; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10716 = btb_502_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_502_bht_T_27 : _GEN_8694; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_503_bht_T = btb_503_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_503_bht_T_1 = io_i_branch_resolve_pack_taken & btb_503_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_503_bht_T_2 = btb_503_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_503_bht_T_3 = io_i_branch_resolve_pack_taken & btb_503_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_503_bht_T_4 = btb_503_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_503_bht_T_5 = io_i_branch_resolve_pack_taken & btb_503_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_503_bht_T_6 = btb_503_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_503_bht_T_7 = io_i_branch_resolve_pack_taken & btb_503_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_503_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_503_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_503_bht_T_13 = _btb_0_bht_T_8 & _btb_503_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_503_bht_T_16 = _btb_0_bht_T_8 & _btb_503_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_503_bht_T_19 = _btb_0_bht_T_8 & _btb_503_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_503_bht_T_20 = _btb_503_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_21 = _btb_503_bht_T_16 ? 2'h0 : _btb_503_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_22 = _btb_503_bht_T_13 ? 2'h0 : _btb_503_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_23 = _btb_503_bht_T_10 ? 2'h0 : _btb_503_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_24 = _btb_503_bht_T_7 ? 2'h3 : _btb_503_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_25 = _btb_503_bht_T_5 ? 2'h3 : _btb_503_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_26 = _btb_503_bht_T_3 ? 2'h3 : _btb_503_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_503_bht_T_27 = _btb_503_bht_T_1 ? 2'h1 : _btb_503_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10718 = btb_503_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7159; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10720 = btb_503_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_503_bht_T_27 : _GEN_8695; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_504_bht_T = btb_504_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_504_bht_T_1 = io_i_branch_resolve_pack_taken & btb_504_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_504_bht_T_2 = btb_504_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_504_bht_T_3 = io_i_branch_resolve_pack_taken & btb_504_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_504_bht_T_4 = btb_504_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_504_bht_T_5 = io_i_branch_resolve_pack_taken & btb_504_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_504_bht_T_6 = btb_504_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_504_bht_T_7 = io_i_branch_resolve_pack_taken & btb_504_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_504_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_504_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_504_bht_T_13 = _btb_0_bht_T_8 & _btb_504_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_504_bht_T_16 = _btb_0_bht_T_8 & _btb_504_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_504_bht_T_19 = _btb_0_bht_T_8 & _btb_504_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_504_bht_T_20 = _btb_504_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_21 = _btb_504_bht_T_16 ? 2'h0 : _btb_504_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_22 = _btb_504_bht_T_13 ? 2'h0 : _btb_504_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_23 = _btb_504_bht_T_10 ? 2'h0 : _btb_504_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_24 = _btb_504_bht_T_7 ? 2'h3 : _btb_504_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_25 = _btb_504_bht_T_5 ? 2'h3 : _btb_504_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_26 = _btb_504_bht_T_3 ? 2'h3 : _btb_504_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_504_bht_T_27 = _btb_504_bht_T_1 ? 2'h1 : _btb_504_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10722 = btb_504_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7160; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10724 = btb_504_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_504_bht_T_27 : _GEN_8696; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_505_bht_T = btb_505_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_505_bht_T_1 = io_i_branch_resolve_pack_taken & btb_505_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_505_bht_T_2 = btb_505_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_505_bht_T_3 = io_i_branch_resolve_pack_taken & btb_505_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_505_bht_T_4 = btb_505_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_505_bht_T_5 = io_i_branch_resolve_pack_taken & btb_505_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_505_bht_T_6 = btb_505_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_505_bht_T_7 = io_i_branch_resolve_pack_taken & btb_505_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_505_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_505_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_505_bht_T_13 = _btb_0_bht_T_8 & _btb_505_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_505_bht_T_16 = _btb_0_bht_T_8 & _btb_505_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_505_bht_T_19 = _btb_0_bht_T_8 & _btb_505_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_505_bht_T_20 = _btb_505_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_21 = _btb_505_bht_T_16 ? 2'h0 : _btb_505_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_22 = _btb_505_bht_T_13 ? 2'h0 : _btb_505_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_23 = _btb_505_bht_T_10 ? 2'h0 : _btb_505_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_24 = _btb_505_bht_T_7 ? 2'h3 : _btb_505_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_25 = _btb_505_bht_T_5 ? 2'h3 : _btb_505_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_26 = _btb_505_bht_T_3 ? 2'h3 : _btb_505_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_505_bht_T_27 = _btb_505_bht_T_1 ? 2'h1 : _btb_505_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10726 = btb_505_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7161; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10728 = btb_505_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_505_bht_T_27 : _GEN_8697; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_506_bht_T = btb_506_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_506_bht_T_1 = io_i_branch_resolve_pack_taken & btb_506_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_506_bht_T_2 = btb_506_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_506_bht_T_3 = io_i_branch_resolve_pack_taken & btb_506_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_506_bht_T_4 = btb_506_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_506_bht_T_5 = io_i_branch_resolve_pack_taken & btb_506_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_506_bht_T_6 = btb_506_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_506_bht_T_7 = io_i_branch_resolve_pack_taken & btb_506_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_506_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_506_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_506_bht_T_13 = _btb_0_bht_T_8 & _btb_506_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_506_bht_T_16 = _btb_0_bht_T_8 & _btb_506_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_506_bht_T_19 = _btb_0_bht_T_8 & _btb_506_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_506_bht_T_20 = _btb_506_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_21 = _btb_506_bht_T_16 ? 2'h0 : _btb_506_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_22 = _btb_506_bht_T_13 ? 2'h0 : _btb_506_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_23 = _btb_506_bht_T_10 ? 2'h0 : _btb_506_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_24 = _btb_506_bht_T_7 ? 2'h3 : _btb_506_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_25 = _btb_506_bht_T_5 ? 2'h3 : _btb_506_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_26 = _btb_506_bht_T_3 ? 2'h3 : _btb_506_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_506_bht_T_27 = _btb_506_bht_T_1 ? 2'h1 : _btb_506_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10730 = btb_506_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7162; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10732 = btb_506_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_506_bht_T_27 : _GEN_8698; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_507_bht_T = btb_507_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_507_bht_T_1 = io_i_branch_resolve_pack_taken & btb_507_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_507_bht_T_2 = btb_507_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_507_bht_T_3 = io_i_branch_resolve_pack_taken & btb_507_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_507_bht_T_4 = btb_507_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_507_bht_T_5 = io_i_branch_resolve_pack_taken & btb_507_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_507_bht_T_6 = btb_507_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_507_bht_T_7 = io_i_branch_resolve_pack_taken & btb_507_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_507_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_507_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_507_bht_T_13 = _btb_0_bht_T_8 & _btb_507_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_507_bht_T_16 = _btb_0_bht_T_8 & _btb_507_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_507_bht_T_19 = _btb_0_bht_T_8 & _btb_507_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_507_bht_T_20 = _btb_507_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_21 = _btb_507_bht_T_16 ? 2'h0 : _btb_507_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_22 = _btb_507_bht_T_13 ? 2'h0 : _btb_507_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_23 = _btb_507_bht_T_10 ? 2'h0 : _btb_507_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_24 = _btb_507_bht_T_7 ? 2'h3 : _btb_507_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_25 = _btb_507_bht_T_5 ? 2'h3 : _btb_507_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_26 = _btb_507_bht_T_3 ? 2'h3 : _btb_507_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_507_bht_T_27 = _btb_507_bht_T_1 ? 2'h1 : _btb_507_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10734 = btb_507_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7163; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10736 = btb_507_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_507_bht_T_27 : _GEN_8699; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_508_bht_T = btb_508_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_508_bht_T_1 = io_i_branch_resolve_pack_taken & btb_508_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_508_bht_T_2 = btb_508_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_508_bht_T_3 = io_i_branch_resolve_pack_taken & btb_508_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_508_bht_T_4 = btb_508_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_508_bht_T_5 = io_i_branch_resolve_pack_taken & btb_508_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_508_bht_T_6 = btb_508_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_508_bht_T_7 = io_i_branch_resolve_pack_taken & btb_508_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_508_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_508_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_508_bht_T_13 = _btb_0_bht_T_8 & _btb_508_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_508_bht_T_16 = _btb_0_bht_T_8 & _btb_508_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_508_bht_T_19 = _btb_0_bht_T_8 & _btb_508_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_508_bht_T_20 = _btb_508_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_21 = _btb_508_bht_T_16 ? 2'h0 : _btb_508_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_22 = _btb_508_bht_T_13 ? 2'h0 : _btb_508_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_23 = _btb_508_bht_T_10 ? 2'h0 : _btb_508_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_24 = _btb_508_bht_T_7 ? 2'h3 : _btb_508_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_25 = _btb_508_bht_T_5 ? 2'h3 : _btb_508_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_26 = _btb_508_bht_T_3 ? 2'h3 : _btb_508_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_508_bht_T_27 = _btb_508_bht_T_1 ? 2'h1 : _btb_508_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10738 = btb_508_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7164; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10740 = btb_508_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_508_bht_T_27 : _GEN_8700; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_509_bht_T = btb_509_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_509_bht_T_1 = io_i_branch_resolve_pack_taken & btb_509_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_509_bht_T_2 = btb_509_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_509_bht_T_3 = io_i_branch_resolve_pack_taken & btb_509_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_509_bht_T_4 = btb_509_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_509_bht_T_5 = io_i_branch_resolve_pack_taken & btb_509_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_509_bht_T_6 = btb_509_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_509_bht_T_7 = io_i_branch_resolve_pack_taken & btb_509_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_509_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_509_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_509_bht_T_13 = _btb_0_bht_T_8 & _btb_509_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_509_bht_T_16 = _btb_0_bht_T_8 & _btb_509_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_509_bht_T_19 = _btb_0_bht_T_8 & _btb_509_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_509_bht_T_20 = _btb_509_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_21 = _btb_509_bht_T_16 ? 2'h0 : _btb_509_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_22 = _btb_509_bht_T_13 ? 2'h0 : _btb_509_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_23 = _btb_509_bht_T_10 ? 2'h0 : _btb_509_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_24 = _btb_509_bht_T_7 ? 2'h3 : _btb_509_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_25 = _btb_509_bht_T_5 ? 2'h3 : _btb_509_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_26 = _btb_509_bht_T_3 ? 2'h3 : _btb_509_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_509_bht_T_27 = _btb_509_bht_T_1 ? 2'h1 : _btb_509_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10741 = btb_509_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_508_tag == io_i_branch_resolve_pack_pc[12:3
    ] | (btb_507_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_506_tag == io_i_branch_resolve_pack_pc[12:3] | (
    btb_505_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_504_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_503_tag
     == io_i_branch_resolve_pack_pc[12:3] | (btb_502_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_501_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_500_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_499_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_498_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_497_tag ==
    io_i_branch_resolve_pack_pc[12:3] | (btb_496_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_495_tag ==
    io_i_branch_resolve_pack_pc[12:3] | _GEN_10681)))))))))))))); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10742 = btb_509_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7165; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10744 = btb_509_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_509_bht_T_27 : _GEN_8701; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_510_bht_T = btb_510_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_510_bht_T_1 = io_i_branch_resolve_pack_taken & btb_510_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_510_bht_T_2 = btb_510_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_510_bht_T_3 = io_i_branch_resolve_pack_taken & btb_510_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_510_bht_T_4 = btb_510_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_510_bht_T_5 = io_i_branch_resolve_pack_taken & btb_510_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_510_bht_T_6 = btb_510_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_510_bht_T_7 = io_i_branch_resolve_pack_taken & btb_510_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_510_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_510_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_510_bht_T_13 = _btb_0_bht_T_8 & _btb_510_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_510_bht_T_16 = _btb_0_bht_T_8 & _btb_510_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_510_bht_T_19 = _btb_0_bht_T_8 & _btb_510_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_510_bht_T_20 = _btb_510_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_21 = _btb_510_bht_T_16 ? 2'h0 : _btb_510_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_22 = _btb_510_bht_T_13 ? 2'h0 : _btb_510_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_23 = _btb_510_bht_T_10 ? 2'h0 : _btb_510_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_24 = _btb_510_bht_T_7 ? 2'h3 : _btb_510_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_25 = _btb_510_bht_T_5 ? 2'h3 : _btb_510_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_26 = _btb_510_bht_T_3 ? 2'h3 : _btb_510_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_510_bht_T_27 = _btb_510_bht_T_1 ? 2'h1 : _btb_510_bht_T_26; // @[Mux.scala 101:16]
  wire [63:0] _GEN_10746 = btb_510_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7166; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10748 = btb_510_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_510_bht_T_27 : _GEN_8702; // @[branch_predictor.scala 79:71 83:32]
  wire  _btb_511_bht_T = btb_511_bht == 2'h0; // @[branch_predictor.scala 84:67]
  wire  _btb_511_bht_T_1 = io_i_branch_resolve_pack_taken & btb_511_bht == 2'h0; // @[branch_predictor.scala 84:53]
  wire  _btb_511_bht_T_2 = btb_511_bht == 2'h1; // @[branch_predictor.scala 85:67]
  wire  _btb_511_bht_T_3 = io_i_branch_resolve_pack_taken & btb_511_bht == 2'h1; // @[branch_predictor.scala 85:53]
  wire  _btb_511_bht_T_4 = btb_511_bht == 2'h2; // @[branch_predictor.scala 86:67]
  wire  _btb_511_bht_T_5 = io_i_branch_resolve_pack_taken & btb_511_bht == 2'h2; // @[branch_predictor.scala 86:53]
  wire  _btb_511_bht_T_6 = btb_511_bht == 2'h3; // @[branch_predictor.scala 87:67]
  wire  _btb_511_bht_T_7 = io_i_branch_resolve_pack_taken & btb_511_bht == 2'h3; // @[branch_predictor.scala 87:53]
  wire  _btb_511_bht_T_10 = ~io_i_branch_resolve_pack_taken & _btb_511_bht_T; // @[branch_predictor.scala 89:54]
  wire  _btb_511_bht_T_13 = _btb_0_bht_T_8 & _btb_511_bht_T_2; // @[branch_predictor.scala 90:54]
  wire  _btb_511_bht_T_16 = _btb_0_bht_T_8 & _btb_511_bht_T_4; // @[branch_predictor.scala 91:54]
  wire  _btb_511_bht_T_19 = _btb_0_bht_T_8 & _btb_511_bht_T_6; // @[branch_predictor.scala 92:54]
  wire [1:0] _btb_511_bht_T_20 = _btb_511_bht_T_19 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_21 = _btb_511_bht_T_16 ? 2'h0 : _btb_511_bht_T_20; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_22 = _btb_511_bht_T_13 ? 2'h0 : _btb_511_bht_T_21; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_23 = _btb_511_bht_T_10 ? 2'h0 : _btb_511_bht_T_22; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_24 = _btb_511_bht_T_7 ? 2'h3 : _btb_511_bht_T_23; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_25 = _btb_511_bht_T_5 ? 2'h3 : _btb_511_bht_T_24; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_26 = _btb_511_bht_T_3 ? 2'h3 : _btb_511_bht_T_25; // @[Mux.scala 101:16]
  wire [1:0] _btb_511_bht_T_27 = _btb_511_bht_T_1 ? 2'h1 : _btb_511_bht_T_26; // @[Mux.scala 101:16]
  wire  _GEN_10749 = btb_511_tag == io_i_branch_resolve_pack_pc[12:3] | (btb_510_tag == io_i_branch_resolve_pack_pc[12:3
    ] | _GEN_10741); // @[branch_predictor.scala 79:71 80:33]
  wire [63:0] _GEN_10750 = btb_511_tag == io_i_branch_resolve_pack_pc[12:3] ? io_i_branch_resolve_pack_target :
    _GEN_7167; // @[branch_predictor.scala 79:71 81:43]
  wire [1:0] _GEN_10752 = btb_511_tag == io_i_branch_resolve_pack_pc[12:3] ? _btb_511_bht_T_27 : _GEN_8703; // @[branch_predictor.scala 79:71 83:32]
  wire  entry_found = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid & _GEN_10749; // @[branch_predictor.scala 76:17 77:87]
  wire [63:0] _GEN_10754 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8706 :
    _GEN_6656; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10756 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8708 :
    _GEN_8192; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10757 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8710 :
    _GEN_6657; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10759 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8712 :
    _GEN_8193; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10760 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8714 :
    _GEN_6658; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10762 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8716 :
    _GEN_8194; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10763 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8718 :
    _GEN_6659; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10765 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8720 :
    _GEN_8195; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10766 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8722 :
    _GEN_6660; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10768 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8724 :
    _GEN_8196; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10769 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8726 :
    _GEN_6661; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10771 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8728 :
    _GEN_8197; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10772 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8730 :
    _GEN_6662; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10774 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8732 :
    _GEN_8198; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10775 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8734 :
    _GEN_6663; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10777 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8736 :
    _GEN_8199; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10778 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8738 :
    _GEN_6664; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10780 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8740 :
    _GEN_8200; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10781 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8742 :
    _GEN_6665; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10783 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8744 :
    _GEN_8201; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10784 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8746 :
    _GEN_6666; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10786 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8748 :
    _GEN_8202; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10787 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8750 :
    _GEN_6667; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10789 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8752 :
    _GEN_8203; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10790 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8754 :
    _GEN_6668; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10792 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8756 :
    _GEN_8204; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10793 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8758 :
    _GEN_6669; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10795 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8760 :
    _GEN_8205; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10796 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8762 :
    _GEN_6670; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10798 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8764 :
    _GEN_8206; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10799 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8766 :
    _GEN_6671; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10801 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8768 :
    _GEN_8207; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10802 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8770 :
    _GEN_6672; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10804 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8772 :
    _GEN_8208; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10805 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8774 :
    _GEN_6673; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10807 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8776 :
    _GEN_8209; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10808 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8778 :
    _GEN_6674; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10810 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8780 :
    _GEN_8210; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10811 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8782 :
    _GEN_6675; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10813 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8784 :
    _GEN_8211; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10814 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8786 :
    _GEN_6676; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10816 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8788 :
    _GEN_8212; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10817 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8790 :
    _GEN_6677; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10819 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8792 :
    _GEN_8213; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10820 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8794 :
    _GEN_6678; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10822 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8796 :
    _GEN_8214; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10823 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8798 :
    _GEN_6679; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10825 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8800 :
    _GEN_8215; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10826 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8802 :
    _GEN_6680; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10828 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8804 :
    _GEN_8216; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10829 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8806 :
    _GEN_6681; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10831 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8808 :
    _GEN_8217; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10832 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8810 :
    _GEN_6682; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10834 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8812 :
    _GEN_8218; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10835 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8814 :
    _GEN_6683; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10837 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8816 :
    _GEN_8219; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10838 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8818 :
    _GEN_6684; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10840 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8820 :
    _GEN_8220; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10841 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8822 :
    _GEN_6685; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10843 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8824 :
    _GEN_8221; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10844 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8826 :
    _GEN_6686; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10846 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8828 :
    _GEN_8222; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10847 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8830 :
    _GEN_6687; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10849 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8832 :
    _GEN_8223; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10850 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8834 :
    _GEN_6688; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10852 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8836 :
    _GEN_8224; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10853 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8838 :
    _GEN_6689; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10855 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8840 :
    _GEN_8225; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10856 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8842 :
    _GEN_6690; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10858 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8844 :
    _GEN_8226; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10859 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8846 :
    _GEN_6691; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10861 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8848 :
    _GEN_8227; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10862 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8850 :
    _GEN_6692; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10864 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8852 :
    _GEN_8228; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10865 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8854 :
    _GEN_6693; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10867 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8856 :
    _GEN_8229; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10868 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8858 :
    _GEN_6694; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10870 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8860 :
    _GEN_8230; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10871 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8862 :
    _GEN_6695; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10873 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8864 :
    _GEN_8231; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10874 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8866 :
    _GEN_6696; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10876 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8868 :
    _GEN_8232; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10877 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8870 :
    _GEN_6697; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10879 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8872 :
    _GEN_8233; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10880 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8874 :
    _GEN_6698; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10882 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8876 :
    _GEN_8234; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10883 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8878 :
    _GEN_6699; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10885 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8880 :
    _GEN_8235; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10886 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8882 :
    _GEN_6700; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10888 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8884 :
    _GEN_8236; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10889 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8886 :
    _GEN_6701; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10891 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8888 :
    _GEN_8237; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10892 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8890 :
    _GEN_6702; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10894 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8892 :
    _GEN_8238; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10895 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8894 :
    _GEN_6703; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10897 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8896 :
    _GEN_8239; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10898 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8898 :
    _GEN_6704; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10900 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8900 :
    _GEN_8240; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10901 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8902 :
    _GEN_6705; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10903 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8904 :
    _GEN_8241; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10904 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8906 :
    _GEN_6706; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10906 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8908 :
    _GEN_8242; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10907 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8910 :
    _GEN_6707; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10909 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8912 :
    _GEN_8243; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10910 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8914 :
    _GEN_6708; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10912 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8916 :
    _GEN_8244; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10913 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8918 :
    _GEN_6709; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10915 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8920 :
    _GEN_8245; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10916 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8922 :
    _GEN_6710; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10918 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8924 :
    _GEN_8246; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10919 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8926 :
    _GEN_6711; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10921 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8928 :
    _GEN_8247; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10922 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8930 :
    _GEN_6712; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10924 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8932 :
    _GEN_8248; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10925 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8934 :
    _GEN_6713; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10927 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8936 :
    _GEN_8249; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10928 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8938 :
    _GEN_6714; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10930 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8940 :
    _GEN_8250; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10931 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8942 :
    _GEN_6715; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10933 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8944 :
    _GEN_8251; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10934 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8946 :
    _GEN_6716; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10936 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8948 :
    _GEN_8252; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10937 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8950 :
    _GEN_6717; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10939 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8952 :
    _GEN_8253; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10940 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8954 :
    _GEN_6718; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10942 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8956 :
    _GEN_8254; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10943 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8958 :
    _GEN_6719; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10945 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8960 :
    _GEN_8255; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10946 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8962 :
    _GEN_6720; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10948 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8964 :
    _GEN_8256; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10949 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8966 :
    _GEN_6721; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10951 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8968 :
    _GEN_8257; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10952 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8970 :
    _GEN_6722; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10954 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8972 :
    _GEN_8258; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10955 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8974 :
    _GEN_6723; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10957 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8976 :
    _GEN_8259; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10958 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8978 :
    _GEN_6724; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10960 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8980 :
    _GEN_8260; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10961 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8982 :
    _GEN_6725; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10963 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8984 :
    _GEN_8261; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10964 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8986 :
    _GEN_6726; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10966 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8988 :
    _GEN_8262; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10967 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8990 :
    _GEN_6727; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10969 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8992 :
    _GEN_8263; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10970 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8994 :
    _GEN_6728; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10972 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8996 :
    _GEN_8264; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10973 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_8998 :
    _GEN_6729; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10975 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9000 :
    _GEN_8265; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10976 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9002 :
    _GEN_6730; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10978 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9004 :
    _GEN_8266; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10979 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9006 :
    _GEN_6731; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10981 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9008 :
    _GEN_8267; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10982 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9010 :
    _GEN_6732; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10984 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9012 :
    _GEN_8268; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10985 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9014 :
    _GEN_6733; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10987 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9016 :
    _GEN_8269; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10988 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9018 :
    _GEN_6734; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10990 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9020 :
    _GEN_8270; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10991 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9022 :
    _GEN_6735; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10993 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9024 :
    _GEN_8271; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10994 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9026 :
    _GEN_6736; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10996 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9028 :
    _GEN_8272; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_10997 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9030 :
    _GEN_6737; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_10999 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9032 :
    _GEN_8273; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11000 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9034 :
    _GEN_6738; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11002 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9036 :
    _GEN_8274; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11003 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9038 :
    _GEN_6739; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11005 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9040 :
    _GEN_8275; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11006 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9042 :
    _GEN_6740; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11008 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9044 :
    _GEN_8276; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11009 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9046 :
    _GEN_6741; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11011 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9048 :
    _GEN_8277; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11012 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9050 :
    _GEN_6742; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11014 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9052 :
    _GEN_8278; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11015 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9054 :
    _GEN_6743; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11017 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9056 :
    _GEN_8279; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11018 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9058 :
    _GEN_6744; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11020 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9060 :
    _GEN_8280; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11021 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9062 :
    _GEN_6745; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11023 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9064 :
    _GEN_8281; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11024 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9066 :
    _GEN_6746; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11026 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9068 :
    _GEN_8282; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11027 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9070 :
    _GEN_6747; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11029 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9072 :
    _GEN_8283; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11030 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9074 :
    _GEN_6748; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11032 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9076 :
    _GEN_8284; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11033 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9078 :
    _GEN_6749; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11035 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9080 :
    _GEN_8285; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11036 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9082 :
    _GEN_6750; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11038 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9084 :
    _GEN_8286; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11039 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9086 :
    _GEN_6751; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11041 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9088 :
    _GEN_8287; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11042 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9090 :
    _GEN_6752; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11044 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9092 :
    _GEN_8288; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11045 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9094 :
    _GEN_6753; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11047 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9096 :
    _GEN_8289; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11048 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9098 :
    _GEN_6754; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11050 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9100 :
    _GEN_8290; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11051 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9102 :
    _GEN_6755; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11053 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9104 :
    _GEN_8291; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11054 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9106 :
    _GEN_6756; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11056 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9108 :
    _GEN_8292; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11057 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9110 :
    _GEN_6757; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11059 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9112 :
    _GEN_8293; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11060 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9114 :
    _GEN_6758; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11062 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9116 :
    _GEN_8294; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11063 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9118 :
    _GEN_6759; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11065 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9120 :
    _GEN_8295; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11066 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9122 :
    _GEN_6760; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11068 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9124 :
    _GEN_8296; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11069 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9126 :
    _GEN_6761; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11071 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9128 :
    _GEN_8297; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11072 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9130 :
    _GEN_6762; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11074 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9132 :
    _GEN_8298; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11075 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9134 :
    _GEN_6763; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11077 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9136 :
    _GEN_8299; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11078 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9138 :
    _GEN_6764; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11080 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9140 :
    _GEN_8300; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11081 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9142 :
    _GEN_6765; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11083 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9144 :
    _GEN_8301; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11084 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9146 :
    _GEN_6766; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11086 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9148 :
    _GEN_8302; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11087 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9150 :
    _GEN_6767; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11089 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9152 :
    _GEN_8303; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11090 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9154 :
    _GEN_6768; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11092 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9156 :
    _GEN_8304; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11093 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9158 :
    _GEN_6769; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11095 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9160 :
    _GEN_8305; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11096 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9162 :
    _GEN_6770; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11098 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9164 :
    _GEN_8306; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11099 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9166 :
    _GEN_6771; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11101 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9168 :
    _GEN_8307; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11102 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9170 :
    _GEN_6772; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11104 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9172 :
    _GEN_8308; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11105 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9174 :
    _GEN_6773; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11107 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9176 :
    _GEN_8309; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11108 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9178 :
    _GEN_6774; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11110 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9180 :
    _GEN_8310; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11111 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9182 :
    _GEN_6775; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11113 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9184 :
    _GEN_8311; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11114 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9186 :
    _GEN_6776; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11116 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9188 :
    _GEN_8312; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11117 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9190 :
    _GEN_6777; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11119 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9192 :
    _GEN_8313; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11120 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9194 :
    _GEN_6778; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11122 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9196 :
    _GEN_8314; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11123 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9198 :
    _GEN_6779; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11125 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9200 :
    _GEN_8315; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11126 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9202 :
    _GEN_6780; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11128 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9204 :
    _GEN_8316; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11129 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9206 :
    _GEN_6781; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11131 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9208 :
    _GEN_8317; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11132 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9210 :
    _GEN_6782; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11134 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9212 :
    _GEN_8318; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11135 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9214 :
    _GEN_6783; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11137 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9216 :
    _GEN_8319; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11138 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9218 :
    _GEN_6784; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11140 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9220 :
    _GEN_8320; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11141 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9222 :
    _GEN_6785; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11143 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9224 :
    _GEN_8321; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11144 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9226 :
    _GEN_6786; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11146 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9228 :
    _GEN_8322; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11147 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9230 :
    _GEN_6787; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11149 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9232 :
    _GEN_8323; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11150 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9234 :
    _GEN_6788; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11152 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9236 :
    _GEN_8324; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11153 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9238 :
    _GEN_6789; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11155 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9240 :
    _GEN_8325; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11156 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9242 :
    _GEN_6790; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11158 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9244 :
    _GEN_8326; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11159 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9246 :
    _GEN_6791; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11161 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9248 :
    _GEN_8327; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11162 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9250 :
    _GEN_6792; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11164 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9252 :
    _GEN_8328; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11165 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9254 :
    _GEN_6793; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11167 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9256 :
    _GEN_8329; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11168 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9258 :
    _GEN_6794; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11170 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9260 :
    _GEN_8330; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11171 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9262 :
    _GEN_6795; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11173 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9264 :
    _GEN_8331; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11174 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9266 :
    _GEN_6796; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11176 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9268 :
    _GEN_8332; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11177 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9270 :
    _GEN_6797; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11179 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9272 :
    _GEN_8333; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11180 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9274 :
    _GEN_6798; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11182 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9276 :
    _GEN_8334; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11183 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9278 :
    _GEN_6799; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11185 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9280 :
    _GEN_8335; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11186 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9282 :
    _GEN_6800; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11188 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9284 :
    _GEN_8336; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11189 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9286 :
    _GEN_6801; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11191 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9288 :
    _GEN_8337; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11192 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9290 :
    _GEN_6802; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11194 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9292 :
    _GEN_8338; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11195 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9294 :
    _GEN_6803; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11197 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9296 :
    _GEN_8339; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11198 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9298 :
    _GEN_6804; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11200 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9300 :
    _GEN_8340; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11201 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9302 :
    _GEN_6805; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11203 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9304 :
    _GEN_8341; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11204 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9306 :
    _GEN_6806; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11206 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9308 :
    _GEN_8342; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11207 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9310 :
    _GEN_6807; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11209 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9312 :
    _GEN_8343; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11210 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9314 :
    _GEN_6808; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11212 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9316 :
    _GEN_8344; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11213 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9318 :
    _GEN_6809; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11215 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9320 :
    _GEN_8345; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11216 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9322 :
    _GEN_6810; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11218 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9324 :
    _GEN_8346; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11219 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9326 :
    _GEN_6811; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11221 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9328 :
    _GEN_8347; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11222 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9330 :
    _GEN_6812; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11224 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9332 :
    _GEN_8348; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11225 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9334 :
    _GEN_6813; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11227 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9336 :
    _GEN_8349; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11228 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9338 :
    _GEN_6814; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11230 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9340 :
    _GEN_8350; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11231 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9342 :
    _GEN_6815; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11233 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9344 :
    _GEN_8351; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11234 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9346 :
    _GEN_6816; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11236 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9348 :
    _GEN_8352; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11237 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9350 :
    _GEN_6817; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11239 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9352 :
    _GEN_8353; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11240 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9354 :
    _GEN_6818; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11242 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9356 :
    _GEN_8354; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11243 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9358 :
    _GEN_6819; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11245 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9360 :
    _GEN_8355; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11246 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9362 :
    _GEN_6820; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11248 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9364 :
    _GEN_8356; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11249 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9366 :
    _GEN_6821; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11251 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9368 :
    _GEN_8357; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11252 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9370 :
    _GEN_6822; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11254 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9372 :
    _GEN_8358; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11255 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9374 :
    _GEN_6823; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11257 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9376 :
    _GEN_8359; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11258 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9378 :
    _GEN_6824; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11260 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9380 :
    _GEN_8360; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11261 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9382 :
    _GEN_6825; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11263 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9384 :
    _GEN_8361; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11264 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9386 :
    _GEN_6826; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11266 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9388 :
    _GEN_8362; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11267 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9390 :
    _GEN_6827; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11269 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9392 :
    _GEN_8363; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11270 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9394 :
    _GEN_6828; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11272 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9396 :
    _GEN_8364; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11273 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9398 :
    _GEN_6829; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11275 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9400 :
    _GEN_8365; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11276 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9402 :
    _GEN_6830; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11278 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9404 :
    _GEN_8366; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11279 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9406 :
    _GEN_6831; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11281 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9408 :
    _GEN_8367; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11282 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9410 :
    _GEN_6832; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11284 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9412 :
    _GEN_8368; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11285 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9414 :
    _GEN_6833; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11287 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9416 :
    _GEN_8369; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11288 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9418 :
    _GEN_6834; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11290 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9420 :
    _GEN_8370; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11291 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9422 :
    _GEN_6835; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11293 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9424 :
    _GEN_8371; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11294 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9426 :
    _GEN_6836; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11296 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9428 :
    _GEN_8372; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11297 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9430 :
    _GEN_6837; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11299 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9432 :
    _GEN_8373; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11300 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9434 :
    _GEN_6838; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11302 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9436 :
    _GEN_8374; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11303 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9438 :
    _GEN_6839; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11305 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9440 :
    _GEN_8375; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11306 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9442 :
    _GEN_6840; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11308 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9444 :
    _GEN_8376; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11309 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9446 :
    _GEN_6841; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11311 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9448 :
    _GEN_8377; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11312 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9450 :
    _GEN_6842; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11314 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9452 :
    _GEN_8378; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11315 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9454 :
    _GEN_6843; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11317 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9456 :
    _GEN_8379; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11318 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9458 :
    _GEN_6844; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11320 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9460 :
    _GEN_8380; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11321 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9462 :
    _GEN_6845; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11323 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9464 :
    _GEN_8381; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11324 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9466 :
    _GEN_6846; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11326 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9468 :
    _GEN_8382; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11327 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9470 :
    _GEN_6847; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11329 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9472 :
    _GEN_8383; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11330 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9474 :
    _GEN_6848; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11332 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9476 :
    _GEN_8384; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11333 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9478 :
    _GEN_6849; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11335 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9480 :
    _GEN_8385; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11336 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9482 :
    _GEN_6850; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11338 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9484 :
    _GEN_8386; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11339 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9486 :
    _GEN_6851; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11341 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9488 :
    _GEN_8387; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11342 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9490 :
    _GEN_6852; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11344 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9492 :
    _GEN_8388; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11345 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9494 :
    _GEN_6853; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11347 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9496 :
    _GEN_8389; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11348 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9498 :
    _GEN_6854; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11350 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9500 :
    _GEN_8390; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11351 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9502 :
    _GEN_6855; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11353 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9504 :
    _GEN_8391; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11354 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9506 :
    _GEN_6856; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11356 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9508 :
    _GEN_8392; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11357 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9510 :
    _GEN_6857; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11359 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9512 :
    _GEN_8393; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11360 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9514 :
    _GEN_6858; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11362 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9516 :
    _GEN_8394; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11363 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9518 :
    _GEN_6859; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11365 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9520 :
    _GEN_8395; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11366 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9522 :
    _GEN_6860; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11368 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9524 :
    _GEN_8396; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11369 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9526 :
    _GEN_6861; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11371 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9528 :
    _GEN_8397; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11372 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9530 :
    _GEN_6862; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11374 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9532 :
    _GEN_8398; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11375 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9534 :
    _GEN_6863; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11377 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9536 :
    _GEN_8399; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11378 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9538 :
    _GEN_6864; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11380 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9540 :
    _GEN_8400; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11381 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9542 :
    _GEN_6865; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11383 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9544 :
    _GEN_8401; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11384 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9546 :
    _GEN_6866; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11386 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9548 :
    _GEN_8402; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11387 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9550 :
    _GEN_6867; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11389 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9552 :
    _GEN_8403; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11390 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9554 :
    _GEN_6868; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11392 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9556 :
    _GEN_8404; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11393 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9558 :
    _GEN_6869; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11395 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9560 :
    _GEN_8405; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11396 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9562 :
    _GEN_6870; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11398 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9564 :
    _GEN_8406; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11399 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9566 :
    _GEN_6871; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11401 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9568 :
    _GEN_8407; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11402 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9570 :
    _GEN_6872; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11404 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9572 :
    _GEN_8408; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11405 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9574 :
    _GEN_6873; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11407 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9576 :
    _GEN_8409; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11408 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9578 :
    _GEN_6874; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11410 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9580 :
    _GEN_8410; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11411 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9582 :
    _GEN_6875; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11413 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9584 :
    _GEN_8411; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11414 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9586 :
    _GEN_6876; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11416 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9588 :
    _GEN_8412; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11417 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9590 :
    _GEN_6877; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11419 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9592 :
    _GEN_8413; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11420 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9594 :
    _GEN_6878; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11422 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9596 :
    _GEN_8414; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11423 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9598 :
    _GEN_6879; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11425 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9600 :
    _GEN_8415; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11426 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9602 :
    _GEN_6880; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11428 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9604 :
    _GEN_8416; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11429 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9606 :
    _GEN_6881; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11431 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9608 :
    _GEN_8417; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11432 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9610 :
    _GEN_6882; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11434 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9612 :
    _GEN_8418; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11435 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9614 :
    _GEN_6883; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11437 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9616 :
    _GEN_8419; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11438 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9618 :
    _GEN_6884; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11440 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9620 :
    _GEN_8420; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11441 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9622 :
    _GEN_6885; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11443 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9624 :
    _GEN_8421; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11444 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9626 :
    _GEN_6886; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11446 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9628 :
    _GEN_8422; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11447 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9630 :
    _GEN_6887; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11449 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9632 :
    _GEN_8423; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11450 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9634 :
    _GEN_6888; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11452 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9636 :
    _GEN_8424; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11453 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9638 :
    _GEN_6889; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11455 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9640 :
    _GEN_8425; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11456 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9642 :
    _GEN_6890; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11458 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9644 :
    _GEN_8426; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11459 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9646 :
    _GEN_6891; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11461 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9648 :
    _GEN_8427; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11462 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9650 :
    _GEN_6892; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11464 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9652 :
    _GEN_8428; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11465 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9654 :
    _GEN_6893; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11467 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9656 :
    _GEN_8429; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11468 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9658 :
    _GEN_6894; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11470 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9660 :
    _GEN_8430; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11471 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9662 :
    _GEN_6895; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11473 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9664 :
    _GEN_8431; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11474 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9666 :
    _GEN_6896; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11476 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9668 :
    _GEN_8432; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11477 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9670 :
    _GEN_6897; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11479 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9672 :
    _GEN_8433; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11480 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9674 :
    _GEN_6898; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11482 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9676 :
    _GEN_8434; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11483 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9678 :
    _GEN_6899; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11485 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9680 :
    _GEN_8435; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11486 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9682 :
    _GEN_6900; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11488 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9684 :
    _GEN_8436; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11489 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9686 :
    _GEN_6901; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11491 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9688 :
    _GEN_8437; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11492 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9690 :
    _GEN_6902; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11494 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9692 :
    _GEN_8438; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11495 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9694 :
    _GEN_6903; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11497 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9696 :
    _GEN_8439; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11498 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9698 :
    _GEN_6904; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11500 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9700 :
    _GEN_8440; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11501 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9702 :
    _GEN_6905; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11503 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9704 :
    _GEN_8441; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11504 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9706 :
    _GEN_6906; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11506 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9708 :
    _GEN_8442; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11507 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9710 :
    _GEN_6907; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11509 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9712 :
    _GEN_8443; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11510 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9714 :
    _GEN_6908; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11512 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9716 :
    _GEN_8444; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11513 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9718 :
    _GEN_6909; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11515 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9720 :
    _GEN_8445; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11516 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9722 :
    _GEN_6910; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11518 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9724 :
    _GEN_8446; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11519 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9726 :
    _GEN_6911; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11521 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9728 :
    _GEN_8447; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11522 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9730 :
    _GEN_6912; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11524 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9732 :
    _GEN_8448; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11525 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9734 :
    _GEN_6913; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11527 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9736 :
    _GEN_8449; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11528 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9738 :
    _GEN_6914; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11530 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9740 :
    _GEN_8450; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11531 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9742 :
    _GEN_6915; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11533 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9744 :
    _GEN_8451; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11534 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9746 :
    _GEN_6916; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11536 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9748 :
    _GEN_8452; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11537 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9750 :
    _GEN_6917; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11539 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9752 :
    _GEN_8453; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11540 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9754 :
    _GEN_6918; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11542 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9756 :
    _GEN_8454; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11543 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9758 :
    _GEN_6919; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11545 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9760 :
    _GEN_8455; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11546 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9762 :
    _GEN_6920; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11548 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9764 :
    _GEN_8456; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11549 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9766 :
    _GEN_6921; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11551 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9768 :
    _GEN_8457; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11552 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9770 :
    _GEN_6922; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11554 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9772 :
    _GEN_8458; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11555 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9774 :
    _GEN_6923; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11557 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9776 :
    _GEN_8459; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11558 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9778 :
    _GEN_6924; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11560 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9780 :
    _GEN_8460; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11561 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9782 :
    _GEN_6925; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11563 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9784 :
    _GEN_8461; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11564 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9786 :
    _GEN_6926; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11566 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9788 :
    _GEN_8462; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11567 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9790 :
    _GEN_6927; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11569 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9792 :
    _GEN_8463; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11570 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9794 :
    _GEN_6928; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11572 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9796 :
    _GEN_8464; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11573 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9798 :
    _GEN_6929; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11575 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9800 :
    _GEN_8465; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11576 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9802 :
    _GEN_6930; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11578 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9804 :
    _GEN_8466; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11579 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9806 :
    _GEN_6931; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11581 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9808 :
    _GEN_8467; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11582 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9810 :
    _GEN_6932; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11584 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9812 :
    _GEN_8468; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11585 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9814 :
    _GEN_6933; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11587 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9816 :
    _GEN_8469; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11588 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9818 :
    _GEN_6934; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11590 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9820 :
    _GEN_8470; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11591 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9822 :
    _GEN_6935; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11593 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9824 :
    _GEN_8471; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11594 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9826 :
    _GEN_6936; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11596 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9828 :
    _GEN_8472; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11597 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9830 :
    _GEN_6937; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11599 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9832 :
    _GEN_8473; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11600 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9834 :
    _GEN_6938; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11602 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9836 :
    _GEN_8474; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11603 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9838 :
    _GEN_6939; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11605 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9840 :
    _GEN_8475; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11606 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9842 :
    _GEN_6940; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11608 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9844 :
    _GEN_8476; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11609 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9846 :
    _GEN_6941; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11611 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9848 :
    _GEN_8477; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11612 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9850 :
    _GEN_6942; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11614 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9852 :
    _GEN_8478; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11615 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9854 :
    _GEN_6943; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11617 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9856 :
    _GEN_8479; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11618 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9858 :
    _GEN_6944; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11620 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9860 :
    _GEN_8480; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11621 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9862 :
    _GEN_6945; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11623 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9864 :
    _GEN_8481; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11624 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9866 :
    _GEN_6946; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11626 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9868 :
    _GEN_8482; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11627 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9870 :
    _GEN_6947; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11629 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9872 :
    _GEN_8483; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11630 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9874 :
    _GEN_6948; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11632 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9876 :
    _GEN_8484; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11633 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9878 :
    _GEN_6949; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11635 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9880 :
    _GEN_8485; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11636 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9882 :
    _GEN_6950; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11638 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9884 :
    _GEN_8486; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11639 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9886 :
    _GEN_6951; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11641 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9888 :
    _GEN_8487; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11642 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9890 :
    _GEN_6952; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11644 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9892 :
    _GEN_8488; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11645 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9894 :
    _GEN_6953; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11647 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9896 :
    _GEN_8489; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11648 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9898 :
    _GEN_6954; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11650 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9900 :
    _GEN_8490; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11651 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9902 :
    _GEN_6955; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11653 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9904 :
    _GEN_8491; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11654 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9906 :
    _GEN_6956; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11656 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9908 :
    _GEN_8492; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11657 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9910 :
    _GEN_6957; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11659 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9912 :
    _GEN_8493; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11660 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9914 :
    _GEN_6958; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11662 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9916 :
    _GEN_8494; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11663 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9918 :
    _GEN_6959; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11665 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9920 :
    _GEN_8495; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11666 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9922 :
    _GEN_6960; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11668 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9924 :
    _GEN_8496; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11669 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9926 :
    _GEN_6961; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11671 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9928 :
    _GEN_8497; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11672 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9930 :
    _GEN_6962; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11674 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9932 :
    _GEN_8498; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11675 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9934 :
    _GEN_6963; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11677 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9936 :
    _GEN_8499; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11678 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9938 :
    _GEN_6964; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11680 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9940 :
    _GEN_8500; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11681 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9942 :
    _GEN_6965; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11683 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9944 :
    _GEN_8501; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11684 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9946 :
    _GEN_6966; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11686 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9948 :
    _GEN_8502; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11687 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9950 :
    _GEN_6967; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11689 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9952 :
    _GEN_8503; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11690 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9954 :
    _GEN_6968; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11692 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9956 :
    _GEN_8504; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11693 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9958 :
    _GEN_6969; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11695 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9960 :
    _GEN_8505; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11696 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9962 :
    _GEN_6970; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11698 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9964 :
    _GEN_8506; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11699 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9966 :
    _GEN_6971; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11701 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9968 :
    _GEN_8507; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11702 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9970 :
    _GEN_6972; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11704 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9972 :
    _GEN_8508; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11705 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9974 :
    _GEN_6973; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11707 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9976 :
    _GEN_8509; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11708 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9978 :
    _GEN_6974; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11710 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9980 :
    _GEN_8510; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11711 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9982 :
    _GEN_6975; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11713 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9984 :
    _GEN_8511; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11714 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9986 :
    _GEN_6976; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11716 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9988 :
    _GEN_8512; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11717 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9990 :
    _GEN_6977; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11719 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9992 :
    _GEN_8513; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11720 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9994 :
    _GEN_6978; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11722 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9996 :
    _GEN_8514; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11723 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_9998 :
    _GEN_6979; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11725 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10000 :
    _GEN_8515; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11726 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10002 :
    _GEN_6980; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11728 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10004 :
    _GEN_8516; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11729 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10006 :
    _GEN_6981; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11731 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10008 :
    _GEN_8517; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11732 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10010 :
    _GEN_6982; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11734 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10012 :
    _GEN_8518; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11735 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10014 :
    _GEN_6983; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11737 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10016 :
    _GEN_8519; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11738 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10018 :
    _GEN_6984; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11740 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10020 :
    _GEN_8520; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11741 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10022 :
    _GEN_6985; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11743 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10024 :
    _GEN_8521; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11744 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10026 :
    _GEN_6986; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11746 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10028 :
    _GEN_8522; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11747 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10030 :
    _GEN_6987; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11749 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10032 :
    _GEN_8523; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11750 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10034 :
    _GEN_6988; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11752 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10036 :
    _GEN_8524; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11753 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10038 :
    _GEN_6989; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11755 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10040 :
    _GEN_8525; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11756 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10042 :
    _GEN_6990; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11758 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10044 :
    _GEN_8526; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11759 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10046 :
    _GEN_6991; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11761 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10048 :
    _GEN_8527; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11762 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10050 :
    _GEN_6992; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11764 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10052 :
    _GEN_8528; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11765 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10054 :
    _GEN_6993; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11767 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10056 :
    _GEN_8529; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11768 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10058 :
    _GEN_6994; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11770 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10060 :
    _GEN_8530; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11771 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10062 :
    _GEN_6995; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11773 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10064 :
    _GEN_8531; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11774 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10066 :
    _GEN_6996; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11776 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10068 :
    _GEN_8532; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11777 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10070 :
    _GEN_6997; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11779 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10072 :
    _GEN_8533; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11780 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10074 :
    _GEN_6998; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11782 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10076 :
    _GEN_8534; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11783 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10078 :
    _GEN_6999; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11785 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10080 :
    _GEN_8535; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11786 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10082 :
    _GEN_7000; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11788 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10084 :
    _GEN_8536; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11789 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10086 :
    _GEN_7001; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11791 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10088 :
    _GEN_8537; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11792 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10090 :
    _GEN_7002; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11794 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10092 :
    _GEN_8538; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11795 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10094 :
    _GEN_7003; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11797 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10096 :
    _GEN_8539; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11798 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10098 :
    _GEN_7004; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11800 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10100 :
    _GEN_8540; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11801 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10102 :
    _GEN_7005; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11803 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10104 :
    _GEN_8541; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11804 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10106 :
    _GEN_7006; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11806 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10108 :
    _GEN_8542; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11807 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10110 :
    _GEN_7007; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11809 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10112 :
    _GEN_8543; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11810 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10114 :
    _GEN_7008; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11812 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10116 :
    _GEN_8544; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11813 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10118 :
    _GEN_7009; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11815 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10120 :
    _GEN_8545; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11816 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10122 :
    _GEN_7010; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11818 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10124 :
    _GEN_8546; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11819 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10126 :
    _GEN_7011; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11821 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10128 :
    _GEN_8547; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11822 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10130 :
    _GEN_7012; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11824 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10132 :
    _GEN_8548; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11825 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10134 :
    _GEN_7013; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11827 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10136 :
    _GEN_8549; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11828 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10138 :
    _GEN_7014; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11830 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10140 :
    _GEN_8550; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11831 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10142 :
    _GEN_7015; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11833 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10144 :
    _GEN_8551; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11834 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10146 :
    _GEN_7016; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11836 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10148 :
    _GEN_8552; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11837 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10150 :
    _GEN_7017; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11839 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10152 :
    _GEN_8553; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11840 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10154 :
    _GEN_7018; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11842 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10156 :
    _GEN_8554; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11843 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10158 :
    _GEN_7019; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11845 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10160 :
    _GEN_8555; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11846 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10162 :
    _GEN_7020; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11848 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10164 :
    _GEN_8556; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11849 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10166 :
    _GEN_7021; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11851 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10168 :
    _GEN_8557; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11852 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10170 :
    _GEN_7022; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11854 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10172 :
    _GEN_8558; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11855 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10174 :
    _GEN_7023; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11857 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10176 :
    _GEN_8559; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11858 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10178 :
    _GEN_7024; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11860 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10180 :
    _GEN_8560; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11861 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10182 :
    _GEN_7025; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11863 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10184 :
    _GEN_8561; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11864 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10186 :
    _GEN_7026; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11866 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10188 :
    _GEN_8562; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11867 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10190 :
    _GEN_7027; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11869 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10192 :
    _GEN_8563; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11870 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10194 :
    _GEN_7028; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11872 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10196 :
    _GEN_8564; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11873 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10198 :
    _GEN_7029; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11875 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10200 :
    _GEN_8565; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11876 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10202 :
    _GEN_7030; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11878 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10204 :
    _GEN_8566; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11879 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10206 :
    _GEN_7031; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11881 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10208 :
    _GEN_8567; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11882 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10210 :
    _GEN_7032; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11884 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10212 :
    _GEN_8568; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11885 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10214 :
    _GEN_7033; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11887 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10216 :
    _GEN_8569; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11888 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10218 :
    _GEN_7034; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11890 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10220 :
    _GEN_8570; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11891 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10222 :
    _GEN_7035; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11893 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10224 :
    _GEN_8571; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11894 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10226 :
    _GEN_7036; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11896 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10228 :
    _GEN_8572; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11897 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10230 :
    _GEN_7037; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11899 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10232 :
    _GEN_8573; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11900 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10234 :
    _GEN_7038; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11902 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10236 :
    _GEN_8574; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11903 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10238 :
    _GEN_7039; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11905 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10240 :
    _GEN_8575; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11906 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10242 :
    _GEN_7040; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11908 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10244 :
    _GEN_8576; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11909 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10246 :
    _GEN_7041; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11911 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10248 :
    _GEN_8577; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11912 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10250 :
    _GEN_7042; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11914 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10252 :
    _GEN_8578; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11915 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10254 :
    _GEN_7043; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11917 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10256 :
    _GEN_8579; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11918 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10258 :
    _GEN_7044; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11920 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10260 :
    _GEN_8580; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11921 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10262 :
    _GEN_7045; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11923 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10264 :
    _GEN_8581; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11924 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10266 :
    _GEN_7046; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11926 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10268 :
    _GEN_8582; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11927 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10270 :
    _GEN_7047; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11929 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10272 :
    _GEN_8583; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11930 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10274 :
    _GEN_7048; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11932 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10276 :
    _GEN_8584; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11933 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10278 :
    _GEN_7049; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11935 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10280 :
    _GEN_8585; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11936 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10282 :
    _GEN_7050; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11938 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10284 :
    _GEN_8586; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11939 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10286 :
    _GEN_7051; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11941 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10288 :
    _GEN_8587; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11942 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10290 :
    _GEN_7052; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11944 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10292 :
    _GEN_8588; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11945 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10294 :
    _GEN_7053; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11947 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10296 :
    _GEN_8589; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11948 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10298 :
    _GEN_7054; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11950 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10300 :
    _GEN_8590; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11951 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10302 :
    _GEN_7055; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11953 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10304 :
    _GEN_8591; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11954 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10306 :
    _GEN_7056; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11956 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10308 :
    _GEN_8592; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11957 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10310 :
    _GEN_7057; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11959 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10312 :
    _GEN_8593; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11960 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10314 :
    _GEN_7058; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11962 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10316 :
    _GEN_8594; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11963 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10318 :
    _GEN_7059; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11965 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10320 :
    _GEN_8595; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11966 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10322 :
    _GEN_7060; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11968 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10324 :
    _GEN_8596; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11969 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10326 :
    _GEN_7061; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11971 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10328 :
    _GEN_8597; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11972 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10330 :
    _GEN_7062; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11974 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10332 :
    _GEN_8598; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11975 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10334 :
    _GEN_7063; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11977 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10336 :
    _GEN_8599; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11978 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10338 :
    _GEN_7064; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11980 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10340 :
    _GEN_8600; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11981 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10342 :
    _GEN_7065; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11983 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10344 :
    _GEN_8601; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11984 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10346 :
    _GEN_7066; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11986 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10348 :
    _GEN_8602; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11987 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10350 :
    _GEN_7067; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11989 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10352 :
    _GEN_8603; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11990 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10354 :
    _GEN_7068; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11992 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10356 :
    _GEN_8604; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11993 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10358 :
    _GEN_7069; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11995 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10360 :
    _GEN_8605; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11996 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10362 :
    _GEN_7070; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_11998 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10364 :
    _GEN_8606; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_11999 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10366 :
    _GEN_7071; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12001 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10368 :
    _GEN_8607; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12002 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10370 :
    _GEN_7072; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12004 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10372 :
    _GEN_8608; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12005 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10374 :
    _GEN_7073; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12007 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10376 :
    _GEN_8609; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12008 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10378 :
    _GEN_7074; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12010 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10380 :
    _GEN_8610; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12011 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10382 :
    _GEN_7075; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12013 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10384 :
    _GEN_8611; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12014 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10386 :
    _GEN_7076; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12016 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10388 :
    _GEN_8612; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12017 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10390 :
    _GEN_7077; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12019 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10392 :
    _GEN_8613; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12020 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10394 :
    _GEN_7078; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12022 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10396 :
    _GEN_8614; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12023 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10398 :
    _GEN_7079; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12025 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10400 :
    _GEN_8615; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12026 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10402 :
    _GEN_7080; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12028 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10404 :
    _GEN_8616; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12029 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10406 :
    _GEN_7081; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12031 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10408 :
    _GEN_8617; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12032 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10410 :
    _GEN_7082; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12034 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10412 :
    _GEN_8618; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12035 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10414 :
    _GEN_7083; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12037 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10416 :
    _GEN_8619; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12038 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10418 :
    _GEN_7084; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12040 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10420 :
    _GEN_8620; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12041 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10422 :
    _GEN_7085; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12043 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10424 :
    _GEN_8621; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12044 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10426 :
    _GEN_7086; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12046 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10428 :
    _GEN_8622; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12047 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10430 :
    _GEN_7087; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12049 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10432 :
    _GEN_8623; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12050 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10434 :
    _GEN_7088; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12052 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10436 :
    _GEN_8624; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12053 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10438 :
    _GEN_7089; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12055 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10440 :
    _GEN_8625; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12056 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10442 :
    _GEN_7090; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12058 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10444 :
    _GEN_8626; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12059 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10446 :
    _GEN_7091; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12061 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10448 :
    _GEN_8627; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12062 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10450 :
    _GEN_7092; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12064 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10452 :
    _GEN_8628; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12065 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10454 :
    _GEN_7093; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12067 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10456 :
    _GEN_8629; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12068 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10458 :
    _GEN_7094; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12070 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10460 :
    _GEN_8630; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12071 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10462 :
    _GEN_7095; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12073 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10464 :
    _GEN_8631; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12074 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10466 :
    _GEN_7096; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12076 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10468 :
    _GEN_8632; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12077 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10470 :
    _GEN_7097; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12079 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10472 :
    _GEN_8633; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12080 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10474 :
    _GEN_7098; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12082 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10476 :
    _GEN_8634; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12083 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10478 :
    _GEN_7099; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12085 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10480 :
    _GEN_8635; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12086 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10482 :
    _GEN_7100; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12088 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10484 :
    _GEN_8636; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12089 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10486 :
    _GEN_7101; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12091 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10488 :
    _GEN_8637; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12092 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10490 :
    _GEN_7102; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12094 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10492 :
    _GEN_8638; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12095 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10494 :
    _GEN_7103; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12097 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10496 :
    _GEN_8639; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12098 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10498 :
    _GEN_7104; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12100 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10500 :
    _GEN_8640; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12101 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10502 :
    _GEN_7105; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12103 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10504 :
    _GEN_8641; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12104 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10506 :
    _GEN_7106; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12106 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10508 :
    _GEN_8642; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12107 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10510 :
    _GEN_7107; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12109 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10512 :
    _GEN_8643; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12110 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10514 :
    _GEN_7108; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12112 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10516 :
    _GEN_8644; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12113 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10518 :
    _GEN_7109; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12115 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10520 :
    _GEN_8645; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12116 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10522 :
    _GEN_7110; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12118 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10524 :
    _GEN_8646; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12119 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10526 :
    _GEN_7111; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12121 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10528 :
    _GEN_8647; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12122 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10530 :
    _GEN_7112; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12124 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10532 :
    _GEN_8648; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12125 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10534 :
    _GEN_7113; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12127 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10536 :
    _GEN_8649; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12128 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10538 :
    _GEN_7114; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12130 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10540 :
    _GEN_8650; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12131 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10542 :
    _GEN_7115; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12133 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10544 :
    _GEN_8651; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12134 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10546 :
    _GEN_7116; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12136 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10548 :
    _GEN_8652; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12137 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10550 :
    _GEN_7117; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12139 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10552 :
    _GEN_8653; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12140 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10554 :
    _GEN_7118; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12142 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10556 :
    _GEN_8654; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12143 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10558 :
    _GEN_7119; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12145 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10560 :
    _GEN_8655; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12146 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10562 :
    _GEN_7120; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12148 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10564 :
    _GEN_8656; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12149 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10566 :
    _GEN_7121; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12151 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10568 :
    _GEN_8657; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12152 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10570 :
    _GEN_7122; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12154 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10572 :
    _GEN_8658; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12155 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10574 :
    _GEN_7123; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12157 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10576 :
    _GEN_8659; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12158 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10578 :
    _GEN_7124; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12160 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10580 :
    _GEN_8660; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12161 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10582 :
    _GEN_7125; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12163 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10584 :
    _GEN_8661; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12164 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10586 :
    _GEN_7126; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12166 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10588 :
    _GEN_8662; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12167 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10590 :
    _GEN_7127; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12169 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10592 :
    _GEN_8663; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12170 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10594 :
    _GEN_7128; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12172 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10596 :
    _GEN_8664; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12173 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10598 :
    _GEN_7129; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12175 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10600 :
    _GEN_8665; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12176 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10602 :
    _GEN_7130; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12178 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10604 :
    _GEN_8666; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12179 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10606 :
    _GEN_7131; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12181 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10608 :
    _GEN_8667; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12182 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10610 :
    _GEN_7132; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12184 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10612 :
    _GEN_8668; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12185 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10614 :
    _GEN_7133; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12187 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10616 :
    _GEN_8669; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12188 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10618 :
    _GEN_7134; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12190 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10620 :
    _GEN_8670; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12191 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10622 :
    _GEN_7135; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12193 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10624 :
    _GEN_8671; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12194 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10626 :
    _GEN_7136; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12196 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10628 :
    _GEN_8672; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12197 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10630 :
    _GEN_7137; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12199 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10632 :
    _GEN_8673; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12200 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10634 :
    _GEN_7138; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12202 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10636 :
    _GEN_8674; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12203 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10638 :
    _GEN_7139; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12205 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10640 :
    _GEN_8675; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12206 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10642 :
    _GEN_7140; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12208 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10644 :
    _GEN_8676; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12209 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10646 :
    _GEN_7141; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12211 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10648 :
    _GEN_8677; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12212 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10650 :
    _GEN_7142; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12214 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10652 :
    _GEN_8678; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12215 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10654 :
    _GEN_7143; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12217 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10656 :
    _GEN_8679; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12218 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10658 :
    _GEN_7144; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12220 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10660 :
    _GEN_8680; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12221 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10662 :
    _GEN_7145; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12223 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10664 :
    _GEN_8681; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12224 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10666 :
    _GEN_7146; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12226 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10668 :
    _GEN_8682; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12227 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10670 :
    _GEN_7147; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12229 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10672 :
    _GEN_8683; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12230 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10674 :
    _GEN_7148; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12232 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10676 :
    _GEN_8684; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12233 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10678 :
    _GEN_7149; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12235 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10680 :
    _GEN_8685; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12236 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10682 :
    _GEN_7150; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12238 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10684 :
    _GEN_8686; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12239 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10686 :
    _GEN_7151; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12241 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10688 :
    _GEN_8687; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12242 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10690 :
    _GEN_7152; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12244 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10692 :
    _GEN_8688; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12245 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10694 :
    _GEN_7153; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12247 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10696 :
    _GEN_8689; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12248 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10698 :
    _GEN_7154; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12250 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10700 :
    _GEN_8690; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12251 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10702 :
    _GEN_7155; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12253 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10704 :
    _GEN_8691; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12254 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10706 :
    _GEN_7156; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12256 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10708 :
    _GEN_8692; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12257 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10710 :
    _GEN_7157; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12259 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10712 :
    _GEN_8693; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12260 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10714 :
    _GEN_7158; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12262 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10716 :
    _GEN_8694; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12263 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10718 :
    _GEN_7159; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12265 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10720 :
    _GEN_8695; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12266 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10722 :
    _GEN_7160; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12268 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10724 :
    _GEN_8696; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12269 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10726 :
    _GEN_7161; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12271 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10728 :
    _GEN_8697; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12272 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10730 :
    _GEN_7162; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12274 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10732 :
    _GEN_8698; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12275 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10734 :
    _GEN_7163; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12277 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10736 :
    _GEN_8699; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12278 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10738 :
    _GEN_7164; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12280 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10740 :
    _GEN_8700; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12281 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10742 :
    _GEN_7165; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12283 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10744 :
    _GEN_8701; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12284 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10746 :
    _GEN_7166; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12286 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10748 :
    _GEN_8702; // @[branch_predictor.scala 77:87]
  wire [63:0] _GEN_12287 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10750 :
    _GEN_7167; // @[branch_predictor.scala 77:87]
  wire [1:0] _GEN_12289 = io_i_branch_resolve_pack_valid & io_i_branch_resolve_pack_prediction_valid ? _GEN_10752 :
    _GEN_8703; // @[branch_predictor.scala 77:87]
  wire  _GEN_12290 = _GEN_19459 | _GEN_5632; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12291 = _GEN_19460 | _GEN_5633; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12292 = _GEN_19461 | _GEN_5634; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12293 = _GEN_19462 | _GEN_5635; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12294 = _GEN_19463 | _GEN_5636; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12295 = _GEN_19464 | _GEN_5637; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12296 = _GEN_19465 | _GEN_5638; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12297 = _GEN_19466 | _GEN_5639; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12298 = _GEN_19467 | _GEN_5640; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12299 = _GEN_19468 | _GEN_5641; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12300 = _GEN_19469 | _GEN_5642; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12301 = _GEN_19470 | _GEN_5643; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12302 = _GEN_19471 | _GEN_5644; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12303 = _GEN_19472 | _GEN_5645; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12304 = _GEN_19473 | _GEN_5646; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12305 = _GEN_19474 | _GEN_5647; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12306 = _GEN_19475 | _GEN_5648; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12307 = _GEN_19476 | _GEN_5649; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12308 = _GEN_19477 | _GEN_5650; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12309 = _GEN_19478 | _GEN_5651; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12310 = _GEN_19479 | _GEN_5652; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12311 = _GEN_19480 | _GEN_5653; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12312 = _GEN_19481 | _GEN_5654; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12313 = _GEN_19482 | _GEN_5655; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12314 = _GEN_19483 | _GEN_5656; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12315 = _GEN_19484 | _GEN_5657; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12316 = _GEN_19485 | _GEN_5658; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12317 = _GEN_19486 | _GEN_5659; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12318 = _GEN_19487 | _GEN_5660; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12319 = _GEN_19488 | _GEN_5661; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12320 = _GEN_19489 | _GEN_5662; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12321 = _GEN_19490 | _GEN_5663; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12322 = _GEN_19491 | _GEN_5664; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12323 = _GEN_19492 | _GEN_5665; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12324 = _GEN_19493 | _GEN_5666; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12325 = _GEN_19494 | _GEN_5667; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12326 = _GEN_19495 | _GEN_5668; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12327 = _GEN_19496 | _GEN_5669; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12328 = _GEN_19497 | _GEN_5670; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12329 = _GEN_19498 | _GEN_5671; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12330 = _GEN_19499 | _GEN_5672; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12331 = _GEN_19500 | _GEN_5673; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12332 = _GEN_19501 | _GEN_5674; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12333 = _GEN_19502 | _GEN_5675; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12334 = _GEN_19503 | _GEN_5676; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12335 = _GEN_19504 | _GEN_5677; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12336 = _GEN_19505 | _GEN_5678; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12337 = _GEN_19506 | _GEN_5679; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12338 = _GEN_19507 | _GEN_5680; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12339 = _GEN_19508 | _GEN_5681; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12340 = _GEN_19509 | _GEN_5682; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12341 = _GEN_19510 | _GEN_5683; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12342 = _GEN_19511 | _GEN_5684; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12343 = _GEN_19512 | _GEN_5685; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12344 = _GEN_19513 | _GEN_5686; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12345 = _GEN_19514 | _GEN_5687; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12346 = _GEN_19515 | _GEN_5688; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12347 = _GEN_19516 | _GEN_5689; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12348 = _GEN_19517 | _GEN_5690; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12349 = _GEN_19518 | _GEN_5691; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12350 = _GEN_19519 | _GEN_5692; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12351 = _GEN_19520 | _GEN_5693; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12352 = _GEN_19521 | _GEN_5694; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12353 = _GEN_19522 | _GEN_5695; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12354 = _GEN_19523 | _GEN_5696; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12355 = _GEN_19524 | _GEN_5697; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12356 = _GEN_19525 | _GEN_5698; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12357 = _GEN_19526 | _GEN_5699; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12358 = _GEN_19527 | _GEN_5700; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12359 = _GEN_19528 | _GEN_5701; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12360 = _GEN_19529 | _GEN_5702; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12361 = _GEN_19530 | _GEN_5703; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12362 = _GEN_19531 | _GEN_5704; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12363 = _GEN_19532 | _GEN_5705; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12364 = _GEN_19533 | _GEN_5706; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12365 = _GEN_19534 | _GEN_5707; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12366 = _GEN_19535 | _GEN_5708; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12367 = _GEN_19536 | _GEN_5709; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12368 = _GEN_19537 | _GEN_5710; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12369 = _GEN_19538 | _GEN_5711; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12370 = _GEN_19539 | _GEN_5712; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12371 = _GEN_19540 | _GEN_5713; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12372 = _GEN_19541 | _GEN_5714; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12373 = _GEN_19542 | _GEN_5715; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12374 = _GEN_19543 | _GEN_5716; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12375 = _GEN_19544 | _GEN_5717; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12376 = _GEN_19545 | _GEN_5718; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12377 = _GEN_19546 | _GEN_5719; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12378 = _GEN_19547 | _GEN_5720; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12379 = _GEN_19548 | _GEN_5721; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12380 = _GEN_19549 | _GEN_5722; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12381 = _GEN_19550 | _GEN_5723; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12382 = _GEN_19551 | _GEN_5724; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12383 = _GEN_19552 | _GEN_5725; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12384 = _GEN_19553 | _GEN_5726; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12385 = _GEN_19554 | _GEN_5727; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12386 = _GEN_19555 | _GEN_5728; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12387 = _GEN_19556 | _GEN_5729; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12388 = _GEN_19557 | _GEN_5730; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12389 = _GEN_19558 | _GEN_5731; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12390 = _GEN_19559 | _GEN_5732; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12391 = _GEN_19560 | _GEN_5733; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12392 = _GEN_19561 | _GEN_5734; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12393 = _GEN_19562 | _GEN_5735; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12394 = _GEN_19563 | _GEN_5736; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12395 = _GEN_19564 | _GEN_5737; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12396 = _GEN_19565 | _GEN_5738; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12397 = _GEN_19566 | _GEN_5739; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12398 = _GEN_19567 | _GEN_5740; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12399 = _GEN_19568 | _GEN_5741; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12400 = _GEN_19569 | _GEN_5742; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12401 = _GEN_19570 | _GEN_5743; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12402 = _GEN_19571 | _GEN_5744; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12403 = _GEN_19572 | _GEN_5745; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12404 = _GEN_19573 | _GEN_5746; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12405 = _GEN_19574 | _GEN_5747; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12406 = _GEN_19575 | _GEN_5748; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12407 = _GEN_19576 | _GEN_5749; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12408 = _GEN_19577 | _GEN_5750; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12409 = _GEN_19578 | _GEN_5751; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12410 = _GEN_19579 | _GEN_5752; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12411 = _GEN_19580 | _GEN_5753; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12412 = _GEN_19581 | _GEN_5754; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12413 = _GEN_19582 | _GEN_5755; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12414 = _GEN_19583 | _GEN_5756; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12415 = _GEN_19584 | _GEN_5757; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12416 = _GEN_19585 | _GEN_5758; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12417 = _GEN_19586 | _GEN_5759; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12418 = _GEN_19587 | _GEN_5760; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12419 = _GEN_19588 | _GEN_5761; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12420 = _GEN_19589 | _GEN_5762; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12421 = _GEN_19590 | _GEN_5763; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12422 = _GEN_19591 | _GEN_5764; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12423 = _GEN_19592 | _GEN_5765; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12424 = _GEN_19593 | _GEN_5766; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12425 = _GEN_19594 | _GEN_5767; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12426 = _GEN_19595 | _GEN_5768; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12427 = _GEN_19596 | _GEN_5769; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12428 = _GEN_19597 | _GEN_5770; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12429 = _GEN_19598 | _GEN_5771; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12430 = _GEN_19599 | _GEN_5772; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12431 = _GEN_19600 | _GEN_5773; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12432 = _GEN_19601 | _GEN_5774; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12433 = _GEN_19602 | _GEN_5775; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12434 = _GEN_19603 | _GEN_5776; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12435 = _GEN_19604 | _GEN_5777; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12436 = _GEN_19605 | _GEN_5778; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12437 = _GEN_19606 | _GEN_5779; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12438 = _GEN_19607 | _GEN_5780; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12439 = _GEN_19608 | _GEN_5781; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12440 = _GEN_19609 | _GEN_5782; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12441 = _GEN_19610 | _GEN_5783; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12442 = _GEN_19611 | _GEN_5784; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12443 = _GEN_19612 | _GEN_5785; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12444 = _GEN_19613 | _GEN_5786; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12445 = _GEN_19614 | _GEN_5787; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12446 = _GEN_19615 | _GEN_5788; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12447 = _GEN_19616 | _GEN_5789; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12448 = _GEN_19617 | _GEN_5790; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12449 = _GEN_19618 | _GEN_5791; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12450 = _GEN_19619 | _GEN_5792; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12451 = _GEN_19620 | _GEN_5793; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12452 = _GEN_19621 | _GEN_5794; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12453 = _GEN_19622 | _GEN_5795; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12454 = _GEN_19623 | _GEN_5796; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12455 = _GEN_19624 | _GEN_5797; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12456 = _GEN_19625 | _GEN_5798; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12457 = _GEN_19626 | _GEN_5799; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12458 = _GEN_19627 | _GEN_5800; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12459 = _GEN_19628 | _GEN_5801; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12460 = _GEN_19629 | _GEN_5802; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12461 = _GEN_19630 | _GEN_5803; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12462 = _GEN_19631 | _GEN_5804; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12463 = _GEN_19632 | _GEN_5805; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12464 = _GEN_19633 | _GEN_5806; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12465 = _GEN_19634 | _GEN_5807; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12466 = _GEN_19635 | _GEN_5808; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12467 = _GEN_19636 | _GEN_5809; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12468 = _GEN_19637 | _GEN_5810; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12469 = _GEN_19638 | _GEN_5811; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12470 = _GEN_19639 | _GEN_5812; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12471 = _GEN_19640 | _GEN_5813; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12472 = _GEN_19641 | _GEN_5814; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12473 = _GEN_19642 | _GEN_5815; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12474 = _GEN_19643 | _GEN_5816; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12475 = _GEN_19644 | _GEN_5817; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12476 = _GEN_19645 | _GEN_5818; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12477 = _GEN_19646 | _GEN_5819; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12478 = _GEN_19647 | _GEN_5820; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12479 = _GEN_19648 | _GEN_5821; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12480 = _GEN_19649 | _GEN_5822; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12481 = _GEN_19650 | _GEN_5823; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12482 = _GEN_19651 | _GEN_5824; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12483 = _GEN_19652 | _GEN_5825; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12484 = _GEN_19653 | _GEN_5826; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12485 = _GEN_19654 | _GEN_5827; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12486 = _GEN_19655 | _GEN_5828; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12487 = _GEN_19656 | _GEN_5829; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12488 = _GEN_19657 | _GEN_5830; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12489 = _GEN_19658 | _GEN_5831; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12490 = _GEN_19659 | _GEN_5832; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12491 = _GEN_19660 | _GEN_5833; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12492 = _GEN_19661 | _GEN_5834; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12493 = _GEN_19662 | _GEN_5835; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12494 = _GEN_19663 | _GEN_5836; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12495 = _GEN_19664 | _GEN_5837; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12496 = _GEN_19665 | _GEN_5838; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12497 = _GEN_19666 | _GEN_5839; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12498 = _GEN_19667 | _GEN_5840; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12499 = _GEN_19668 | _GEN_5841; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12500 = _GEN_19669 | _GEN_5842; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12501 = _GEN_19670 | _GEN_5843; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12502 = _GEN_19671 | _GEN_5844; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12503 = _GEN_19672 | _GEN_5845; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12504 = _GEN_19673 | _GEN_5846; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12505 = _GEN_19674 | _GEN_5847; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12506 = _GEN_19675 | _GEN_5848; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12507 = _GEN_19676 | _GEN_5849; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12508 = _GEN_19677 | _GEN_5850; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12509 = _GEN_19678 | _GEN_5851; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12510 = _GEN_19679 | _GEN_5852; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12511 = _GEN_19680 | _GEN_5853; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12512 = _GEN_19681 | _GEN_5854; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12513 = _GEN_19682 | _GEN_5855; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12514 = _GEN_19683 | _GEN_5856; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12515 = _GEN_19684 | _GEN_5857; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12516 = _GEN_19685 | _GEN_5858; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12517 = _GEN_19686 | _GEN_5859; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12518 = _GEN_19687 | _GEN_5860; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12519 = _GEN_19688 | _GEN_5861; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12520 = _GEN_19689 | _GEN_5862; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12521 = _GEN_19690 | _GEN_5863; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12522 = _GEN_19691 | _GEN_5864; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12523 = _GEN_19692 | _GEN_5865; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12524 = _GEN_19693 | _GEN_5866; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12525 = _GEN_19694 | _GEN_5867; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12526 = _GEN_19695 | _GEN_5868; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12527 = _GEN_19696 | _GEN_5869; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12528 = _GEN_19697 | _GEN_5870; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12529 = _GEN_19698 | _GEN_5871; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12530 = _GEN_19699 | _GEN_5872; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12531 = _GEN_19700 | _GEN_5873; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12532 = _GEN_19701 | _GEN_5874; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12533 = _GEN_19702 | _GEN_5875; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12534 = _GEN_19703 | _GEN_5876; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12535 = _GEN_19704 | _GEN_5877; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12536 = _GEN_19705 | _GEN_5878; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12537 = _GEN_19706 | _GEN_5879; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12538 = _GEN_19707 | _GEN_5880; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12539 = _GEN_19708 | _GEN_5881; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12540 = _GEN_19709 | _GEN_5882; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12541 = _GEN_19710 | _GEN_5883; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12542 = _GEN_19711 | _GEN_5884; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12543 = _GEN_19712 | _GEN_5885; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12544 = _GEN_19713 | _GEN_5886; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12545 = _GEN_19714 | _GEN_5887; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12546 = _GEN_19715 | _GEN_5888; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12547 = _GEN_19716 | _GEN_5889; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12548 = _GEN_19717 | _GEN_5890; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12549 = _GEN_19718 | _GEN_5891; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12550 = _GEN_19719 | _GEN_5892; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12551 = _GEN_19720 | _GEN_5893; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12552 = _GEN_19721 | _GEN_5894; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12553 = _GEN_19722 | _GEN_5895; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12554 = _GEN_19723 | _GEN_5896; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12555 = _GEN_19724 | _GEN_5897; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12556 = _GEN_19725 | _GEN_5898; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12557 = _GEN_19726 | _GEN_5899; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12558 = _GEN_19727 | _GEN_5900; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12559 = _GEN_19728 | _GEN_5901; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12560 = _GEN_19729 | _GEN_5902; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12561 = _GEN_19730 | _GEN_5903; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12562 = _GEN_19731 | _GEN_5904; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12563 = _GEN_19732 | _GEN_5905; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12564 = _GEN_19733 | _GEN_5906; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12565 = _GEN_19734 | _GEN_5907; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12566 = _GEN_19735 | _GEN_5908; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12567 = _GEN_19736 | _GEN_5909; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12568 = _GEN_19737 | _GEN_5910; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12569 = _GEN_19738 | _GEN_5911; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12570 = _GEN_19739 | _GEN_5912; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12571 = _GEN_19740 | _GEN_5913; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12572 = _GEN_19741 | _GEN_5914; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12573 = _GEN_19742 | _GEN_5915; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12574 = _GEN_19743 | _GEN_5916; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12575 = _GEN_19744 | _GEN_5917; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12576 = _GEN_19745 | _GEN_5918; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12577 = _GEN_19746 | _GEN_5919; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12578 = _GEN_19747 | _GEN_5920; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12579 = _GEN_19748 | _GEN_5921; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12580 = _GEN_19749 | _GEN_5922; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12581 = _GEN_19750 | _GEN_5923; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12582 = _GEN_19751 | _GEN_5924; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12583 = _GEN_19752 | _GEN_5925; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12584 = _GEN_19753 | _GEN_5926; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12585 = _GEN_19754 | _GEN_5927; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12586 = _GEN_19755 | _GEN_5928; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12587 = _GEN_19756 | _GEN_5929; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12588 = _GEN_19757 | _GEN_5930; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12589 = _GEN_19758 | _GEN_5931; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12590 = _GEN_19759 | _GEN_5932; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12591 = _GEN_19760 | _GEN_5933; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12592 = _GEN_19761 | _GEN_5934; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12593 = _GEN_19762 | _GEN_5935; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12594 = _GEN_19763 | _GEN_5936; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12595 = _GEN_19764 | _GEN_5937; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12596 = _GEN_19765 | _GEN_5938; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12597 = _GEN_19766 | _GEN_5939; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12598 = _GEN_19767 | _GEN_5940; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12599 = _GEN_19768 | _GEN_5941; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12600 = _GEN_19769 | _GEN_5942; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12601 = _GEN_19770 | _GEN_5943; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12602 = _GEN_19771 | _GEN_5944; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12603 = _GEN_19772 | _GEN_5945; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12604 = _GEN_19773 | _GEN_5946; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12605 = _GEN_19774 | _GEN_5947; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12606 = _GEN_19775 | _GEN_5948; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12607 = _GEN_19776 | _GEN_5949; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12608 = _GEN_19777 | _GEN_5950; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12609 = _GEN_19778 | _GEN_5951; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12610 = _GEN_19779 | _GEN_5952; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12611 = _GEN_19780 | _GEN_5953; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12612 = _GEN_19781 | _GEN_5954; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12613 = _GEN_19782 | _GEN_5955; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12614 = _GEN_19783 | _GEN_5956; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12615 = _GEN_19784 | _GEN_5957; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12616 = _GEN_19785 | _GEN_5958; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12617 = _GEN_19786 | _GEN_5959; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12618 = _GEN_19787 | _GEN_5960; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12619 = _GEN_19788 | _GEN_5961; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12620 = _GEN_19789 | _GEN_5962; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12621 = _GEN_19790 | _GEN_5963; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12622 = _GEN_19791 | _GEN_5964; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12623 = _GEN_19792 | _GEN_5965; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12624 = _GEN_19793 | _GEN_5966; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12625 = _GEN_19794 | _GEN_5967; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12626 = _GEN_19795 | _GEN_5968; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12627 = _GEN_19796 | _GEN_5969; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12628 = _GEN_19797 | _GEN_5970; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12629 = _GEN_19798 | _GEN_5971; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12630 = _GEN_19799 | _GEN_5972; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12631 = _GEN_19800 | _GEN_5973; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12632 = _GEN_19801 | _GEN_5974; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12633 = _GEN_19802 | _GEN_5975; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12634 = _GEN_19803 | _GEN_5976; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12635 = _GEN_19804 | _GEN_5977; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12636 = _GEN_19805 | _GEN_5978; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12637 = _GEN_19806 | _GEN_5979; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12638 = _GEN_19807 | _GEN_5980; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12639 = _GEN_19808 | _GEN_5981; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12640 = _GEN_19809 | _GEN_5982; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12641 = _GEN_19810 | _GEN_5983; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12642 = _GEN_19811 | _GEN_5984; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12643 = _GEN_19812 | _GEN_5985; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12644 = _GEN_19813 | _GEN_5986; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12645 = _GEN_19814 | _GEN_5987; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12646 = _GEN_19815 | _GEN_5988; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12647 = _GEN_19816 | _GEN_5989; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12648 = _GEN_19817 | _GEN_5990; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12649 = _GEN_19818 | _GEN_5991; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12650 = _GEN_19819 | _GEN_5992; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12651 = _GEN_19820 | _GEN_5993; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12652 = _GEN_19821 | _GEN_5994; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12653 = _GEN_19822 | _GEN_5995; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12654 = _GEN_19823 | _GEN_5996; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12655 = _GEN_19824 | _GEN_5997; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12656 = _GEN_19825 | _GEN_5998; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12657 = _GEN_19826 | _GEN_5999; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12658 = _GEN_19827 | _GEN_6000; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12659 = _GEN_19828 | _GEN_6001; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12660 = _GEN_19829 | _GEN_6002; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12661 = _GEN_19830 | _GEN_6003; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12662 = _GEN_19831 | _GEN_6004; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12663 = _GEN_19832 | _GEN_6005; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12664 = _GEN_19833 | _GEN_6006; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12665 = _GEN_19834 | _GEN_6007; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12666 = _GEN_19835 | _GEN_6008; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12667 = _GEN_19836 | _GEN_6009; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12668 = _GEN_19837 | _GEN_6010; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12669 = _GEN_19838 | _GEN_6011; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12670 = _GEN_19839 | _GEN_6012; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12671 = _GEN_19840 | _GEN_6013; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12672 = _GEN_19841 | _GEN_6014; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12673 = _GEN_19842 | _GEN_6015; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12674 = _GEN_19843 | _GEN_6016; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12675 = _GEN_19844 | _GEN_6017; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12676 = _GEN_19845 | _GEN_6018; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12677 = _GEN_19846 | _GEN_6019; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12678 = _GEN_19847 | _GEN_6020; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12679 = _GEN_19848 | _GEN_6021; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12680 = _GEN_19849 | _GEN_6022; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12681 = _GEN_19850 | _GEN_6023; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12682 = _GEN_19851 | _GEN_6024; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12683 = _GEN_19852 | _GEN_6025; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12684 = _GEN_19853 | _GEN_6026; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12685 = _GEN_19854 | _GEN_6027; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12686 = _GEN_19855 | _GEN_6028; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12687 = _GEN_19856 | _GEN_6029; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12688 = _GEN_19857 | _GEN_6030; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12689 = _GEN_19858 | _GEN_6031; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12690 = _GEN_19859 | _GEN_6032; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12691 = _GEN_19860 | _GEN_6033; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12692 = _GEN_19861 | _GEN_6034; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12693 = _GEN_19862 | _GEN_6035; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12694 = _GEN_19863 | _GEN_6036; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12695 = _GEN_19864 | _GEN_6037; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12696 = _GEN_19865 | _GEN_6038; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12697 = _GEN_19866 | _GEN_6039; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12698 = _GEN_19867 | _GEN_6040; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12699 = _GEN_19868 | _GEN_6041; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12700 = _GEN_19869 | _GEN_6042; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12701 = _GEN_19870 | _GEN_6043; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12702 = _GEN_19871 | _GEN_6044; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12703 = _GEN_19872 | _GEN_6045; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12704 = _GEN_19873 | _GEN_6046; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12705 = _GEN_19874 | _GEN_6047; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12706 = _GEN_19875 | _GEN_6048; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12707 = _GEN_19876 | _GEN_6049; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12708 = _GEN_19877 | _GEN_6050; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12709 = _GEN_19878 | _GEN_6051; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12710 = _GEN_19879 | _GEN_6052; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12711 = _GEN_19880 | _GEN_6053; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12712 = _GEN_19881 | _GEN_6054; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12713 = _GEN_19882 | _GEN_6055; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12714 = _GEN_19883 | _GEN_6056; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12715 = _GEN_19884 | _GEN_6057; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12716 = _GEN_19885 | _GEN_6058; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12717 = _GEN_19886 | _GEN_6059; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12718 = _GEN_19887 | _GEN_6060; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12719 = _GEN_19888 | _GEN_6061; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12720 = _GEN_19889 | _GEN_6062; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12721 = _GEN_19890 | _GEN_6063; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12722 = _GEN_19891 | _GEN_6064; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12723 = _GEN_19892 | _GEN_6065; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12724 = _GEN_19893 | _GEN_6066; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12725 = _GEN_19894 | _GEN_6067; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12726 = _GEN_19895 | _GEN_6068; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12727 = _GEN_19896 | _GEN_6069; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12728 = _GEN_19897 | _GEN_6070; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12729 = _GEN_19898 | _GEN_6071; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12730 = _GEN_19899 | _GEN_6072; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12731 = _GEN_19900 | _GEN_6073; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12732 = _GEN_19901 | _GEN_6074; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12733 = _GEN_19902 | _GEN_6075; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12734 = _GEN_19903 | _GEN_6076; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12735 = _GEN_19904 | _GEN_6077; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12736 = _GEN_19905 | _GEN_6078; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12737 = _GEN_19906 | _GEN_6079; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12738 = _GEN_19907 | _GEN_6080; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12739 = _GEN_19908 | _GEN_6081; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12740 = _GEN_19909 | _GEN_6082; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12741 = _GEN_19910 | _GEN_6083; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12742 = _GEN_19911 | _GEN_6084; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12743 = _GEN_19912 | _GEN_6085; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12744 = _GEN_19913 | _GEN_6086; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12745 = _GEN_19914 | _GEN_6087; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12746 = _GEN_19915 | _GEN_6088; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12747 = _GEN_19916 | _GEN_6089; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12748 = _GEN_19917 | _GEN_6090; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12749 = _GEN_19918 | _GEN_6091; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12750 = _GEN_19919 | _GEN_6092; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12751 = _GEN_19920 | _GEN_6093; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12752 = _GEN_19921 | _GEN_6094; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12753 = _GEN_19922 | _GEN_6095; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12754 = _GEN_19923 | _GEN_6096; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12755 = _GEN_19924 | _GEN_6097; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12756 = _GEN_19925 | _GEN_6098; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12757 = _GEN_19926 | _GEN_6099; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12758 = _GEN_19927 | _GEN_6100; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12759 = _GEN_19928 | _GEN_6101; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12760 = _GEN_19929 | _GEN_6102; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12761 = _GEN_19930 | _GEN_6103; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12762 = _GEN_19931 | _GEN_6104; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12763 = _GEN_19932 | _GEN_6105; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12764 = _GEN_19933 | _GEN_6106; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12765 = _GEN_19934 | _GEN_6107; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12766 = _GEN_19935 | _GEN_6108; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12767 = _GEN_19936 | _GEN_6109; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12768 = _GEN_19937 | _GEN_6110; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12769 = _GEN_19938 | _GEN_6111; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12770 = _GEN_19939 | _GEN_6112; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12771 = _GEN_19940 | _GEN_6113; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12772 = _GEN_19941 | _GEN_6114; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12773 = _GEN_19942 | _GEN_6115; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12774 = _GEN_19943 | _GEN_6116; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12775 = _GEN_19944 | _GEN_6117; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12776 = _GEN_19945 | _GEN_6118; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12777 = _GEN_19946 | _GEN_6119; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12778 = _GEN_19947 | _GEN_6120; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12779 = _GEN_19948 | _GEN_6121; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12780 = _GEN_19949 | _GEN_6122; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12781 = _GEN_19950 | _GEN_6123; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12782 = _GEN_19951 | _GEN_6124; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12783 = _GEN_19952 | _GEN_6125; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12784 = _GEN_19953 | _GEN_6126; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12785 = _GEN_19954 | _GEN_6127; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12786 = _GEN_19955 | _GEN_6128; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12787 = _GEN_19956 | _GEN_6129; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12788 = _GEN_19957 | _GEN_6130; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12789 = _GEN_19958 | _GEN_6131; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12790 = _GEN_19959 | _GEN_6132; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12791 = _GEN_19960 | _GEN_6133; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12792 = _GEN_19961 | _GEN_6134; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12793 = _GEN_19962 | _GEN_6135; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12794 = _GEN_19963 | _GEN_6136; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12795 = _GEN_19964 | _GEN_6137; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12796 = _GEN_19965 | _GEN_6138; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12797 = _GEN_19966 | _GEN_6139; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12798 = _GEN_19967 | _GEN_6140; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12799 = _GEN_19968 | _GEN_6141; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12800 = _GEN_19969 | _GEN_6142; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_12801 = _GEN_19970 | _GEN_6143; // @[branch_predictor.scala 99:{35,35}]
  wire  _GEN_15362 = _T_1027 & ~entry_found ? _GEN_12290 : _GEN_5632; // @[branch_predictor.scala 98:103]
  wire  _GEN_15363 = _T_1027 & ~entry_found ? _GEN_12291 : _GEN_5633; // @[branch_predictor.scala 98:103]
  wire  _GEN_15364 = _T_1027 & ~entry_found ? _GEN_12292 : _GEN_5634; // @[branch_predictor.scala 98:103]
  wire  _GEN_15365 = _T_1027 & ~entry_found ? _GEN_12293 : _GEN_5635; // @[branch_predictor.scala 98:103]
  wire  _GEN_15366 = _T_1027 & ~entry_found ? _GEN_12294 : _GEN_5636; // @[branch_predictor.scala 98:103]
  wire  _GEN_15367 = _T_1027 & ~entry_found ? _GEN_12295 : _GEN_5637; // @[branch_predictor.scala 98:103]
  wire  _GEN_15368 = _T_1027 & ~entry_found ? _GEN_12296 : _GEN_5638; // @[branch_predictor.scala 98:103]
  wire  _GEN_15369 = _T_1027 & ~entry_found ? _GEN_12297 : _GEN_5639; // @[branch_predictor.scala 98:103]
  wire  _GEN_15370 = _T_1027 & ~entry_found ? _GEN_12298 : _GEN_5640; // @[branch_predictor.scala 98:103]
  wire  _GEN_15371 = _T_1027 & ~entry_found ? _GEN_12299 : _GEN_5641; // @[branch_predictor.scala 98:103]
  wire  _GEN_15372 = _T_1027 & ~entry_found ? _GEN_12300 : _GEN_5642; // @[branch_predictor.scala 98:103]
  wire  _GEN_15373 = _T_1027 & ~entry_found ? _GEN_12301 : _GEN_5643; // @[branch_predictor.scala 98:103]
  wire  _GEN_15374 = _T_1027 & ~entry_found ? _GEN_12302 : _GEN_5644; // @[branch_predictor.scala 98:103]
  wire  _GEN_15375 = _T_1027 & ~entry_found ? _GEN_12303 : _GEN_5645; // @[branch_predictor.scala 98:103]
  wire  _GEN_15376 = _T_1027 & ~entry_found ? _GEN_12304 : _GEN_5646; // @[branch_predictor.scala 98:103]
  wire  _GEN_15377 = _T_1027 & ~entry_found ? _GEN_12305 : _GEN_5647; // @[branch_predictor.scala 98:103]
  wire  _GEN_15378 = _T_1027 & ~entry_found ? _GEN_12306 : _GEN_5648; // @[branch_predictor.scala 98:103]
  wire  _GEN_15379 = _T_1027 & ~entry_found ? _GEN_12307 : _GEN_5649; // @[branch_predictor.scala 98:103]
  wire  _GEN_15380 = _T_1027 & ~entry_found ? _GEN_12308 : _GEN_5650; // @[branch_predictor.scala 98:103]
  wire  _GEN_15381 = _T_1027 & ~entry_found ? _GEN_12309 : _GEN_5651; // @[branch_predictor.scala 98:103]
  wire  _GEN_15382 = _T_1027 & ~entry_found ? _GEN_12310 : _GEN_5652; // @[branch_predictor.scala 98:103]
  wire  _GEN_15383 = _T_1027 & ~entry_found ? _GEN_12311 : _GEN_5653; // @[branch_predictor.scala 98:103]
  wire  _GEN_15384 = _T_1027 & ~entry_found ? _GEN_12312 : _GEN_5654; // @[branch_predictor.scala 98:103]
  wire  _GEN_15385 = _T_1027 & ~entry_found ? _GEN_12313 : _GEN_5655; // @[branch_predictor.scala 98:103]
  wire  _GEN_15386 = _T_1027 & ~entry_found ? _GEN_12314 : _GEN_5656; // @[branch_predictor.scala 98:103]
  wire  _GEN_15387 = _T_1027 & ~entry_found ? _GEN_12315 : _GEN_5657; // @[branch_predictor.scala 98:103]
  wire  _GEN_15388 = _T_1027 & ~entry_found ? _GEN_12316 : _GEN_5658; // @[branch_predictor.scala 98:103]
  wire  _GEN_15389 = _T_1027 & ~entry_found ? _GEN_12317 : _GEN_5659; // @[branch_predictor.scala 98:103]
  wire  _GEN_15390 = _T_1027 & ~entry_found ? _GEN_12318 : _GEN_5660; // @[branch_predictor.scala 98:103]
  wire  _GEN_15391 = _T_1027 & ~entry_found ? _GEN_12319 : _GEN_5661; // @[branch_predictor.scala 98:103]
  wire  _GEN_15392 = _T_1027 & ~entry_found ? _GEN_12320 : _GEN_5662; // @[branch_predictor.scala 98:103]
  wire  _GEN_15393 = _T_1027 & ~entry_found ? _GEN_12321 : _GEN_5663; // @[branch_predictor.scala 98:103]
  wire  _GEN_15394 = _T_1027 & ~entry_found ? _GEN_12322 : _GEN_5664; // @[branch_predictor.scala 98:103]
  wire  _GEN_15395 = _T_1027 & ~entry_found ? _GEN_12323 : _GEN_5665; // @[branch_predictor.scala 98:103]
  wire  _GEN_15396 = _T_1027 & ~entry_found ? _GEN_12324 : _GEN_5666; // @[branch_predictor.scala 98:103]
  wire  _GEN_15397 = _T_1027 & ~entry_found ? _GEN_12325 : _GEN_5667; // @[branch_predictor.scala 98:103]
  wire  _GEN_15398 = _T_1027 & ~entry_found ? _GEN_12326 : _GEN_5668; // @[branch_predictor.scala 98:103]
  wire  _GEN_15399 = _T_1027 & ~entry_found ? _GEN_12327 : _GEN_5669; // @[branch_predictor.scala 98:103]
  wire  _GEN_15400 = _T_1027 & ~entry_found ? _GEN_12328 : _GEN_5670; // @[branch_predictor.scala 98:103]
  wire  _GEN_15401 = _T_1027 & ~entry_found ? _GEN_12329 : _GEN_5671; // @[branch_predictor.scala 98:103]
  wire  _GEN_15402 = _T_1027 & ~entry_found ? _GEN_12330 : _GEN_5672; // @[branch_predictor.scala 98:103]
  wire  _GEN_15403 = _T_1027 & ~entry_found ? _GEN_12331 : _GEN_5673; // @[branch_predictor.scala 98:103]
  wire  _GEN_15404 = _T_1027 & ~entry_found ? _GEN_12332 : _GEN_5674; // @[branch_predictor.scala 98:103]
  wire  _GEN_15405 = _T_1027 & ~entry_found ? _GEN_12333 : _GEN_5675; // @[branch_predictor.scala 98:103]
  wire  _GEN_15406 = _T_1027 & ~entry_found ? _GEN_12334 : _GEN_5676; // @[branch_predictor.scala 98:103]
  wire  _GEN_15407 = _T_1027 & ~entry_found ? _GEN_12335 : _GEN_5677; // @[branch_predictor.scala 98:103]
  wire  _GEN_15408 = _T_1027 & ~entry_found ? _GEN_12336 : _GEN_5678; // @[branch_predictor.scala 98:103]
  wire  _GEN_15409 = _T_1027 & ~entry_found ? _GEN_12337 : _GEN_5679; // @[branch_predictor.scala 98:103]
  wire  _GEN_15410 = _T_1027 & ~entry_found ? _GEN_12338 : _GEN_5680; // @[branch_predictor.scala 98:103]
  wire  _GEN_15411 = _T_1027 & ~entry_found ? _GEN_12339 : _GEN_5681; // @[branch_predictor.scala 98:103]
  wire  _GEN_15412 = _T_1027 & ~entry_found ? _GEN_12340 : _GEN_5682; // @[branch_predictor.scala 98:103]
  wire  _GEN_15413 = _T_1027 & ~entry_found ? _GEN_12341 : _GEN_5683; // @[branch_predictor.scala 98:103]
  wire  _GEN_15414 = _T_1027 & ~entry_found ? _GEN_12342 : _GEN_5684; // @[branch_predictor.scala 98:103]
  wire  _GEN_15415 = _T_1027 & ~entry_found ? _GEN_12343 : _GEN_5685; // @[branch_predictor.scala 98:103]
  wire  _GEN_15416 = _T_1027 & ~entry_found ? _GEN_12344 : _GEN_5686; // @[branch_predictor.scala 98:103]
  wire  _GEN_15417 = _T_1027 & ~entry_found ? _GEN_12345 : _GEN_5687; // @[branch_predictor.scala 98:103]
  wire  _GEN_15418 = _T_1027 & ~entry_found ? _GEN_12346 : _GEN_5688; // @[branch_predictor.scala 98:103]
  wire  _GEN_15419 = _T_1027 & ~entry_found ? _GEN_12347 : _GEN_5689; // @[branch_predictor.scala 98:103]
  wire  _GEN_15420 = _T_1027 & ~entry_found ? _GEN_12348 : _GEN_5690; // @[branch_predictor.scala 98:103]
  wire  _GEN_15421 = _T_1027 & ~entry_found ? _GEN_12349 : _GEN_5691; // @[branch_predictor.scala 98:103]
  wire  _GEN_15422 = _T_1027 & ~entry_found ? _GEN_12350 : _GEN_5692; // @[branch_predictor.scala 98:103]
  wire  _GEN_15423 = _T_1027 & ~entry_found ? _GEN_12351 : _GEN_5693; // @[branch_predictor.scala 98:103]
  wire  _GEN_15424 = _T_1027 & ~entry_found ? _GEN_12352 : _GEN_5694; // @[branch_predictor.scala 98:103]
  wire  _GEN_15425 = _T_1027 & ~entry_found ? _GEN_12353 : _GEN_5695; // @[branch_predictor.scala 98:103]
  wire  _GEN_15426 = _T_1027 & ~entry_found ? _GEN_12354 : _GEN_5696; // @[branch_predictor.scala 98:103]
  wire  _GEN_15427 = _T_1027 & ~entry_found ? _GEN_12355 : _GEN_5697; // @[branch_predictor.scala 98:103]
  wire  _GEN_15428 = _T_1027 & ~entry_found ? _GEN_12356 : _GEN_5698; // @[branch_predictor.scala 98:103]
  wire  _GEN_15429 = _T_1027 & ~entry_found ? _GEN_12357 : _GEN_5699; // @[branch_predictor.scala 98:103]
  wire  _GEN_15430 = _T_1027 & ~entry_found ? _GEN_12358 : _GEN_5700; // @[branch_predictor.scala 98:103]
  wire  _GEN_15431 = _T_1027 & ~entry_found ? _GEN_12359 : _GEN_5701; // @[branch_predictor.scala 98:103]
  wire  _GEN_15432 = _T_1027 & ~entry_found ? _GEN_12360 : _GEN_5702; // @[branch_predictor.scala 98:103]
  wire  _GEN_15433 = _T_1027 & ~entry_found ? _GEN_12361 : _GEN_5703; // @[branch_predictor.scala 98:103]
  wire  _GEN_15434 = _T_1027 & ~entry_found ? _GEN_12362 : _GEN_5704; // @[branch_predictor.scala 98:103]
  wire  _GEN_15435 = _T_1027 & ~entry_found ? _GEN_12363 : _GEN_5705; // @[branch_predictor.scala 98:103]
  wire  _GEN_15436 = _T_1027 & ~entry_found ? _GEN_12364 : _GEN_5706; // @[branch_predictor.scala 98:103]
  wire  _GEN_15437 = _T_1027 & ~entry_found ? _GEN_12365 : _GEN_5707; // @[branch_predictor.scala 98:103]
  wire  _GEN_15438 = _T_1027 & ~entry_found ? _GEN_12366 : _GEN_5708; // @[branch_predictor.scala 98:103]
  wire  _GEN_15439 = _T_1027 & ~entry_found ? _GEN_12367 : _GEN_5709; // @[branch_predictor.scala 98:103]
  wire  _GEN_15440 = _T_1027 & ~entry_found ? _GEN_12368 : _GEN_5710; // @[branch_predictor.scala 98:103]
  wire  _GEN_15441 = _T_1027 & ~entry_found ? _GEN_12369 : _GEN_5711; // @[branch_predictor.scala 98:103]
  wire  _GEN_15442 = _T_1027 & ~entry_found ? _GEN_12370 : _GEN_5712; // @[branch_predictor.scala 98:103]
  wire  _GEN_15443 = _T_1027 & ~entry_found ? _GEN_12371 : _GEN_5713; // @[branch_predictor.scala 98:103]
  wire  _GEN_15444 = _T_1027 & ~entry_found ? _GEN_12372 : _GEN_5714; // @[branch_predictor.scala 98:103]
  wire  _GEN_15445 = _T_1027 & ~entry_found ? _GEN_12373 : _GEN_5715; // @[branch_predictor.scala 98:103]
  wire  _GEN_15446 = _T_1027 & ~entry_found ? _GEN_12374 : _GEN_5716; // @[branch_predictor.scala 98:103]
  wire  _GEN_15447 = _T_1027 & ~entry_found ? _GEN_12375 : _GEN_5717; // @[branch_predictor.scala 98:103]
  wire  _GEN_15448 = _T_1027 & ~entry_found ? _GEN_12376 : _GEN_5718; // @[branch_predictor.scala 98:103]
  wire  _GEN_15449 = _T_1027 & ~entry_found ? _GEN_12377 : _GEN_5719; // @[branch_predictor.scala 98:103]
  wire  _GEN_15450 = _T_1027 & ~entry_found ? _GEN_12378 : _GEN_5720; // @[branch_predictor.scala 98:103]
  wire  _GEN_15451 = _T_1027 & ~entry_found ? _GEN_12379 : _GEN_5721; // @[branch_predictor.scala 98:103]
  wire  _GEN_15452 = _T_1027 & ~entry_found ? _GEN_12380 : _GEN_5722; // @[branch_predictor.scala 98:103]
  wire  _GEN_15453 = _T_1027 & ~entry_found ? _GEN_12381 : _GEN_5723; // @[branch_predictor.scala 98:103]
  wire  _GEN_15454 = _T_1027 & ~entry_found ? _GEN_12382 : _GEN_5724; // @[branch_predictor.scala 98:103]
  wire  _GEN_15455 = _T_1027 & ~entry_found ? _GEN_12383 : _GEN_5725; // @[branch_predictor.scala 98:103]
  wire  _GEN_15456 = _T_1027 & ~entry_found ? _GEN_12384 : _GEN_5726; // @[branch_predictor.scala 98:103]
  wire  _GEN_15457 = _T_1027 & ~entry_found ? _GEN_12385 : _GEN_5727; // @[branch_predictor.scala 98:103]
  wire  _GEN_15458 = _T_1027 & ~entry_found ? _GEN_12386 : _GEN_5728; // @[branch_predictor.scala 98:103]
  wire  _GEN_15459 = _T_1027 & ~entry_found ? _GEN_12387 : _GEN_5729; // @[branch_predictor.scala 98:103]
  wire  _GEN_15460 = _T_1027 & ~entry_found ? _GEN_12388 : _GEN_5730; // @[branch_predictor.scala 98:103]
  wire  _GEN_15461 = _T_1027 & ~entry_found ? _GEN_12389 : _GEN_5731; // @[branch_predictor.scala 98:103]
  wire  _GEN_15462 = _T_1027 & ~entry_found ? _GEN_12390 : _GEN_5732; // @[branch_predictor.scala 98:103]
  wire  _GEN_15463 = _T_1027 & ~entry_found ? _GEN_12391 : _GEN_5733; // @[branch_predictor.scala 98:103]
  wire  _GEN_15464 = _T_1027 & ~entry_found ? _GEN_12392 : _GEN_5734; // @[branch_predictor.scala 98:103]
  wire  _GEN_15465 = _T_1027 & ~entry_found ? _GEN_12393 : _GEN_5735; // @[branch_predictor.scala 98:103]
  wire  _GEN_15466 = _T_1027 & ~entry_found ? _GEN_12394 : _GEN_5736; // @[branch_predictor.scala 98:103]
  wire  _GEN_15467 = _T_1027 & ~entry_found ? _GEN_12395 : _GEN_5737; // @[branch_predictor.scala 98:103]
  wire  _GEN_15468 = _T_1027 & ~entry_found ? _GEN_12396 : _GEN_5738; // @[branch_predictor.scala 98:103]
  wire  _GEN_15469 = _T_1027 & ~entry_found ? _GEN_12397 : _GEN_5739; // @[branch_predictor.scala 98:103]
  wire  _GEN_15470 = _T_1027 & ~entry_found ? _GEN_12398 : _GEN_5740; // @[branch_predictor.scala 98:103]
  wire  _GEN_15471 = _T_1027 & ~entry_found ? _GEN_12399 : _GEN_5741; // @[branch_predictor.scala 98:103]
  wire  _GEN_15472 = _T_1027 & ~entry_found ? _GEN_12400 : _GEN_5742; // @[branch_predictor.scala 98:103]
  wire  _GEN_15473 = _T_1027 & ~entry_found ? _GEN_12401 : _GEN_5743; // @[branch_predictor.scala 98:103]
  wire  _GEN_15474 = _T_1027 & ~entry_found ? _GEN_12402 : _GEN_5744; // @[branch_predictor.scala 98:103]
  wire  _GEN_15475 = _T_1027 & ~entry_found ? _GEN_12403 : _GEN_5745; // @[branch_predictor.scala 98:103]
  wire  _GEN_15476 = _T_1027 & ~entry_found ? _GEN_12404 : _GEN_5746; // @[branch_predictor.scala 98:103]
  wire  _GEN_15477 = _T_1027 & ~entry_found ? _GEN_12405 : _GEN_5747; // @[branch_predictor.scala 98:103]
  wire  _GEN_15478 = _T_1027 & ~entry_found ? _GEN_12406 : _GEN_5748; // @[branch_predictor.scala 98:103]
  wire  _GEN_15479 = _T_1027 & ~entry_found ? _GEN_12407 : _GEN_5749; // @[branch_predictor.scala 98:103]
  wire  _GEN_15480 = _T_1027 & ~entry_found ? _GEN_12408 : _GEN_5750; // @[branch_predictor.scala 98:103]
  wire  _GEN_15481 = _T_1027 & ~entry_found ? _GEN_12409 : _GEN_5751; // @[branch_predictor.scala 98:103]
  wire  _GEN_15482 = _T_1027 & ~entry_found ? _GEN_12410 : _GEN_5752; // @[branch_predictor.scala 98:103]
  wire  _GEN_15483 = _T_1027 & ~entry_found ? _GEN_12411 : _GEN_5753; // @[branch_predictor.scala 98:103]
  wire  _GEN_15484 = _T_1027 & ~entry_found ? _GEN_12412 : _GEN_5754; // @[branch_predictor.scala 98:103]
  wire  _GEN_15485 = _T_1027 & ~entry_found ? _GEN_12413 : _GEN_5755; // @[branch_predictor.scala 98:103]
  wire  _GEN_15486 = _T_1027 & ~entry_found ? _GEN_12414 : _GEN_5756; // @[branch_predictor.scala 98:103]
  wire  _GEN_15487 = _T_1027 & ~entry_found ? _GEN_12415 : _GEN_5757; // @[branch_predictor.scala 98:103]
  wire  _GEN_15488 = _T_1027 & ~entry_found ? _GEN_12416 : _GEN_5758; // @[branch_predictor.scala 98:103]
  wire  _GEN_15489 = _T_1027 & ~entry_found ? _GEN_12417 : _GEN_5759; // @[branch_predictor.scala 98:103]
  wire  _GEN_15490 = _T_1027 & ~entry_found ? _GEN_12418 : _GEN_5760; // @[branch_predictor.scala 98:103]
  wire  _GEN_15491 = _T_1027 & ~entry_found ? _GEN_12419 : _GEN_5761; // @[branch_predictor.scala 98:103]
  wire  _GEN_15492 = _T_1027 & ~entry_found ? _GEN_12420 : _GEN_5762; // @[branch_predictor.scala 98:103]
  wire  _GEN_15493 = _T_1027 & ~entry_found ? _GEN_12421 : _GEN_5763; // @[branch_predictor.scala 98:103]
  wire  _GEN_15494 = _T_1027 & ~entry_found ? _GEN_12422 : _GEN_5764; // @[branch_predictor.scala 98:103]
  wire  _GEN_15495 = _T_1027 & ~entry_found ? _GEN_12423 : _GEN_5765; // @[branch_predictor.scala 98:103]
  wire  _GEN_15496 = _T_1027 & ~entry_found ? _GEN_12424 : _GEN_5766; // @[branch_predictor.scala 98:103]
  wire  _GEN_15497 = _T_1027 & ~entry_found ? _GEN_12425 : _GEN_5767; // @[branch_predictor.scala 98:103]
  wire  _GEN_15498 = _T_1027 & ~entry_found ? _GEN_12426 : _GEN_5768; // @[branch_predictor.scala 98:103]
  wire  _GEN_15499 = _T_1027 & ~entry_found ? _GEN_12427 : _GEN_5769; // @[branch_predictor.scala 98:103]
  wire  _GEN_15500 = _T_1027 & ~entry_found ? _GEN_12428 : _GEN_5770; // @[branch_predictor.scala 98:103]
  wire  _GEN_15501 = _T_1027 & ~entry_found ? _GEN_12429 : _GEN_5771; // @[branch_predictor.scala 98:103]
  wire  _GEN_15502 = _T_1027 & ~entry_found ? _GEN_12430 : _GEN_5772; // @[branch_predictor.scala 98:103]
  wire  _GEN_15503 = _T_1027 & ~entry_found ? _GEN_12431 : _GEN_5773; // @[branch_predictor.scala 98:103]
  wire  _GEN_15504 = _T_1027 & ~entry_found ? _GEN_12432 : _GEN_5774; // @[branch_predictor.scala 98:103]
  wire  _GEN_15505 = _T_1027 & ~entry_found ? _GEN_12433 : _GEN_5775; // @[branch_predictor.scala 98:103]
  wire  _GEN_15506 = _T_1027 & ~entry_found ? _GEN_12434 : _GEN_5776; // @[branch_predictor.scala 98:103]
  wire  _GEN_15507 = _T_1027 & ~entry_found ? _GEN_12435 : _GEN_5777; // @[branch_predictor.scala 98:103]
  wire  _GEN_15508 = _T_1027 & ~entry_found ? _GEN_12436 : _GEN_5778; // @[branch_predictor.scala 98:103]
  wire  _GEN_15509 = _T_1027 & ~entry_found ? _GEN_12437 : _GEN_5779; // @[branch_predictor.scala 98:103]
  wire  _GEN_15510 = _T_1027 & ~entry_found ? _GEN_12438 : _GEN_5780; // @[branch_predictor.scala 98:103]
  wire  _GEN_15511 = _T_1027 & ~entry_found ? _GEN_12439 : _GEN_5781; // @[branch_predictor.scala 98:103]
  wire  _GEN_15512 = _T_1027 & ~entry_found ? _GEN_12440 : _GEN_5782; // @[branch_predictor.scala 98:103]
  wire  _GEN_15513 = _T_1027 & ~entry_found ? _GEN_12441 : _GEN_5783; // @[branch_predictor.scala 98:103]
  wire  _GEN_15514 = _T_1027 & ~entry_found ? _GEN_12442 : _GEN_5784; // @[branch_predictor.scala 98:103]
  wire  _GEN_15515 = _T_1027 & ~entry_found ? _GEN_12443 : _GEN_5785; // @[branch_predictor.scala 98:103]
  wire  _GEN_15516 = _T_1027 & ~entry_found ? _GEN_12444 : _GEN_5786; // @[branch_predictor.scala 98:103]
  wire  _GEN_15517 = _T_1027 & ~entry_found ? _GEN_12445 : _GEN_5787; // @[branch_predictor.scala 98:103]
  wire  _GEN_15518 = _T_1027 & ~entry_found ? _GEN_12446 : _GEN_5788; // @[branch_predictor.scala 98:103]
  wire  _GEN_15519 = _T_1027 & ~entry_found ? _GEN_12447 : _GEN_5789; // @[branch_predictor.scala 98:103]
  wire  _GEN_15520 = _T_1027 & ~entry_found ? _GEN_12448 : _GEN_5790; // @[branch_predictor.scala 98:103]
  wire  _GEN_15521 = _T_1027 & ~entry_found ? _GEN_12449 : _GEN_5791; // @[branch_predictor.scala 98:103]
  wire  _GEN_15522 = _T_1027 & ~entry_found ? _GEN_12450 : _GEN_5792; // @[branch_predictor.scala 98:103]
  wire  _GEN_15523 = _T_1027 & ~entry_found ? _GEN_12451 : _GEN_5793; // @[branch_predictor.scala 98:103]
  wire  _GEN_15524 = _T_1027 & ~entry_found ? _GEN_12452 : _GEN_5794; // @[branch_predictor.scala 98:103]
  wire  _GEN_15525 = _T_1027 & ~entry_found ? _GEN_12453 : _GEN_5795; // @[branch_predictor.scala 98:103]
  wire  _GEN_15526 = _T_1027 & ~entry_found ? _GEN_12454 : _GEN_5796; // @[branch_predictor.scala 98:103]
  wire  _GEN_15527 = _T_1027 & ~entry_found ? _GEN_12455 : _GEN_5797; // @[branch_predictor.scala 98:103]
  wire  _GEN_15528 = _T_1027 & ~entry_found ? _GEN_12456 : _GEN_5798; // @[branch_predictor.scala 98:103]
  wire  _GEN_15529 = _T_1027 & ~entry_found ? _GEN_12457 : _GEN_5799; // @[branch_predictor.scala 98:103]
  wire  _GEN_15530 = _T_1027 & ~entry_found ? _GEN_12458 : _GEN_5800; // @[branch_predictor.scala 98:103]
  wire  _GEN_15531 = _T_1027 & ~entry_found ? _GEN_12459 : _GEN_5801; // @[branch_predictor.scala 98:103]
  wire  _GEN_15532 = _T_1027 & ~entry_found ? _GEN_12460 : _GEN_5802; // @[branch_predictor.scala 98:103]
  wire  _GEN_15533 = _T_1027 & ~entry_found ? _GEN_12461 : _GEN_5803; // @[branch_predictor.scala 98:103]
  wire  _GEN_15534 = _T_1027 & ~entry_found ? _GEN_12462 : _GEN_5804; // @[branch_predictor.scala 98:103]
  wire  _GEN_15535 = _T_1027 & ~entry_found ? _GEN_12463 : _GEN_5805; // @[branch_predictor.scala 98:103]
  wire  _GEN_15536 = _T_1027 & ~entry_found ? _GEN_12464 : _GEN_5806; // @[branch_predictor.scala 98:103]
  wire  _GEN_15537 = _T_1027 & ~entry_found ? _GEN_12465 : _GEN_5807; // @[branch_predictor.scala 98:103]
  wire  _GEN_15538 = _T_1027 & ~entry_found ? _GEN_12466 : _GEN_5808; // @[branch_predictor.scala 98:103]
  wire  _GEN_15539 = _T_1027 & ~entry_found ? _GEN_12467 : _GEN_5809; // @[branch_predictor.scala 98:103]
  wire  _GEN_15540 = _T_1027 & ~entry_found ? _GEN_12468 : _GEN_5810; // @[branch_predictor.scala 98:103]
  wire  _GEN_15541 = _T_1027 & ~entry_found ? _GEN_12469 : _GEN_5811; // @[branch_predictor.scala 98:103]
  wire  _GEN_15542 = _T_1027 & ~entry_found ? _GEN_12470 : _GEN_5812; // @[branch_predictor.scala 98:103]
  wire  _GEN_15543 = _T_1027 & ~entry_found ? _GEN_12471 : _GEN_5813; // @[branch_predictor.scala 98:103]
  wire  _GEN_15544 = _T_1027 & ~entry_found ? _GEN_12472 : _GEN_5814; // @[branch_predictor.scala 98:103]
  wire  _GEN_15545 = _T_1027 & ~entry_found ? _GEN_12473 : _GEN_5815; // @[branch_predictor.scala 98:103]
  wire  _GEN_15546 = _T_1027 & ~entry_found ? _GEN_12474 : _GEN_5816; // @[branch_predictor.scala 98:103]
  wire  _GEN_15547 = _T_1027 & ~entry_found ? _GEN_12475 : _GEN_5817; // @[branch_predictor.scala 98:103]
  wire  _GEN_15548 = _T_1027 & ~entry_found ? _GEN_12476 : _GEN_5818; // @[branch_predictor.scala 98:103]
  wire  _GEN_15549 = _T_1027 & ~entry_found ? _GEN_12477 : _GEN_5819; // @[branch_predictor.scala 98:103]
  wire  _GEN_15550 = _T_1027 & ~entry_found ? _GEN_12478 : _GEN_5820; // @[branch_predictor.scala 98:103]
  wire  _GEN_15551 = _T_1027 & ~entry_found ? _GEN_12479 : _GEN_5821; // @[branch_predictor.scala 98:103]
  wire  _GEN_15552 = _T_1027 & ~entry_found ? _GEN_12480 : _GEN_5822; // @[branch_predictor.scala 98:103]
  wire  _GEN_15553 = _T_1027 & ~entry_found ? _GEN_12481 : _GEN_5823; // @[branch_predictor.scala 98:103]
  wire  _GEN_15554 = _T_1027 & ~entry_found ? _GEN_12482 : _GEN_5824; // @[branch_predictor.scala 98:103]
  wire  _GEN_15555 = _T_1027 & ~entry_found ? _GEN_12483 : _GEN_5825; // @[branch_predictor.scala 98:103]
  wire  _GEN_15556 = _T_1027 & ~entry_found ? _GEN_12484 : _GEN_5826; // @[branch_predictor.scala 98:103]
  wire  _GEN_15557 = _T_1027 & ~entry_found ? _GEN_12485 : _GEN_5827; // @[branch_predictor.scala 98:103]
  wire  _GEN_15558 = _T_1027 & ~entry_found ? _GEN_12486 : _GEN_5828; // @[branch_predictor.scala 98:103]
  wire  _GEN_15559 = _T_1027 & ~entry_found ? _GEN_12487 : _GEN_5829; // @[branch_predictor.scala 98:103]
  wire  _GEN_15560 = _T_1027 & ~entry_found ? _GEN_12488 : _GEN_5830; // @[branch_predictor.scala 98:103]
  wire  _GEN_15561 = _T_1027 & ~entry_found ? _GEN_12489 : _GEN_5831; // @[branch_predictor.scala 98:103]
  wire  _GEN_15562 = _T_1027 & ~entry_found ? _GEN_12490 : _GEN_5832; // @[branch_predictor.scala 98:103]
  wire  _GEN_15563 = _T_1027 & ~entry_found ? _GEN_12491 : _GEN_5833; // @[branch_predictor.scala 98:103]
  wire  _GEN_15564 = _T_1027 & ~entry_found ? _GEN_12492 : _GEN_5834; // @[branch_predictor.scala 98:103]
  wire  _GEN_15565 = _T_1027 & ~entry_found ? _GEN_12493 : _GEN_5835; // @[branch_predictor.scala 98:103]
  wire  _GEN_15566 = _T_1027 & ~entry_found ? _GEN_12494 : _GEN_5836; // @[branch_predictor.scala 98:103]
  wire  _GEN_15567 = _T_1027 & ~entry_found ? _GEN_12495 : _GEN_5837; // @[branch_predictor.scala 98:103]
  wire  _GEN_15568 = _T_1027 & ~entry_found ? _GEN_12496 : _GEN_5838; // @[branch_predictor.scala 98:103]
  wire  _GEN_15569 = _T_1027 & ~entry_found ? _GEN_12497 : _GEN_5839; // @[branch_predictor.scala 98:103]
  wire  _GEN_15570 = _T_1027 & ~entry_found ? _GEN_12498 : _GEN_5840; // @[branch_predictor.scala 98:103]
  wire  _GEN_15571 = _T_1027 & ~entry_found ? _GEN_12499 : _GEN_5841; // @[branch_predictor.scala 98:103]
  wire  _GEN_15572 = _T_1027 & ~entry_found ? _GEN_12500 : _GEN_5842; // @[branch_predictor.scala 98:103]
  wire  _GEN_15573 = _T_1027 & ~entry_found ? _GEN_12501 : _GEN_5843; // @[branch_predictor.scala 98:103]
  wire  _GEN_15574 = _T_1027 & ~entry_found ? _GEN_12502 : _GEN_5844; // @[branch_predictor.scala 98:103]
  wire  _GEN_15575 = _T_1027 & ~entry_found ? _GEN_12503 : _GEN_5845; // @[branch_predictor.scala 98:103]
  wire  _GEN_15576 = _T_1027 & ~entry_found ? _GEN_12504 : _GEN_5846; // @[branch_predictor.scala 98:103]
  wire  _GEN_15577 = _T_1027 & ~entry_found ? _GEN_12505 : _GEN_5847; // @[branch_predictor.scala 98:103]
  wire  _GEN_15578 = _T_1027 & ~entry_found ? _GEN_12506 : _GEN_5848; // @[branch_predictor.scala 98:103]
  wire  _GEN_15579 = _T_1027 & ~entry_found ? _GEN_12507 : _GEN_5849; // @[branch_predictor.scala 98:103]
  wire  _GEN_15580 = _T_1027 & ~entry_found ? _GEN_12508 : _GEN_5850; // @[branch_predictor.scala 98:103]
  wire  _GEN_15581 = _T_1027 & ~entry_found ? _GEN_12509 : _GEN_5851; // @[branch_predictor.scala 98:103]
  wire  _GEN_15582 = _T_1027 & ~entry_found ? _GEN_12510 : _GEN_5852; // @[branch_predictor.scala 98:103]
  wire  _GEN_15583 = _T_1027 & ~entry_found ? _GEN_12511 : _GEN_5853; // @[branch_predictor.scala 98:103]
  wire  _GEN_15584 = _T_1027 & ~entry_found ? _GEN_12512 : _GEN_5854; // @[branch_predictor.scala 98:103]
  wire  _GEN_15585 = _T_1027 & ~entry_found ? _GEN_12513 : _GEN_5855; // @[branch_predictor.scala 98:103]
  wire  _GEN_15586 = _T_1027 & ~entry_found ? _GEN_12514 : _GEN_5856; // @[branch_predictor.scala 98:103]
  wire  _GEN_15587 = _T_1027 & ~entry_found ? _GEN_12515 : _GEN_5857; // @[branch_predictor.scala 98:103]
  wire  _GEN_15588 = _T_1027 & ~entry_found ? _GEN_12516 : _GEN_5858; // @[branch_predictor.scala 98:103]
  wire  _GEN_15589 = _T_1027 & ~entry_found ? _GEN_12517 : _GEN_5859; // @[branch_predictor.scala 98:103]
  wire  _GEN_15590 = _T_1027 & ~entry_found ? _GEN_12518 : _GEN_5860; // @[branch_predictor.scala 98:103]
  wire  _GEN_15591 = _T_1027 & ~entry_found ? _GEN_12519 : _GEN_5861; // @[branch_predictor.scala 98:103]
  wire  _GEN_15592 = _T_1027 & ~entry_found ? _GEN_12520 : _GEN_5862; // @[branch_predictor.scala 98:103]
  wire  _GEN_15593 = _T_1027 & ~entry_found ? _GEN_12521 : _GEN_5863; // @[branch_predictor.scala 98:103]
  wire  _GEN_15594 = _T_1027 & ~entry_found ? _GEN_12522 : _GEN_5864; // @[branch_predictor.scala 98:103]
  wire  _GEN_15595 = _T_1027 & ~entry_found ? _GEN_12523 : _GEN_5865; // @[branch_predictor.scala 98:103]
  wire  _GEN_15596 = _T_1027 & ~entry_found ? _GEN_12524 : _GEN_5866; // @[branch_predictor.scala 98:103]
  wire  _GEN_15597 = _T_1027 & ~entry_found ? _GEN_12525 : _GEN_5867; // @[branch_predictor.scala 98:103]
  wire  _GEN_15598 = _T_1027 & ~entry_found ? _GEN_12526 : _GEN_5868; // @[branch_predictor.scala 98:103]
  wire  _GEN_15599 = _T_1027 & ~entry_found ? _GEN_12527 : _GEN_5869; // @[branch_predictor.scala 98:103]
  wire  _GEN_15600 = _T_1027 & ~entry_found ? _GEN_12528 : _GEN_5870; // @[branch_predictor.scala 98:103]
  wire  _GEN_15601 = _T_1027 & ~entry_found ? _GEN_12529 : _GEN_5871; // @[branch_predictor.scala 98:103]
  wire  _GEN_15602 = _T_1027 & ~entry_found ? _GEN_12530 : _GEN_5872; // @[branch_predictor.scala 98:103]
  wire  _GEN_15603 = _T_1027 & ~entry_found ? _GEN_12531 : _GEN_5873; // @[branch_predictor.scala 98:103]
  wire  _GEN_15604 = _T_1027 & ~entry_found ? _GEN_12532 : _GEN_5874; // @[branch_predictor.scala 98:103]
  wire  _GEN_15605 = _T_1027 & ~entry_found ? _GEN_12533 : _GEN_5875; // @[branch_predictor.scala 98:103]
  wire  _GEN_15606 = _T_1027 & ~entry_found ? _GEN_12534 : _GEN_5876; // @[branch_predictor.scala 98:103]
  wire  _GEN_15607 = _T_1027 & ~entry_found ? _GEN_12535 : _GEN_5877; // @[branch_predictor.scala 98:103]
  wire  _GEN_15608 = _T_1027 & ~entry_found ? _GEN_12536 : _GEN_5878; // @[branch_predictor.scala 98:103]
  wire  _GEN_15609 = _T_1027 & ~entry_found ? _GEN_12537 : _GEN_5879; // @[branch_predictor.scala 98:103]
  wire  _GEN_15610 = _T_1027 & ~entry_found ? _GEN_12538 : _GEN_5880; // @[branch_predictor.scala 98:103]
  wire  _GEN_15611 = _T_1027 & ~entry_found ? _GEN_12539 : _GEN_5881; // @[branch_predictor.scala 98:103]
  wire  _GEN_15612 = _T_1027 & ~entry_found ? _GEN_12540 : _GEN_5882; // @[branch_predictor.scala 98:103]
  wire  _GEN_15613 = _T_1027 & ~entry_found ? _GEN_12541 : _GEN_5883; // @[branch_predictor.scala 98:103]
  wire  _GEN_15614 = _T_1027 & ~entry_found ? _GEN_12542 : _GEN_5884; // @[branch_predictor.scala 98:103]
  wire  _GEN_15615 = _T_1027 & ~entry_found ? _GEN_12543 : _GEN_5885; // @[branch_predictor.scala 98:103]
  wire  _GEN_15616 = _T_1027 & ~entry_found ? _GEN_12544 : _GEN_5886; // @[branch_predictor.scala 98:103]
  wire  _GEN_15617 = _T_1027 & ~entry_found ? _GEN_12545 : _GEN_5887; // @[branch_predictor.scala 98:103]
  wire  _GEN_15618 = _T_1027 & ~entry_found ? _GEN_12546 : _GEN_5888; // @[branch_predictor.scala 98:103]
  wire  _GEN_15619 = _T_1027 & ~entry_found ? _GEN_12547 : _GEN_5889; // @[branch_predictor.scala 98:103]
  wire  _GEN_15620 = _T_1027 & ~entry_found ? _GEN_12548 : _GEN_5890; // @[branch_predictor.scala 98:103]
  wire  _GEN_15621 = _T_1027 & ~entry_found ? _GEN_12549 : _GEN_5891; // @[branch_predictor.scala 98:103]
  wire  _GEN_15622 = _T_1027 & ~entry_found ? _GEN_12550 : _GEN_5892; // @[branch_predictor.scala 98:103]
  wire  _GEN_15623 = _T_1027 & ~entry_found ? _GEN_12551 : _GEN_5893; // @[branch_predictor.scala 98:103]
  wire  _GEN_15624 = _T_1027 & ~entry_found ? _GEN_12552 : _GEN_5894; // @[branch_predictor.scala 98:103]
  wire  _GEN_15625 = _T_1027 & ~entry_found ? _GEN_12553 : _GEN_5895; // @[branch_predictor.scala 98:103]
  wire  _GEN_15626 = _T_1027 & ~entry_found ? _GEN_12554 : _GEN_5896; // @[branch_predictor.scala 98:103]
  wire  _GEN_15627 = _T_1027 & ~entry_found ? _GEN_12555 : _GEN_5897; // @[branch_predictor.scala 98:103]
  wire  _GEN_15628 = _T_1027 & ~entry_found ? _GEN_12556 : _GEN_5898; // @[branch_predictor.scala 98:103]
  wire  _GEN_15629 = _T_1027 & ~entry_found ? _GEN_12557 : _GEN_5899; // @[branch_predictor.scala 98:103]
  wire  _GEN_15630 = _T_1027 & ~entry_found ? _GEN_12558 : _GEN_5900; // @[branch_predictor.scala 98:103]
  wire  _GEN_15631 = _T_1027 & ~entry_found ? _GEN_12559 : _GEN_5901; // @[branch_predictor.scala 98:103]
  wire  _GEN_15632 = _T_1027 & ~entry_found ? _GEN_12560 : _GEN_5902; // @[branch_predictor.scala 98:103]
  wire  _GEN_15633 = _T_1027 & ~entry_found ? _GEN_12561 : _GEN_5903; // @[branch_predictor.scala 98:103]
  wire  _GEN_15634 = _T_1027 & ~entry_found ? _GEN_12562 : _GEN_5904; // @[branch_predictor.scala 98:103]
  wire  _GEN_15635 = _T_1027 & ~entry_found ? _GEN_12563 : _GEN_5905; // @[branch_predictor.scala 98:103]
  wire  _GEN_15636 = _T_1027 & ~entry_found ? _GEN_12564 : _GEN_5906; // @[branch_predictor.scala 98:103]
  wire  _GEN_15637 = _T_1027 & ~entry_found ? _GEN_12565 : _GEN_5907; // @[branch_predictor.scala 98:103]
  wire  _GEN_15638 = _T_1027 & ~entry_found ? _GEN_12566 : _GEN_5908; // @[branch_predictor.scala 98:103]
  wire  _GEN_15639 = _T_1027 & ~entry_found ? _GEN_12567 : _GEN_5909; // @[branch_predictor.scala 98:103]
  wire  _GEN_15640 = _T_1027 & ~entry_found ? _GEN_12568 : _GEN_5910; // @[branch_predictor.scala 98:103]
  wire  _GEN_15641 = _T_1027 & ~entry_found ? _GEN_12569 : _GEN_5911; // @[branch_predictor.scala 98:103]
  wire  _GEN_15642 = _T_1027 & ~entry_found ? _GEN_12570 : _GEN_5912; // @[branch_predictor.scala 98:103]
  wire  _GEN_15643 = _T_1027 & ~entry_found ? _GEN_12571 : _GEN_5913; // @[branch_predictor.scala 98:103]
  wire  _GEN_15644 = _T_1027 & ~entry_found ? _GEN_12572 : _GEN_5914; // @[branch_predictor.scala 98:103]
  wire  _GEN_15645 = _T_1027 & ~entry_found ? _GEN_12573 : _GEN_5915; // @[branch_predictor.scala 98:103]
  wire  _GEN_15646 = _T_1027 & ~entry_found ? _GEN_12574 : _GEN_5916; // @[branch_predictor.scala 98:103]
  wire  _GEN_15647 = _T_1027 & ~entry_found ? _GEN_12575 : _GEN_5917; // @[branch_predictor.scala 98:103]
  wire  _GEN_15648 = _T_1027 & ~entry_found ? _GEN_12576 : _GEN_5918; // @[branch_predictor.scala 98:103]
  wire  _GEN_15649 = _T_1027 & ~entry_found ? _GEN_12577 : _GEN_5919; // @[branch_predictor.scala 98:103]
  wire  _GEN_15650 = _T_1027 & ~entry_found ? _GEN_12578 : _GEN_5920; // @[branch_predictor.scala 98:103]
  wire  _GEN_15651 = _T_1027 & ~entry_found ? _GEN_12579 : _GEN_5921; // @[branch_predictor.scala 98:103]
  wire  _GEN_15652 = _T_1027 & ~entry_found ? _GEN_12580 : _GEN_5922; // @[branch_predictor.scala 98:103]
  wire  _GEN_15653 = _T_1027 & ~entry_found ? _GEN_12581 : _GEN_5923; // @[branch_predictor.scala 98:103]
  wire  _GEN_15654 = _T_1027 & ~entry_found ? _GEN_12582 : _GEN_5924; // @[branch_predictor.scala 98:103]
  wire  _GEN_15655 = _T_1027 & ~entry_found ? _GEN_12583 : _GEN_5925; // @[branch_predictor.scala 98:103]
  wire  _GEN_15656 = _T_1027 & ~entry_found ? _GEN_12584 : _GEN_5926; // @[branch_predictor.scala 98:103]
  wire  _GEN_15657 = _T_1027 & ~entry_found ? _GEN_12585 : _GEN_5927; // @[branch_predictor.scala 98:103]
  wire  _GEN_15658 = _T_1027 & ~entry_found ? _GEN_12586 : _GEN_5928; // @[branch_predictor.scala 98:103]
  wire  _GEN_15659 = _T_1027 & ~entry_found ? _GEN_12587 : _GEN_5929; // @[branch_predictor.scala 98:103]
  wire  _GEN_15660 = _T_1027 & ~entry_found ? _GEN_12588 : _GEN_5930; // @[branch_predictor.scala 98:103]
  wire  _GEN_15661 = _T_1027 & ~entry_found ? _GEN_12589 : _GEN_5931; // @[branch_predictor.scala 98:103]
  wire  _GEN_15662 = _T_1027 & ~entry_found ? _GEN_12590 : _GEN_5932; // @[branch_predictor.scala 98:103]
  wire  _GEN_15663 = _T_1027 & ~entry_found ? _GEN_12591 : _GEN_5933; // @[branch_predictor.scala 98:103]
  wire  _GEN_15664 = _T_1027 & ~entry_found ? _GEN_12592 : _GEN_5934; // @[branch_predictor.scala 98:103]
  wire  _GEN_15665 = _T_1027 & ~entry_found ? _GEN_12593 : _GEN_5935; // @[branch_predictor.scala 98:103]
  wire  _GEN_15666 = _T_1027 & ~entry_found ? _GEN_12594 : _GEN_5936; // @[branch_predictor.scala 98:103]
  wire  _GEN_15667 = _T_1027 & ~entry_found ? _GEN_12595 : _GEN_5937; // @[branch_predictor.scala 98:103]
  wire  _GEN_15668 = _T_1027 & ~entry_found ? _GEN_12596 : _GEN_5938; // @[branch_predictor.scala 98:103]
  wire  _GEN_15669 = _T_1027 & ~entry_found ? _GEN_12597 : _GEN_5939; // @[branch_predictor.scala 98:103]
  wire  _GEN_15670 = _T_1027 & ~entry_found ? _GEN_12598 : _GEN_5940; // @[branch_predictor.scala 98:103]
  wire  _GEN_15671 = _T_1027 & ~entry_found ? _GEN_12599 : _GEN_5941; // @[branch_predictor.scala 98:103]
  wire  _GEN_15672 = _T_1027 & ~entry_found ? _GEN_12600 : _GEN_5942; // @[branch_predictor.scala 98:103]
  wire  _GEN_15673 = _T_1027 & ~entry_found ? _GEN_12601 : _GEN_5943; // @[branch_predictor.scala 98:103]
  wire  _GEN_15674 = _T_1027 & ~entry_found ? _GEN_12602 : _GEN_5944; // @[branch_predictor.scala 98:103]
  wire  _GEN_15675 = _T_1027 & ~entry_found ? _GEN_12603 : _GEN_5945; // @[branch_predictor.scala 98:103]
  wire  _GEN_15676 = _T_1027 & ~entry_found ? _GEN_12604 : _GEN_5946; // @[branch_predictor.scala 98:103]
  wire  _GEN_15677 = _T_1027 & ~entry_found ? _GEN_12605 : _GEN_5947; // @[branch_predictor.scala 98:103]
  wire  _GEN_15678 = _T_1027 & ~entry_found ? _GEN_12606 : _GEN_5948; // @[branch_predictor.scala 98:103]
  wire  _GEN_15679 = _T_1027 & ~entry_found ? _GEN_12607 : _GEN_5949; // @[branch_predictor.scala 98:103]
  wire  _GEN_15680 = _T_1027 & ~entry_found ? _GEN_12608 : _GEN_5950; // @[branch_predictor.scala 98:103]
  wire  _GEN_15681 = _T_1027 & ~entry_found ? _GEN_12609 : _GEN_5951; // @[branch_predictor.scala 98:103]
  wire  _GEN_15682 = _T_1027 & ~entry_found ? _GEN_12610 : _GEN_5952; // @[branch_predictor.scala 98:103]
  wire  _GEN_15683 = _T_1027 & ~entry_found ? _GEN_12611 : _GEN_5953; // @[branch_predictor.scala 98:103]
  wire  _GEN_15684 = _T_1027 & ~entry_found ? _GEN_12612 : _GEN_5954; // @[branch_predictor.scala 98:103]
  wire  _GEN_15685 = _T_1027 & ~entry_found ? _GEN_12613 : _GEN_5955; // @[branch_predictor.scala 98:103]
  wire  _GEN_15686 = _T_1027 & ~entry_found ? _GEN_12614 : _GEN_5956; // @[branch_predictor.scala 98:103]
  wire  _GEN_15687 = _T_1027 & ~entry_found ? _GEN_12615 : _GEN_5957; // @[branch_predictor.scala 98:103]
  wire  _GEN_15688 = _T_1027 & ~entry_found ? _GEN_12616 : _GEN_5958; // @[branch_predictor.scala 98:103]
  wire  _GEN_15689 = _T_1027 & ~entry_found ? _GEN_12617 : _GEN_5959; // @[branch_predictor.scala 98:103]
  wire  _GEN_15690 = _T_1027 & ~entry_found ? _GEN_12618 : _GEN_5960; // @[branch_predictor.scala 98:103]
  wire  _GEN_15691 = _T_1027 & ~entry_found ? _GEN_12619 : _GEN_5961; // @[branch_predictor.scala 98:103]
  wire  _GEN_15692 = _T_1027 & ~entry_found ? _GEN_12620 : _GEN_5962; // @[branch_predictor.scala 98:103]
  wire  _GEN_15693 = _T_1027 & ~entry_found ? _GEN_12621 : _GEN_5963; // @[branch_predictor.scala 98:103]
  wire  _GEN_15694 = _T_1027 & ~entry_found ? _GEN_12622 : _GEN_5964; // @[branch_predictor.scala 98:103]
  wire  _GEN_15695 = _T_1027 & ~entry_found ? _GEN_12623 : _GEN_5965; // @[branch_predictor.scala 98:103]
  wire  _GEN_15696 = _T_1027 & ~entry_found ? _GEN_12624 : _GEN_5966; // @[branch_predictor.scala 98:103]
  wire  _GEN_15697 = _T_1027 & ~entry_found ? _GEN_12625 : _GEN_5967; // @[branch_predictor.scala 98:103]
  wire  _GEN_15698 = _T_1027 & ~entry_found ? _GEN_12626 : _GEN_5968; // @[branch_predictor.scala 98:103]
  wire  _GEN_15699 = _T_1027 & ~entry_found ? _GEN_12627 : _GEN_5969; // @[branch_predictor.scala 98:103]
  wire  _GEN_15700 = _T_1027 & ~entry_found ? _GEN_12628 : _GEN_5970; // @[branch_predictor.scala 98:103]
  wire  _GEN_15701 = _T_1027 & ~entry_found ? _GEN_12629 : _GEN_5971; // @[branch_predictor.scala 98:103]
  wire  _GEN_15702 = _T_1027 & ~entry_found ? _GEN_12630 : _GEN_5972; // @[branch_predictor.scala 98:103]
  wire  _GEN_15703 = _T_1027 & ~entry_found ? _GEN_12631 : _GEN_5973; // @[branch_predictor.scala 98:103]
  wire  _GEN_15704 = _T_1027 & ~entry_found ? _GEN_12632 : _GEN_5974; // @[branch_predictor.scala 98:103]
  wire  _GEN_15705 = _T_1027 & ~entry_found ? _GEN_12633 : _GEN_5975; // @[branch_predictor.scala 98:103]
  wire  _GEN_15706 = _T_1027 & ~entry_found ? _GEN_12634 : _GEN_5976; // @[branch_predictor.scala 98:103]
  wire  _GEN_15707 = _T_1027 & ~entry_found ? _GEN_12635 : _GEN_5977; // @[branch_predictor.scala 98:103]
  wire  _GEN_15708 = _T_1027 & ~entry_found ? _GEN_12636 : _GEN_5978; // @[branch_predictor.scala 98:103]
  wire  _GEN_15709 = _T_1027 & ~entry_found ? _GEN_12637 : _GEN_5979; // @[branch_predictor.scala 98:103]
  wire  _GEN_15710 = _T_1027 & ~entry_found ? _GEN_12638 : _GEN_5980; // @[branch_predictor.scala 98:103]
  wire  _GEN_15711 = _T_1027 & ~entry_found ? _GEN_12639 : _GEN_5981; // @[branch_predictor.scala 98:103]
  wire  _GEN_15712 = _T_1027 & ~entry_found ? _GEN_12640 : _GEN_5982; // @[branch_predictor.scala 98:103]
  wire  _GEN_15713 = _T_1027 & ~entry_found ? _GEN_12641 : _GEN_5983; // @[branch_predictor.scala 98:103]
  wire  _GEN_15714 = _T_1027 & ~entry_found ? _GEN_12642 : _GEN_5984; // @[branch_predictor.scala 98:103]
  wire  _GEN_15715 = _T_1027 & ~entry_found ? _GEN_12643 : _GEN_5985; // @[branch_predictor.scala 98:103]
  wire  _GEN_15716 = _T_1027 & ~entry_found ? _GEN_12644 : _GEN_5986; // @[branch_predictor.scala 98:103]
  wire  _GEN_15717 = _T_1027 & ~entry_found ? _GEN_12645 : _GEN_5987; // @[branch_predictor.scala 98:103]
  wire  _GEN_15718 = _T_1027 & ~entry_found ? _GEN_12646 : _GEN_5988; // @[branch_predictor.scala 98:103]
  wire  _GEN_15719 = _T_1027 & ~entry_found ? _GEN_12647 : _GEN_5989; // @[branch_predictor.scala 98:103]
  wire  _GEN_15720 = _T_1027 & ~entry_found ? _GEN_12648 : _GEN_5990; // @[branch_predictor.scala 98:103]
  wire  _GEN_15721 = _T_1027 & ~entry_found ? _GEN_12649 : _GEN_5991; // @[branch_predictor.scala 98:103]
  wire  _GEN_15722 = _T_1027 & ~entry_found ? _GEN_12650 : _GEN_5992; // @[branch_predictor.scala 98:103]
  wire  _GEN_15723 = _T_1027 & ~entry_found ? _GEN_12651 : _GEN_5993; // @[branch_predictor.scala 98:103]
  wire  _GEN_15724 = _T_1027 & ~entry_found ? _GEN_12652 : _GEN_5994; // @[branch_predictor.scala 98:103]
  wire  _GEN_15725 = _T_1027 & ~entry_found ? _GEN_12653 : _GEN_5995; // @[branch_predictor.scala 98:103]
  wire  _GEN_15726 = _T_1027 & ~entry_found ? _GEN_12654 : _GEN_5996; // @[branch_predictor.scala 98:103]
  wire  _GEN_15727 = _T_1027 & ~entry_found ? _GEN_12655 : _GEN_5997; // @[branch_predictor.scala 98:103]
  wire  _GEN_15728 = _T_1027 & ~entry_found ? _GEN_12656 : _GEN_5998; // @[branch_predictor.scala 98:103]
  wire  _GEN_15729 = _T_1027 & ~entry_found ? _GEN_12657 : _GEN_5999; // @[branch_predictor.scala 98:103]
  wire  _GEN_15730 = _T_1027 & ~entry_found ? _GEN_12658 : _GEN_6000; // @[branch_predictor.scala 98:103]
  wire  _GEN_15731 = _T_1027 & ~entry_found ? _GEN_12659 : _GEN_6001; // @[branch_predictor.scala 98:103]
  wire  _GEN_15732 = _T_1027 & ~entry_found ? _GEN_12660 : _GEN_6002; // @[branch_predictor.scala 98:103]
  wire  _GEN_15733 = _T_1027 & ~entry_found ? _GEN_12661 : _GEN_6003; // @[branch_predictor.scala 98:103]
  wire  _GEN_15734 = _T_1027 & ~entry_found ? _GEN_12662 : _GEN_6004; // @[branch_predictor.scala 98:103]
  wire  _GEN_15735 = _T_1027 & ~entry_found ? _GEN_12663 : _GEN_6005; // @[branch_predictor.scala 98:103]
  wire  _GEN_15736 = _T_1027 & ~entry_found ? _GEN_12664 : _GEN_6006; // @[branch_predictor.scala 98:103]
  wire  _GEN_15737 = _T_1027 & ~entry_found ? _GEN_12665 : _GEN_6007; // @[branch_predictor.scala 98:103]
  wire  _GEN_15738 = _T_1027 & ~entry_found ? _GEN_12666 : _GEN_6008; // @[branch_predictor.scala 98:103]
  wire  _GEN_15739 = _T_1027 & ~entry_found ? _GEN_12667 : _GEN_6009; // @[branch_predictor.scala 98:103]
  wire  _GEN_15740 = _T_1027 & ~entry_found ? _GEN_12668 : _GEN_6010; // @[branch_predictor.scala 98:103]
  wire  _GEN_15741 = _T_1027 & ~entry_found ? _GEN_12669 : _GEN_6011; // @[branch_predictor.scala 98:103]
  wire  _GEN_15742 = _T_1027 & ~entry_found ? _GEN_12670 : _GEN_6012; // @[branch_predictor.scala 98:103]
  wire  _GEN_15743 = _T_1027 & ~entry_found ? _GEN_12671 : _GEN_6013; // @[branch_predictor.scala 98:103]
  wire  _GEN_15744 = _T_1027 & ~entry_found ? _GEN_12672 : _GEN_6014; // @[branch_predictor.scala 98:103]
  wire  _GEN_15745 = _T_1027 & ~entry_found ? _GEN_12673 : _GEN_6015; // @[branch_predictor.scala 98:103]
  wire  _GEN_15746 = _T_1027 & ~entry_found ? _GEN_12674 : _GEN_6016; // @[branch_predictor.scala 98:103]
  wire  _GEN_15747 = _T_1027 & ~entry_found ? _GEN_12675 : _GEN_6017; // @[branch_predictor.scala 98:103]
  wire  _GEN_15748 = _T_1027 & ~entry_found ? _GEN_12676 : _GEN_6018; // @[branch_predictor.scala 98:103]
  wire  _GEN_15749 = _T_1027 & ~entry_found ? _GEN_12677 : _GEN_6019; // @[branch_predictor.scala 98:103]
  wire  _GEN_15750 = _T_1027 & ~entry_found ? _GEN_12678 : _GEN_6020; // @[branch_predictor.scala 98:103]
  wire  _GEN_15751 = _T_1027 & ~entry_found ? _GEN_12679 : _GEN_6021; // @[branch_predictor.scala 98:103]
  wire  _GEN_15752 = _T_1027 & ~entry_found ? _GEN_12680 : _GEN_6022; // @[branch_predictor.scala 98:103]
  wire  _GEN_15753 = _T_1027 & ~entry_found ? _GEN_12681 : _GEN_6023; // @[branch_predictor.scala 98:103]
  wire  _GEN_15754 = _T_1027 & ~entry_found ? _GEN_12682 : _GEN_6024; // @[branch_predictor.scala 98:103]
  wire  _GEN_15755 = _T_1027 & ~entry_found ? _GEN_12683 : _GEN_6025; // @[branch_predictor.scala 98:103]
  wire  _GEN_15756 = _T_1027 & ~entry_found ? _GEN_12684 : _GEN_6026; // @[branch_predictor.scala 98:103]
  wire  _GEN_15757 = _T_1027 & ~entry_found ? _GEN_12685 : _GEN_6027; // @[branch_predictor.scala 98:103]
  wire  _GEN_15758 = _T_1027 & ~entry_found ? _GEN_12686 : _GEN_6028; // @[branch_predictor.scala 98:103]
  wire  _GEN_15759 = _T_1027 & ~entry_found ? _GEN_12687 : _GEN_6029; // @[branch_predictor.scala 98:103]
  wire  _GEN_15760 = _T_1027 & ~entry_found ? _GEN_12688 : _GEN_6030; // @[branch_predictor.scala 98:103]
  wire  _GEN_15761 = _T_1027 & ~entry_found ? _GEN_12689 : _GEN_6031; // @[branch_predictor.scala 98:103]
  wire  _GEN_15762 = _T_1027 & ~entry_found ? _GEN_12690 : _GEN_6032; // @[branch_predictor.scala 98:103]
  wire  _GEN_15763 = _T_1027 & ~entry_found ? _GEN_12691 : _GEN_6033; // @[branch_predictor.scala 98:103]
  wire  _GEN_15764 = _T_1027 & ~entry_found ? _GEN_12692 : _GEN_6034; // @[branch_predictor.scala 98:103]
  wire  _GEN_15765 = _T_1027 & ~entry_found ? _GEN_12693 : _GEN_6035; // @[branch_predictor.scala 98:103]
  wire  _GEN_15766 = _T_1027 & ~entry_found ? _GEN_12694 : _GEN_6036; // @[branch_predictor.scala 98:103]
  wire  _GEN_15767 = _T_1027 & ~entry_found ? _GEN_12695 : _GEN_6037; // @[branch_predictor.scala 98:103]
  wire  _GEN_15768 = _T_1027 & ~entry_found ? _GEN_12696 : _GEN_6038; // @[branch_predictor.scala 98:103]
  wire  _GEN_15769 = _T_1027 & ~entry_found ? _GEN_12697 : _GEN_6039; // @[branch_predictor.scala 98:103]
  wire  _GEN_15770 = _T_1027 & ~entry_found ? _GEN_12698 : _GEN_6040; // @[branch_predictor.scala 98:103]
  wire  _GEN_15771 = _T_1027 & ~entry_found ? _GEN_12699 : _GEN_6041; // @[branch_predictor.scala 98:103]
  wire  _GEN_15772 = _T_1027 & ~entry_found ? _GEN_12700 : _GEN_6042; // @[branch_predictor.scala 98:103]
  wire  _GEN_15773 = _T_1027 & ~entry_found ? _GEN_12701 : _GEN_6043; // @[branch_predictor.scala 98:103]
  wire  _GEN_15774 = _T_1027 & ~entry_found ? _GEN_12702 : _GEN_6044; // @[branch_predictor.scala 98:103]
  wire  _GEN_15775 = _T_1027 & ~entry_found ? _GEN_12703 : _GEN_6045; // @[branch_predictor.scala 98:103]
  wire  _GEN_15776 = _T_1027 & ~entry_found ? _GEN_12704 : _GEN_6046; // @[branch_predictor.scala 98:103]
  wire  _GEN_15777 = _T_1027 & ~entry_found ? _GEN_12705 : _GEN_6047; // @[branch_predictor.scala 98:103]
  wire  _GEN_15778 = _T_1027 & ~entry_found ? _GEN_12706 : _GEN_6048; // @[branch_predictor.scala 98:103]
  wire  _GEN_15779 = _T_1027 & ~entry_found ? _GEN_12707 : _GEN_6049; // @[branch_predictor.scala 98:103]
  wire  _GEN_15780 = _T_1027 & ~entry_found ? _GEN_12708 : _GEN_6050; // @[branch_predictor.scala 98:103]
  wire  _GEN_15781 = _T_1027 & ~entry_found ? _GEN_12709 : _GEN_6051; // @[branch_predictor.scala 98:103]
  wire  _GEN_15782 = _T_1027 & ~entry_found ? _GEN_12710 : _GEN_6052; // @[branch_predictor.scala 98:103]
  wire  _GEN_15783 = _T_1027 & ~entry_found ? _GEN_12711 : _GEN_6053; // @[branch_predictor.scala 98:103]
  wire  _GEN_15784 = _T_1027 & ~entry_found ? _GEN_12712 : _GEN_6054; // @[branch_predictor.scala 98:103]
  wire  _GEN_15785 = _T_1027 & ~entry_found ? _GEN_12713 : _GEN_6055; // @[branch_predictor.scala 98:103]
  wire  _GEN_15786 = _T_1027 & ~entry_found ? _GEN_12714 : _GEN_6056; // @[branch_predictor.scala 98:103]
  wire  _GEN_15787 = _T_1027 & ~entry_found ? _GEN_12715 : _GEN_6057; // @[branch_predictor.scala 98:103]
  wire  _GEN_15788 = _T_1027 & ~entry_found ? _GEN_12716 : _GEN_6058; // @[branch_predictor.scala 98:103]
  wire  _GEN_15789 = _T_1027 & ~entry_found ? _GEN_12717 : _GEN_6059; // @[branch_predictor.scala 98:103]
  wire  _GEN_15790 = _T_1027 & ~entry_found ? _GEN_12718 : _GEN_6060; // @[branch_predictor.scala 98:103]
  wire  _GEN_15791 = _T_1027 & ~entry_found ? _GEN_12719 : _GEN_6061; // @[branch_predictor.scala 98:103]
  wire  _GEN_15792 = _T_1027 & ~entry_found ? _GEN_12720 : _GEN_6062; // @[branch_predictor.scala 98:103]
  wire  _GEN_15793 = _T_1027 & ~entry_found ? _GEN_12721 : _GEN_6063; // @[branch_predictor.scala 98:103]
  wire  _GEN_15794 = _T_1027 & ~entry_found ? _GEN_12722 : _GEN_6064; // @[branch_predictor.scala 98:103]
  wire  _GEN_15795 = _T_1027 & ~entry_found ? _GEN_12723 : _GEN_6065; // @[branch_predictor.scala 98:103]
  wire  _GEN_15796 = _T_1027 & ~entry_found ? _GEN_12724 : _GEN_6066; // @[branch_predictor.scala 98:103]
  wire  _GEN_15797 = _T_1027 & ~entry_found ? _GEN_12725 : _GEN_6067; // @[branch_predictor.scala 98:103]
  wire  _GEN_15798 = _T_1027 & ~entry_found ? _GEN_12726 : _GEN_6068; // @[branch_predictor.scala 98:103]
  wire  _GEN_15799 = _T_1027 & ~entry_found ? _GEN_12727 : _GEN_6069; // @[branch_predictor.scala 98:103]
  wire  _GEN_15800 = _T_1027 & ~entry_found ? _GEN_12728 : _GEN_6070; // @[branch_predictor.scala 98:103]
  wire  _GEN_15801 = _T_1027 & ~entry_found ? _GEN_12729 : _GEN_6071; // @[branch_predictor.scala 98:103]
  wire  _GEN_15802 = _T_1027 & ~entry_found ? _GEN_12730 : _GEN_6072; // @[branch_predictor.scala 98:103]
  wire  _GEN_15803 = _T_1027 & ~entry_found ? _GEN_12731 : _GEN_6073; // @[branch_predictor.scala 98:103]
  wire  _GEN_15804 = _T_1027 & ~entry_found ? _GEN_12732 : _GEN_6074; // @[branch_predictor.scala 98:103]
  wire  _GEN_15805 = _T_1027 & ~entry_found ? _GEN_12733 : _GEN_6075; // @[branch_predictor.scala 98:103]
  wire  _GEN_15806 = _T_1027 & ~entry_found ? _GEN_12734 : _GEN_6076; // @[branch_predictor.scala 98:103]
  wire  _GEN_15807 = _T_1027 & ~entry_found ? _GEN_12735 : _GEN_6077; // @[branch_predictor.scala 98:103]
  wire  _GEN_15808 = _T_1027 & ~entry_found ? _GEN_12736 : _GEN_6078; // @[branch_predictor.scala 98:103]
  wire  _GEN_15809 = _T_1027 & ~entry_found ? _GEN_12737 : _GEN_6079; // @[branch_predictor.scala 98:103]
  wire  _GEN_15810 = _T_1027 & ~entry_found ? _GEN_12738 : _GEN_6080; // @[branch_predictor.scala 98:103]
  wire  _GEN_15811 = _T_1027 & ~entry_found ? _GEN_12739 : _GEN_6081; // @[branch_predictor.scala 98:103]
  wire  _GEN_15812 = _T_1027 & ~entry_found ? _GEN_12740 : _GEN_6082; // @[branch_predictor.scala 98:103]
  wire  _GEN_15813 = _T_1027 & ~entry_found ? _GEN_12741 : _GEN_6083; // @[branch_predictor.scala 98:103]
  wire  _GEN_15814 = _T_1027 & ~entry_found ? _GEN_12742 : _GEN_6084; // @[branch_predictor.scala 98:103]
  wire  _GEN_15815 = _T_1027 & ~entry_found ? _GEN_12743 : _GEN_6085; // @[branch_predictor.scala 98:103]
  wire  _GEN_15816 = _T_1027 & ~entry_found ? _GEN_12744 : _GEN_6086; // @[branch_predictor.scala 98:103]
  wire  _GEN_15817 = _T_1027 & ~entry_found ? _GEN_12745 : _GEN_6087; // @[branch_predictor.scala 98:103]
  wire  _GEN_15818 = _T_1027 & ~entry_found ? _GEN_12746 : _GEN_6088; // @[branch_predictor.scala 98:103]
  wire  _GEN_15819 = _T_1027 & ~entry_found ? _GEN_12747 : _GEN_6089; // @[branch_predictor.scala 98:103]
  wire  _GEN_15820 = _T_1027 & ~entry_found ? _GEN_12748 : _GEN_6090; // @[branch_predictor.scala 98:103]
  wire  _GEN_15821 = _T_1027 & ~entry_found ? _GEN_12749 : _GEN_6091; // @[branch_predictor.scala 98:103]
  wire  _GEN_15822 = _T_1027 & ~entry_found ? _GEN_12750 : _GEN_6092; // @[branch_predictor.scala 98:103]
  wire  _GEN_15823 = _T_1027 & ~entry_found ? _GEN_12751 : _GEN_6093; // @[branch_predictor.scala 98:103]
  wire  _GEN_15824 = _T_1027 & ~entry_found ? _GEN_12752 : _GEN_6094; // @[branch_predictor.scala 98:103]
  wire  _GEN_15825 = _T_1027 & ~entry_found ? _GEN_12753 : _GEN_6095; // @[branch_predictor.scala 98:103]
  wire  _GEN_15826 = _T_1027 & ~entry_found ? _GEN_12754 : _GEN_6096; // @[branch_predictor.scala 98:103]
  wire  _GEN_15827 = _T_1027 & ~entry_found ? _GEN_12755 : _GEN_6097; // @[branch_predictor.scala 98:103]
  wire  _GEN_15828 = _T_1027 & ~entry_found ? _GEN_12756 : _GEN_6098; // @[branch_predictor.scala 98:103]
  wire  _GEN_15829 = _T_1027 & ~entry_found ? _GEN_12757 : _GEN_6099; // @[branch_predictor.scala 98:103]
  wire  _GEN_15830 = _T_1027 & ~entry_found ? _GEN_12758 : _GEN_6100; // @[branch_predictor.scala 98:103]
  wire  _GEN_15831 = _T_1027 & ~entry_found ? _GEN_12759 : _GEN_6101; // @[branch_predictor.scala 98:103]
  wire  _GEN_15832 = _T_1027 & ~entry_found ? _GEN_12760 : _GEN_6102; // @[branch_predictor.scala 98:103]
  wire  _GEN_15833 = _T_1027 & ~entry_found ? _GEN_12761 : _GEN_6103; // @[branch_predictor.scala 98:103]
  wire  _GEN_15834 = _T_1027 & ~entry_found ? _GEN_12762 : _GEN_6104; // @[branch_predictor.scala 98:103]
  wire  _GEN_15835 = _T_1027 & ~entry_found ? _GEN_12763 : _GEN_6105; // @[branch_predictor.scala 98:103]
  wire  _GEN_15836 = _T_1027 & ~entry_found ? _GEN_12764 : _GEN_6106; // @[branch_predictor.scala 98:103]
  wire  _GEN_15837 = _T_1027 & ~entry_found ? _GEN_12765 : _GEN_6107; // @[branch_predictor.scala 98:103]
  wire  _GEN_15838 = _T_1027 & ~entry_found ? _GEN_12766 : _GEN_6108; // @[branch_predictor.scala 98:103]
  wire  _GEN_15839 = _T_1027 & ~entry_found ? _GEN_12767 : _GEN_6109; // @[branch_predictor.scala 98:103]
  wire  _GEN_15840 = _T_1027 & ~entry_found ? _GEN_12768 : _GEN_6110; // @[branch_predictor.scala 98:103]
  wire  _GEN_15841 = _T_1027 & ~entry_found ? _GEN_12769 : _GEN_6111; // @[branch_predictor.scala 98:103]
  wire  _GEN_15842 = _T_1027 & ~entry_found ? _GEN_12770 : _GEN_6112; // @[branch_predictor.scala 98:103]
  wire  _GEN_15843 = _T_1027 & ~entry_found ? _GEN_12771 : _GEN_6113; // @[branch_predictor.scala 98:103]
  wire  _GEN_15844 = _T_1027 & ~entry_found ? _GEN_12772 : _GEN_6114; // @[branch_predictor.scala 98:103]
  wire  _GEN_15845 = _T_1027 & ~entry_found ? _GEN_12773 : _GEN_6115; // @[branch_predictor.scala 98:103]
  wire  _GEN_15846 = _T_1027 & ~entry_found ? _GEN_12774 : _GEN_6116; // @[branch_predictor.scala 98:103]
  wire  _GEN_15847 = _T_1027 & ~entry_found ? _GEN_12775 : _GEN_6117; // @[branch_predictor.scala 98:103]
  wire  _GEN_15848 = _T_1027 & ~entry_found ? _GEN_12776 : _GEN_6118; // @[branch_predictor.scala 98:103]
  wire  _GEN_15849 = _T_1027 & ~entry_found ? _GEN_12777 : _GEN_6119; // @[branch_predictor.scala 98:103]
  wire  _GEN_15850 = _T_1027 & ~entry_found ? _GEN_12778 : _GEN_6120; // @[branch_predictor.scala 98:103]
  wire  _GEN_15851 = _T_1027 & ~entry_found ? _GEN_12779 : _GEN_6121; // @[branch_predictor.scala 98:103]
  wire  _GEN_15852 = _T_1027 & ~entry_found ? _GEN_12780 : _GEN_6122; // @[branch_predictor.scala 98:103]
  wire  _GEN_15853 = _T_1027 & ~entry_found ? _GEN_12781 : _GEN_6123; // @[branch_predictor.scala 98:103]
  wire  _GEN_15854 = _T_1027 & ~entry_found ? _GEN_12782 : _GEN_6124; // @[branch_predictor.scala 98:103]
  wire  _GEN_15855 = _T_1027 & ~entry_found ? _GEN_12783 : _GEN_6125; // @[branch_predictor.scala 98:103]
  wire  _GEN_15856 = _T_1027 & ~entry_found ? _GEN_12784 : _GEN_6126; // @[branch_predictor.scala 98:103]
  wire  _GEN_15857 = _T_1027 & ~entry_found ? _GEN_12785 : _GEN_6127; // @[branch_predictor.scala 98:103]
  wire  _GEN_15858 = _T_1027 & ~entry_found ? _GEN_12786 : _GEN_6128; // @[branch_predictor.scala 98:103]
  wire  _GEN_15859 = _T_1027 & ~entry_found ? _GEN_12787 : _GEN_6129; // @[branch_predictor.scala 98:103]
  wire  _GEN_15860 = _T_1027 & ~entry_found ? _GEN_12788 : _GEN_6130; // @[branch_predictor.scala 98:103]
  wire  _GEN_15861 = _T_1027 & ~entry_found ? _GEN_12789 : _GEN_6131; // @[branch_predictor.scala 98:103]
  wire  _GEN_15862 = _T_1027 & ~entry_found ? _GEN_12790 : _GEN_6132; // @[branch_predictor.scala 98:103]
  wire  _GEN_15863 = _T_1027 & ~entry_found ? _GEN_12791 : _GEN_6133; // @[branch_predictor.scala 98:103]
  wire  _GEN_15864 = _T_1027 & ~entry_found ? _GEN_12792 : _GEN_6134; // @[branch_predictor.scala 98:103]
  wire  _GEN_15865 = _T_1027 & ~entry_found ? _GEN_12793 : _GEN_6135; // @[branch_predictor.scala 98:103]
  wire  _GEN_15866 = _T_1027 & ~entry_found ? _GEN_12794 : _GEN_6136; // @[branch_predictor.scala 98:103]
  wire  _GEN_15867 = _T_1027 & ~entry_found ? _GEN_12795 : _GEN_6137; // @[branch_predictor.scala 98:103]
  wire  _GEN_15868 = _T_1027 & ~entry_found ? _GEN_12796 : _GEN_6138; // @[branch_predictor.scala 98:103]
  wire  _GEN_15869 = _T_1027 & ~entry_found ? _GEN_12797 : _GEN_6139; // @[branch_predictor.scala 98:103]
  wire  _GEN_15870 = _T_1027 & ~entry_found ? _GEN_12798 : _GEN_6140; // @[branch_predictor.scala 98:103]
  wire  _GEN_15871 = _T_1027 & ~entry_found ? _GEN_12799 : _GEN_6141; // @[branch_predictor.scala 98:103]
  wire  _GEN_15872 = _T_1027 & ~entry_found ? _GEN_12800 : _GEN_6142; // @[branch_predictor.scala 98:103]
  wire  _GEN_15873 = _T_1027 & ~entry_found ? _GEN_12801 : _GEN_6143; // @[branch_predictor.scala 98:103]
  assign io_o_branch_predict_pack_valid = btb_511_tag == io_i_addr[12:3] ? btb_511_valid : _GEN_2550; // @[branch_predictor.scala 40:45 41:44]
  assign io_o_branch_predict_pack_target = btb_511_tag == io_i_addr[12:3] ? btb_511_target_address : _GEN_2551; // @[branch_predictor.scala 40:45 42:45]
  assign io_o_branch_predict_pack_taken = btb_511_tag == io_i_addr[12:3] ? ~btb_511_bht[1] : _GEN_2554; // @[branch_predictor.scala 40:45 45:44]
  always @(posedge clock) begin
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_0_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_0_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_0_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_0_valid <= _GEN_15362;
      end
    end else begin
      btb_0_valid <= _GEN_15362;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_0_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_0_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_0_tag <= _GEN_6144;
      end
    end else begin
      btb_0_tag <= _GEN_6144;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_0_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_0_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_0_target_address <= _GEN_10754;
      end
    end else begin
      btb_0_target_address <= _GEN_10754;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_0_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_0_bht <= 2'h1;
        end else begin
          btb_0_bht <= 2'h0;
        end
      end else begin
        btb_0_bht <= _GEN_10756;
      end
    end else begin
      btb_0_bht <= _GEN_10756;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_1_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_1_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_1_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_1_valid <= _GEN_15363;
      end
    end else begin
      btb_1_valid <= _GEN_15363;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_1_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_1_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_1_tag <= _GEN_6145;
      end
    end else begin
      btb_1_tag <= _GEN_6145;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_1_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_1_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_1_target_address <= _GEN_10757;
      end
    end else begin
      btb_1_target_address <= _GEN_10757;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_1_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_1_bht <= 2'h1;
        end else begin
          btb_1_bht <= 2'h0;
        end
      end else begin
        btb_1_bht <= _GEN_10759;
      end
    end else begin
      btb_1_bht <= _GEN_10759;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_2_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_2_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_2_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_2_valid <= _GEN_15364;
      end
    end else begin
      btb_2_valid <= _GEN_15364;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_2_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_2_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_2_tag <= _GEN_6146;
      end
    end else begin
      btb_2_tag <= _GEN_6146;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_2_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_2_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_2_target_address <= _GEN_10760;
      end
    end else begin
      btb_2_target_address <= _GEN_10760;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_2_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_2_bht <= 2'h1;
        end else begin
          btb_2_bht <= 2'h0;
        end
      end else begin
        btb_2_bht <= _GEN_10762;
      end
    end else begin
      btb_2_bht <= _GEN_10762;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_3_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_3_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_3_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_3_valid <= _GEN_15365;
      end
    end else begin
      btb_3_valid <= _GEN_15365;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_3_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_3_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_3_tag <= _GEN_6147;
      end
    end else begin
      btb_3_tag <= _GEN_6147;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_3_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_3_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_3_target_address <= _GEN_10763;
      end
    end else begin
      btb_3_target_address <= _GEN_10763;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_3_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_3_bht <= 2'h1;
        end else begin
          btb_3_bht <= 2'h0;
        end
      end else begin
        btb_3_bht <= _GEN_10765;
      end
    end else begin
      btb_3_bht <= _GEN_10765;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_4_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_4_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_4_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_4_valid <= _GEN_15366;
      end
    end else begin
      btb_4_valid <= _GEN_15366;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_4_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_4_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_4_tag <= _GEN_6148;
      end
    end else begin
      btb_4_tag <= _GEN_6148;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_4_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_4_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_4_target_address <= _GEN_10766;
      end
    end else begin
      btb_4_target_address <= _GEN_10766;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_4_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_4_bht <= 2'h1;
        end else begin
          btb_4_bht <= 2'h0;
        end
      end else begin
        btb_4_bht <= _GEN_10768;
      end
    end else begin
      btb_4_bht <= _GEN_10768;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_5_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_5_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_5_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_5_valid <= _GEN_15367;
      end
    end else begin
      btb_5_valid <= _GEN_15367;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_5_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_5_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_5_tag <= _GEN_6149;
      end
    end else begin
      btb_5_tag <= _GEN_6149;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_5_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_5_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_5_target_address <= _GEN_10769;
      end
    end else begin
      btb_5_target_address <= _GEN_10769;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_5_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_5_bht <= 2'h1;
        end else begin
          btb_5_bht <= 2'h0;
        end
      end else begin
        btb_5_bht <= _GEN_10771;
      end
    end else begin
      btb_5_bht <= _GEN_10771;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_6_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_6_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_6_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_6_valid <= _GEN_15368;
      end
    end else begin
      btb_6_valid <= _GEN_15368;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_6_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_6_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_6_tag <= _GEN_6150;
      end
    end else begin
      btb_6_tag <= _GEN_6150;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_6_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_6_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_6_target_address <= _GEN_10772;
      end
    end else begin
      btb_6_target_address <= _GEN_10772;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_6_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_6_bht <= 2'h1;
        end else begin
          btb_6_bht <= 2'h0;
        end
      end else begin
        btb_6_bht <= _GEN_10774;
      end
    end else begin
      btb_6_bht <= _GEN_10774;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_7_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_7_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_7_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_7_valid <= _GEN_15369;
      end
    end else begin
      btb_7_valid <= _GEN_15369;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_7_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_7_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_7_tag <= _GEN_6151;
      end
    end else begin
      btb_7_tag <= _GEN_6151;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_7_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_7_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_7_target_address <= _GEN_10775;
      end
    end else begin
      btb_7_target_address <= _GEN_10775;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_7_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_7_bht <= 2'h1;
        end else begin
          btb_7_bht <= 2'h0;
        end
      end else begin
        btb_7_bht <= _GEN_10777;
      end
    end else begin
      btb_7_bht <= _GEN_10777;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_8_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_8_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_8_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_8_valid <= _GEN_15370;
      end
    end else begin
      btb_8_valid <= _GEN_15370;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_8_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_8_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_8_tag <= _GEN_6152;
      end
    end else begin
      btb_8_tag <= _GEN_6152;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_8_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_8_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_8_target_address <= _GEN_10778;
      end
    end else begin
      btb_8_target_address <= _GEN_10778;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_8_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_8_bht <= 2'h1;
        end else begin
          btb_8_bht <= 2'h0;
        end
      end else begin
        btb_8_bht <= _GEN_10780;
      end
    end else begin
      btb_8_bht <= _GEN_10780;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_9_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_9_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_9_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_9_valid <= _GEN_15371;
      end
    end else begin
      btb_9_valid <= _GEN_15371;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_9_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_9_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_9_tag <= _GEN_6153;
      end
    end else begin
      btb_9_tag <= _GEN_6153;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_9_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_9_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_9_target_address <= _GEN_10781;
      end
    end else begin
      btb_9_target_address <= _GEN_10781;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_9_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_9_bht <= 2'h1;
        end else begin
          btb_9_bht <= 2'h0;
        end
      end else begin
        btb_9_bht <= _GEN_10783;
      end
    end else begin
      btb_9_bht <= _GEN_10783;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_10_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_10_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_10_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_10_valid <= _GEN_15372;
      end
    end else begin
      btb_10_valid <= _GEN_15372;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_10_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_10_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_10_tag <= _GEN_6154;
      end
    end else begin
      btb_10_tag <= _GEN_6154;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_10_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_10_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_10_target_address <= _GEN_10784;
      end
    end else begin
      btb_10_target_address <= _GEN_10784;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_10_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_10_bht <= 2'h1;
        end else begin
          btb_10_bht <= 2'h0;
        end
      end else begin
        btb_10_bht <= _GEN_10786;
      end
    end else begin
      btb_10_bht <= _GEN_10786;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_11_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_11_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_11_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_11_valid <= _GEN_15373;
      end
    end else begin
      btb_11_valid <= _GEN_15373;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_11_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_11_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_11_tag <= _GEN_6155;
      end
    end else begin
      btb_11_tag <= _GEN_6155;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_11_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_11_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_11_target_address <= _GEN_10787;
      end
    end else begin
      btb_11_target_address <= _GEN_10787;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_11_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_11_bht <= 2'h1;
        end else begin
          btb_11_bht <= 2'h0;
        end
      end else begin
        btb_11_bht <= _GEN_10789;
      end
    end else begin
      btb_11_bht <= _GEN_10789;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_12_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_12_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_12_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_12_valid <= _GEN_15374;
      end
    end else begin
      btb_12_valid <= _GEN_15374;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_12_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_12_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_12_tag <= _GEN_6156;
      end
    end else begin
      btb_12_tag <= _GEN_6156;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_12_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_12_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_12_target_address <= _GEN_10790;
      end
    end else begin
      btb_12_target_address <= _GEN_10790;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_12_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_12_bht <= 2'h1;
        end else begin
          btb_12_bht <= 2'h0;
        end
      end else begin
        btb_12_bht <= _GEN_10792;
      end
    end else begin
      btb_12_bht <= _GEN_10792;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_13_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_13_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_13_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_13_valid <= _GEN_15375;
      end
    end else begin
      btb_13_valid <= _GEN_15375;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_13_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_13_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_13_tag <= _GEN_6157;
      end
    end else begin
      btb_13_tag <= _GEN_6157;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_13_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_13_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_13_target_address <= _GEN_10793;
      end
    end else begin
      btb_13_target_address <= _GEN_10793;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_13_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_13_bht <= 2'h1;
        end else begin
          btb_13_bht <= 2'h0;
        end
      end else begin
        btb_13_bht <= _GEN_10795;
      end
    end else begin
      btb_13_bht <= _GEN_10795;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_14_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_14_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_14_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_14_valid <= _GEN_15376;
      end
    end else begin
      btb_14_valid <= _GEN_15376;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_14_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_14_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_14_tag <= _GEN_6158;
      end
    end else begin
      btb_14_tag <= _GEN_6158;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_14_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_14_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_14_target_address <= _GEN_10796;
      end
    end else begin
      btb_14_target_address <= _GEN_10796;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_14_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_14_bht <= 2'h1;
        end else begin
          btb_14_bht <= 2'h0;
        end
      end else begin
        btb_14_bht <= _GEN_10798;
      end
    end else begin
      btb_14_bht <= _GEN_10798;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_15_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_15_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_15_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_15_valid <= _GEN_15377;
      end
    end else begin
      btb_15_valid <= _GEN_15377;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_15_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_15_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_15_tag <= _GEN_6159;
      end
    end else begin
      btb_15_tag <= _GEN_6159;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_15_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_15_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_15_target_address <= _GEN_10799;
      end
    end else begin
      btb_15_target_address <= _GEN_10799;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_15_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_15_bht <= 2'h1;
        end else begin
          btb_15_bht <= 2'h0;
        end
      end else begin
        btb_15_bht <= _GEN_10801;
      end
    end else begin
      btb_15_bht <= _GEN_10801;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_16_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_16_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_16_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_16_valid <= _GEN_15378;
      end
    end else begin
      btb_16_valid <= _GEN_15378;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_16_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_16_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_16_tag <= _GEN_6160;
      end
    end else begin
      btb_16_tag <= _GEN_6160;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_16_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_16_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_16_target_address <= _GEN_10802;
      end
    end else begin
      btb_16_target_address <= _GEN_10802;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_16_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_16_bht <= 2'h1;
        end else begin
          btb_16_bht <= 2'h0;
        end
      end else begin
        btb_16_bht <= _GEN_10804;
      end
    end else begin
      btb_16_bht <= _GEN_10804;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_17_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_17_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_17_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_17_valid <= _GEN_15379;
      end
    end else begin
      btb_17_valid <= _GEN_15379;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_17_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_17_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_17_tag <= _GEN_6161;
      end
    end else begin
      btb_17_tag <= _GEN_6161;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_17_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_17_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_17_target_address <= _GEN_10805;
      end
    end else begin
      btb_17_target_address <= _GEN_10805;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_17_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_17_bht <= 2'h1;
        end else begin
          btb_17_bht <= 2'h0;
        end
      end else begin
        btb_17_bht <= _GEN_10807;
      end
    end else begin
      btb_17_bht <= _GEN_10807;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_18_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_18_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_18_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_18_valid <= _GEN_15380;
      end
    end else begin
      btb_18_valid <= _GEN_15380;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_18_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_18_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_18_tag <= _GEN_6162;
      end
    end else begin
      btb_18_tag <= _GEN_6162;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_18_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_18_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_18_target_address <= _GEN_10808;
      end
    end else begin
      btb_18_target_address <= _GEN_10808;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_18_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_18_bht <= 2'h1;
        end else begin
          btb_18_bht <= 2'h0;
        end
      end else begin
        btb_18_bht <= _GEN_10810;
      end
    end else begin
      btb_18_bht <= _GEN_10810;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_19_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_19_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_19_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_19_valid <= _GEN_15381;
      end
    end else begin
      btb_19_valid <= _GEN_15381;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_19_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_19_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_19_tag <= _GEN_6163;
      end
    end else begin
      btb_19_tag <= _GEN_6163;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_19_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_19_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_19_target_address <= _GEN_10811;
      end
    end else begin
      btb_19_target_address <= _GEN_10811;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_19_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_19_bht <= 2'h1;
        end else begin
          btb_19_bht <= 2'h0;
        end
      end else begin
        btb_19_bht <= _GEN_10813;
      end
    end else begin
      btb_19_bht <= _GEN_10813;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_20_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_20_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_20_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_20_valid <= _GEN_15382;
      end
    end else begin
      btb_20_valid <= _GEN_15382;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_20_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_20_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_20_tag <= _GEN_6164;
      end
    end else begin
      btb_20_tag <= _GEN_6164;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_20_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_20_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_20_target_address <= _GEN_10814;
      end
    end else begin
      btb_20_target_address <= _GEN_10814;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_20_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_20_bht <= 2'h1;
        end else begin
          btb_20_bht <= 2'h0;
        end
      end else begin
        btb_20_bht <= _GEN_10816;
      end
    end else begin
      btb_20_bht <= _GEN_10816;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_21_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_21_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_21_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_21_valid <= _GEN_15383;
      end
    end else begin
      btb_21_valid <= _GEN_15383;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_21_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_21_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_21_tag <= _GEN_6165;
      end
    end else begin
      btb_21_tag <= _GEN_6165;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_21_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_21_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_21_target_address <= _GEN_10817;
      end
    end else begin
      btb_21_target_address <= _GEN_10817;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_21_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_21_bht <= 2'h1;
        end else begin
          btb_21_bht <= 2'h0;
        end
      end else begin
        btb_21_bht <= _GEN_10819;
      end
    end else begin
      btb_21_bht <= _GEN_10819;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_22_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_22_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_22_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_22_valid <= _GEN_15384;
      end
    end else begin
      btb_22_valid <= _GEN_15384;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_22_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_22_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_22_tag <= _GEN_6166;
      end
    end else begin
      btb_22_tag <= _GEN_6166;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_22_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_22_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_22_target_address <= _GEN_10820;
      end
    end else begin
      btb_22_target_address <= _GEN_10820;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_22_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_22_bht <= 2'h1;
        end else begin
          btb_22_bht <= 2'h0;
        end
      end else begin
        btb_22_bht <= _GEN_10822;
      end
    end else begin
      btb_22_bht <= _GEN_10822;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_23_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_23_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_23_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_23_valid <= _GEN_15385;
      end
    end else begin
      btb_23_valid <= _GEN_15385;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_23_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_23_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_23_tag <= _GEN_6167;
      end
    end else begin
      btb_23_tag <= _GEN_6167;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_23_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_23_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_23_target_address <= _GEN_10823;
      end
    end else begin
      btb_23_target_address <= _GEN_10823;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_23_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_23_bht <= 2'h1;
        end else begin
          btb_23_bht <= 2'h0;
        end
      end else begin
        btb_23_bht <= _GEN_10825;
      end
    end else begin
      btb_23_bht <= _GEN_10825;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_24_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_24_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_24_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_24_valid <= _GEN_15386;
      end
    end else begin
      btb_24_valid <= _GEN_15386;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_24_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_24_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_24_tag <= _GEN_6168;
      end
    end else begin
      btb_24_tag <= _GEN_6168;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_24_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_24_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_24_target_address <= _GEN_10826;
      end
    end else begin
      btb_24_target_address <= _GEN_10826;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_24_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_24_bht <= 2'h1;
        end else begin
          btb_24_bht <= 2'h0;
        end
      end else begin
        btb_24_bht <= _GEN_10828;
      end
    end else begin
      btb_24_bht <= _GEN_10828;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_25_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_25_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_25_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_25_valid <= _GEN_15387;
      end
    end else begin
      btb_25_valid <= _GEN_15387;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_25_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_25_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_25_tag <= _GEN_6169;
      end
    end else begin
      btb_25_tag <= _GEN_6169;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_25_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_25_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_25_target_address <= _GEN_10829;
      end
    end else begin
      btb_25_target_address <= _GEN_10829;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_25_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_25_bht <= 2'h1;
        end else begin
          btb_25_bht <= 2'h0;
        end
      end else begin
        btb_25_bht <= _GEN_10831;
      end
    end else begin
      btb_25_bht <= _GEN_10831;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_26_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_26_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_26_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_26_valid <= _GEN_15388;
      end
    end else begin
      btb_26_valid <= _GEN_15388;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_26_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_26_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_26_tag <= _GEN_6170;
      end
    end else begin
      btb_26_tag <= _GEN_6170;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_26_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_26_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_26_target_address <= _GEN_10832;
      end
    end else begin
      btb_26_target_address <= _GEN_10832;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_26_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_26_bht <= 2'h1;
        end else begin
          btb_26_bht <= 2'h0;
        end
      end else begin
        btb_26_bht <= _GEN_10834;
      end
    end else begin
      btb_26_bht <= _GEN_10834;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_27_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_27_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_27_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_27_valid <= _GEN_15389;
      end
    end else begin
      btb_27_valid <= _GEN_15389;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_27_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_27_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_27_tag <= _GEN_6171;
      end
    end else begin
      btb_27_tag <= _GEN_6171;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_27_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_27_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_27_target_address <= _GEN_10835;
      end
    end else begin
      btb_27_target_address <= _GEN_10835;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_27_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_27_bht <= 2'h1;
        end else begin
          btb_27_bht <= 2'h0;
        end
      end else begin
        btb_27_bht <= _GEN_10837;
      end
    end else begin
      btb_27_bht <= _GEN_10837;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_28_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_28_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_28_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_28_valid <= _GEN_15390;
      end
    end else begin
      btb_28_valid <= _GEN_15390;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_28_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_28_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_28_tag <= _GEN_6172;
      end
    end else begin
      btb_28_tag <= _GEN_6172;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_28_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_28_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_28_target_address <= _GEN_10838;
      end
    end else begin
      btb_28_target_address <= _GEN_10838;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_28_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_28_bht <= 2'h1;
        end else begin
          btb_28_bht <= 2'h0;
        end
      end else begin
        btb_28_bht <= _GEN_10840;
      end
    end else begin
      btb_28_bht <= _GEN_10840;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_29_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_29_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_29_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_29_valid <= _GEN_15391;
      end
    end else begin
      btb_29_valid <= _GEN_15391;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_29_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_29_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_29_tag <= _GEN_6173;
      end
    end else begin
      btb_29_tag <= _GEN_6173;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_29_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_29_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_29_target_address <= _GEN_10841;
      end
    end else begin
      btb_29_target_address <= _GEN_10841;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_29_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_29_bht <= 2'h1;
        end else begin
          btb_29_bht <= 2'h0;
        end
      end else begin
        btb_29_bht <= _GEN_10843;
      end
    end else begin
      btb_29_bht <= _GEN_10843;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_30_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_30_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_30_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_30_valid <= _GEN_15392;
      end
    end else begin
      btb_30_valid <= _GEN_15392;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_30_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_30_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_30_tag <= _GEN_6174;
      end
    end else begin
      btb_30_tag <= _GEN_6174;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_30_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_30_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_30_target_address <= _GEN_10844;
      end
    end else begin
      btb_30_target_address <= _GEN_10844;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_30_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_30_bht <= 2'h1;
        end else begin
          btb_30_bht <= 2'h0;
        end
      end else begin
        btb_30_bht <= _GEN_10846;
      end
    end else begin
      btb_30_bht <= _GEN_10846;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_31_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_31_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_31_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_31_valid <= _GEN_15393;
      end
    end else begin
      btb_31_valid <= _GEN_15393;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_31_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_31_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_31_tag <= _GEN_6175;
      end
    end else begin
      btb_31_tag <= _GEN_6175;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_31_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_31_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_31_target_address <= _GEN_10847;
      end
    end else begin
      btb_31_target_address <= _GEN_10847;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_31_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_31_bht <= 2'h1;
        end else begin
          btb_31_bht <= 2'h0;
        end
      end else begin
        btb_31_bht <= _GEN_10849;
      end
    end else begin
      btb_31_bht <= _GEN_10849;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_32_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_32_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_32_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_32_valid <= _GEN_15394;
      end
    end else begin
      btb_32_valid <= _GEN_15394;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_32_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h20 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_32_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_32_tag <= _GEN_6176;
      end
    end else begin
      btb_32_tag <= _GEN_6176;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_32_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h20 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_32_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_32_target_address <= _GEN_10850;
      end
    end else begin
      btb_32_target_address <= _GEN_10850;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_32_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h20 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_32_bht <= 2'h1;
        end else begin
          btb_32_bht <= 2'h0;
        end
      end else begin
        btb_32_bht <= _GEN_10852;
      end
    end else begin
      btb_32_bht <= _GEN_10852;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_33_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_33_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_33_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_33_valid <= _GEN_15395;
      end
    end else begin
      btb_33_valid <= _GEN_15395;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_33_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h21 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_33_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_33_tag <= _GEN_6177;
      end
    end else begin
      btb_33_tag <= _GEN_6177;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_33_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h21 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_33_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_33_target_address <= _GEN_10853;
      end
    end else begin
      btb_33_target_address <= _GEN_10853;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_33_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h21 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_33_bht <= 2'h1;
        end else begin
          btb_33_bht <= 2'h0;
        end
      end else begin
        btb_33_bht <= _GEN_10855;
      end
    end else begin
      btb_33_bht <= _GEN_10855;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_34_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_34_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_34_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_34_valid <= _GEN_15396;
      end
    end else begin
      btb_34_valid <= _GEN_15396;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_34_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h22 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_34_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_34_tag <= _GEN_6178;
      end
    end else begin
      btb_34_tag <= _GEN_6178;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_34_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h22 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_34_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_34_target_address <= _GEN_10856;
      end
    end else begin
      btb_34_target_address <= _GEN_10856;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_34_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h22 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_34_bht <= 2'h1;
        end else begin
          btb_34_bht <= 2'h0;
        end
      end else begin
        btb_34_bht <= _GEN_10858;
      end
    end else begin
      btb_34_bht <= _GEN_10858;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_35_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_35_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_35_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_35_valid <= _GEN_15397;
      end
    end else begin
      btb_35_valid <= _GEN_15397;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_35_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h23 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_35_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_35_tag <= _GEN_6179;
      end
    end else begin
      btb_35_tag <= _GEN_6179;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_35_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h23 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_35_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_35_target_address <= _GEN_10859;
      end
    end else begin
      btb_35_target_address <= _GEN_10859;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_35_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h23 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_35_bht <= 2'h1;
        end else begin
          btb_35_bht <= 2'h0;
        end
      end else begin
        btb_35_bht <= _GEN_10861;
      end
    end else begin
      btb_35_bht <= _GEN_10861;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_36_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_36_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_36_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_36_valid <= _GEN_15398;
      end
    end else begin
      btb_36_valid <= _GEN_15398;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_36_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h24 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_36_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_36_tag <= _GEN_6180;
      end
    end else begin
      btb_36_tag <= _GEN_6180;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_36_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h24 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_36_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_36_target_address <= _GEN_10862;
      end
    end else begin
      btb_36_target_address <= _GEN_10862;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_36_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h24 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_36_bht <= 2'h1;
        end else begin
          btb_36_bht <= 2'h0;
        end
      end else begin
        btb_36_bht <= _GEN_10864;
      end
    end else begin
      btb_36_bht <= _GEN_10864;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_37_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_37_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_37_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_37_valid <= _GEN_15399;
      end
    end else begin
      btb_37_valid <= _GEN_15399;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_37_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h25 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_37_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_37_tag <= _GEN_6181;
      end
    end else begin
      btb_37_tag <= _GEN_6181;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_37_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h25 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_37_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_37_target_address <= _GEN_10865;
      end
    end else begin
      btb_37_target_address <= _GEN_10865;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_37_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h25 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_37_bht <= 2'h1;
        end else begin
          btb_37_bht <= 2'h0;
        end
      end else begin
        btb_37_bht <= _GEN_10867;
      end
    end else begin
      btb_37_bht <= _GEN_10867;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_38_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_38_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_38_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_38_valid <= _GEN_15400;
      end
    end else begin
      btb_38_valid <= _GEN_15400;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_38_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h26 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_38_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_38_tag <= _GEN_6182;
      end
    end else begin
      btb_38_tag <= _GEN_6182;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_38_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h26 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_38_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_38_target_address <= _GEN_10868;
      end
    end else begin
      btb_38_target_address <= _GEN_10868;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_38_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h26 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_38_bht <= 2'h1;
        end else begin
          btb_38_bht <= 2'h0;
        end
      end else begin
        btb_38_bht <= _GEN_10870;
      end
    end else begin
      btb_38_bht <= _GEN_10870;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_39_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_39_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_39_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_39_valid <= _GEN_15401;
      end
    end else begin
      btb_39_valid <= _GEN_15401;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_39_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h27 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_39_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_39_tag <= _GEN_6183;
      end
    end else begin
      btb_39_tag <= _GEN_6183;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_39_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h27 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_39_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_39_target_address <= _GEN_10871;
      end
    end else begin
      btb_39_target_address <= _GEN_10871;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_39_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h27 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_39_bht <= 2'h1;
        end else begin
          btb_39_bht <= 2'h0;
        end
      end else begin
        btb_39_bht <= _GEN_10873;
      end
    end else begin
      btb_39_bht <= _GEN_10873;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_40_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_40_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_40_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_40_valid <= _GEN_15402;
      end
    end else begin
      btb_40_valid <= _GEN_15402;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_40_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h28 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_40_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_40_tag <= _GEN_6184;
      end
    end else begin
      btb_40_tag <= _GEN_6184;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_40_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h28 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_40_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_40_target_address <= _GEN_10874;
      end
    end else begin
      btb_40_target_address <= _GEN_10874;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_40_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h28 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_40_bht <= 2'h1;
        end else begin
          btb_40_bht <= 2'h0;
        end
      end else begin
        btb_40_bht <= _GEN_10876;
      end
    end else begin
      btb_40_bht <= _GEN_10876;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_41_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_41_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_41_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_41_valid <= _GEN_15403;
      end
    end else begin
      btb_41_valid <= _GEN_15403;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_41_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h29 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_41_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_41_tag <= _GEN_6185;
      end
    end else begin
      btb_41_tag <= _GEN_6185;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_41_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h29 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_41_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_41_target_address <= _GEN_10877;
      end
    end else begin
      btb_41_target_address <= _GEN_10877;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_41_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h29 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_41_bht <= 2'h1;
        end else begin
          btb_41_bht <= 2'h0;
        end
      end else begin
        btb_41_bht <= _GEN_10879;
      end
    end else begin
      btb_41_bht <= _GEN_10879;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_42_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_42_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_42_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_42_valid <= _GEN_15404;
      end
    end else begin
      btb_42_valid <= _GEN_15404;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_42_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_42_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_42_tag <= _GEN_6186;
      end
    end else begin
      btb_42_tag <= _GEN_6186;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_42_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_42_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_42_target_address <= _GEN_10880;
      end
    end else begin
      btb_42_target_address <= _GEN_10880;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_42_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_42_bht <= 2'h1;
        end else begin
          btb_42_bht <= 2'h0;
        end
      end else begin
        btb_42_bht <= _GEN_10882;
      end
    end else begin
      btb_42_bht <= _GEN_10882;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_43_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_43_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_43_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_43_valid <= _GEN_15405;
      end
    end else begin
      btb_43_valid <= _GEN_15405;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_43_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_43_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_43_tag <= _GEN_6187;
      end
    end else begin
      btb_43_tag <= _GEN_6187;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_43_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_43_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_43_target_address <= _GEN_10883;
      end
    end else begin
      btb_43_target_address <= _GEN_10883;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_43_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_43_bht <= 2'h1;
        end else begin
          btb_43_bht <= 2'h0;
        end
      end else begin
        btb_43_bht <= _GEN_10885;
      end
    end else begin
      btb_43_bht <= _GEN_10885;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_44_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_44_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_44_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_44_valid <= _GEN_15406;
      end
    end else begin
      btb_44_valid <= _GEN_15406;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_44_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_44_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_44_tag <= _GEN_6188;
      end
    end else begin
      btb_44_tag <= _GEN_6188;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_44_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_44_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_44_target_address <= _GEN_10886;
      end
    end else begin
      btb_44_target_address <= _GEN_10886;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_44_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_44_bht <= 2'h1;
        end else begin
          btb_44_bht <= 2'h0;
        end
      end else begin
        btb_44_bht <= _GEN_10888;
      end
    end else begin
      btb_44_bht <= _GEN_10888;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_45_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_45_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_45_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_45_valid <= _GEN_15407;
      end
    end else begin
      btb_45_valid <= _GEN_15407;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_45_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_45_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_45_tag <= _GEN_6189;
      end
    end else begin
      btb_45_tag <= _GEN_6189;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_45_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_45_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_45_target_address <= _GEN_10889;
      end
    end else begin
      btb_45_target_address <= _GEN_10889;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_45_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_45_bht <= 2'h1;
        end else begin
          btb_45_bht <= 2'h0;
        end
      end else begin
        btb_45_bht <= _GEN_10891;
      end
    end else begin
      btb_45_bht <= _GEN_10891;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_46_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_46_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_46_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_46_valid <= _GEN_15408;
      end
    end else begin
      btb_46_valid <= _GEN_15408;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_46_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_46_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_46_tag <= _GEN_6190;
      end
    end else begin
      btb_46_tag <= _GEN_6190;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_46_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_46_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_46_target_address <= _GEN_10892;
      end
    end else begin
      btb_46_target_address <= _GEN_10892;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_46_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_46_bht <= 2'h1;
        end else begin
          btb_46_bht <= 2'h0;
        end
      end else begin
        btb_46_bht <= _GEN_10894;
      end
    end else begin
      btb_46_bht <= _GEN_10894;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_47_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_47_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_47_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_47_valid <= _GEN_15409;
      end
    end else begin
      btb_47_valid <= _GEN_15409;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_47_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_47_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_47_tag <= _GEN_6191;
      end
    end else begin
      btb_47_tag <= _GEN_6191;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_47_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_47_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_47_target_address <= _GEN_10895;
      end
    end else begin
      btb_47_target_address <= _GEN_10895;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_47_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h2f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_47_bht <= 2'h1;
        end else begin
          btb_47_bht <= 2'h0;
        end
      end else begin
        btb_47_bht <= _GEN_10897;
      end
    end else begin
      btb_47_bht <= _GEN_10897;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_48_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_48_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_48_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_48_valid <= _GEN_15410;
      end
    end else begin
      btb_48_valid <= _GEN_15410;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_48_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h30 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_48_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_48_tag <= _GEN_6192;
      end
    end else begin
      btb_48_tag <= _GEN_6192;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_48_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h30 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_48_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_48_target_address <= _GEN_10898;
      end
    end else begin
      btb_48_target_address <= _GEN_10898;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_48_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h30 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_48_bht <= 2'h1;
        end else begin
          btb_48_bht <= 2'h0;
        end
      end else begin
        btb_48_bht <= _GEN_10900;
      end
    end else begin
      btb_48_bht <= _GEN_10900;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_49_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_49_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_49_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_49_valid <= _GEN_15411;
      end
    end else begin
      btb_49_valid <= _GEN_15411;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_49_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h31 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_49_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_49_tag <= _GEN_6193;
      end
    end else begin
      btb_49_tag <= _GEN_6193;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_49_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h31 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_49_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_49_target_address <= _GEN_10901;
      end
    end else begin
      btb_49_target_address <= _GEN_10901;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_49_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h31 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_49_bht <= 2'h1;
        end else begin
          btb_49_bht <= 2'h0;
        end
      end else begin
        btb_49_bht <= _GEN_10903;
      end
    end else begin
      btb_49_bht <= _GEN_10903;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_50_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_50_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_50_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_50_valid <= _GEN_15412;
      end
    end else begin
      btb_50_valid <= _GEN_15412;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_50_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h32 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_50_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_50_tag <= _GEN_6194;
      end
    end else begin
      btb_50_tag <= _GEN_6194;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_50_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h32 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_50_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_50_target_address <= _GEN_10904;
      end
    end else begin
      btb_50_target_address <= _GEN_10904;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_50_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h32 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_50_bht <= 2'h1;
        end else begin
          btb_50_bht <= 2'h0;
        end
      end else begin
        btb_50_bht <= _GEN_10906;
      end
    end else begin
      btb_50_bht <= _GEN_10906;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_51_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_51_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_51_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_51_valid <= _GEN_15413;
      end
    end else begin
      btb_51_valid <= _GEN_15413;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_51_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h33 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_51_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_51_tag <= _GEN_6195;
      end
    end else begin
      btb_51_tag <= _GEN_6195;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_51_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h33 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_51_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_51_target_address <= _GEN_10907;
      end
    end else begin
      btb_51_target_address <= _GEN_10907;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_51_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h33 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_51_bht <= 2'h1;
        end else begin
          btb_51_bht <= 2'h0;
        end
      end else begin
        btb_51_bht <= _GEN_10909;
      end
    end else begin
      btb_51_bht <= _GEN_10909;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_52_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_52_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_52_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_52_valid <= _GEN_15414;
      end
    end else begin
      btb_52_valid <= _GEN_15414;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_52_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h34 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_52_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_52_tag <= _GEN_6196;
      end
    end else begin
      btb_52_tag <= _GEN_6196;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_52_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h34 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_52_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_52_target_address <= _GEN_10910;
      end
    end else begin
      btb_52_target_address <= _GEN_10910;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_52_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h34 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_52_bht <= 2'h1;
        end else begin
          btb_52_bht <= 2'h0;
        end
      end else begin
        btb_52_bht <= _GEN_10912;
      end
    end else begin
      btb_52_bht <= _GEN_10912;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_53_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_53_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_53_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_53_valid <= _GEN_15415;
      end
    end else begin
      btb_53_valid <= _GEN_15415;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_53_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h35 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_53_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_53_tag <= _GEN_6197;
      end
    end else begin
      btb_53_tag <= _GEN_6197;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_53_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h35 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_53_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_53_target_address <= _GEN_10913;
      end
    end else begin
      btb_53_target_address <= _GEN_10913;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_53_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h35 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_53_bht <= 2'h1;
        end else begin
          btb_53_bht <= 2'h0;
        end
      end else begin
        btb_53_bht <= _GEN_10915;
      end
    end else begin
      btb_53_bht <= _GEN_10915;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_54_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_54_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_54_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_54_valid <= _GEN_15416;
      end
    end else begin
      btb_54_valid <= _GEN_15416;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_54_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h36 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_54_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_54_tag <= _GEN_6198;
      end
    end else begin
      btb_54_tag <= _GEN_6198;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_54_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h36 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_54_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_54_target_address <= _GEN_10916;
      end
    end else begin
      btb_54_target_address <= _GEN_10916;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_54_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h36 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_54_bht <= 2'h1;
        end else begin
          btb_54_bht <= 2'h0;
        end
      end else begin
        btb_54_bht <= _GEN_10918;
      end
    end else begin
      btb_54_bht <= _GEN_10918;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_55_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_55_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_55_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_55_valid <= _GEN_15417;
      end
    end else begin
      btb_55_valid <= _GEN_15417;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_55_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h37 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_55_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_55_tag <= _GEN_6199;
      end
    end else begin
      btb_55_tag <= _GEN_6199;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_55_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h37 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_55_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_55_target_address <= _GEN_10919;
      end
    end else begin
      btb_55_target_address <= _GEN_10919;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_55_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h37 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_55_bht <= 2'h1;
        end else begin
          btb_55_bht <= 2'h0;
        end
      end else begin
        btb_55_bht <= _GEN_10921;
      end
    end else begin
      btb_55_bht <= _GEN_10921;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_56_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_56_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_56_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_56_valid <= _GEN_15418;
      end
    end else begin
      btb_56_valid <= _GEN_15418;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_56_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h38 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_56_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_56_tag <= _GEN_6200;
      end
    end else begin
      btb_56_tag <= _GEN_6200;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_56_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h38 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_56_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_56_target_address <= _GEN_10922;
      end
    end else begin
      btb_56_target_address <= _GEN_10922;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_56_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h38 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_56_bht <= 2'h1;
        end else begin
          btb_56_bht <= 2'h0;
        end
      end else begin
        btb_56_bht <= _GEN_10924;
      end
    end else begin
      btb_56_bht <= _GEN_10924;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_57_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_57_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_57_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_57_valid <= _GEN_15419;
      end
    end else begin
      btb_57_valid <= _GEN_15419;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_57_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h39 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_57_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_57_tag <= _GEN_6201;
      end
    end else begin
      btb_57_tag <= _GEN_6201;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_57_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h39 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_57_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_57_target_address <= _GEN_10925;
      end
    end else begin
      btb_57_target_address <= _GEN_10925;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_57_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h39 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_57_bht <= 2'h1;
        end else begin
          btb_57_bht <= 2'h0;
        end
      end else begin
        btb_57_bht <= _GEN_10927;
      end
    end else begin
      btb_57_bht <= _GEN_10927;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_58_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_58_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_58_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_58_valid <= _GEN_15420;
      end
    end else begin
      btb_58_valid <= _GEN_15420;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_58_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_58_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_58_tag <= _GEN_6202;
      end
    end else begin
      btb_58_tag <= _GEN_6202;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_58_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_58_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_58_target_address <= _GEN_10928;
      end
    end else begin
      btb_58_target_address <= _GEN_10928;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_58_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_58_bht <= 2'h1;
        end else begin
          btb_58_bht <= 2'h0;
        end
      end else begin
        btb_58_bht <= _GEN_10930;
      end
    end else begin
      btb_58_bht <= _GEN_10930;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_59_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_59_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_59_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_59_valid <= _GEN_15421;
      end
    end else begin
      btb_59_valid <= _GEN_15421;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_59_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_59_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_59_tag <= _GEN_6203;
      end
    end else begin
      btb_59_tag <= _GEN_6203;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_59_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_59_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_59_target_address <= _GEN_10931;
      end
    end else begin
      btb_59_target_address <= _GEN_10931;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_59_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_59_bht <= 2'h1;
        end else begin
          btb_59_bht <= 2'h0;
        end
      end else begin
        btb_59_bht <= _GEN_10933;
      end
    end else begin
      btb_59_bht <= _GEN_10933;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_60_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_60_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_60_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_60_valid <= _GEN_15422;
      end
    end else begin
      btb_60_valid <= _GEN_15422;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_60_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_60_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_60_tag <= _GEN_6204;
      end
    end else begin
      btb_60_tag <= _GEN_6204;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_60_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_60_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_60_target_address <= _GEN_10934;
      end
    end else begin
      btb_60_target_address <= _GEN_10934;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_60_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_60_bht <= 2'h1;
        end else begin
          btb_60_bht <= 2'h0;
        end
      end else begin
        btb_60_bht <= _GEN_10936;
      end
    end else begin
      btb_60_bht <= _GEN_10936;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_61_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_61_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_61_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_61_valid <= _GEN_15423;
      end
    end else begin
      btb_61_valid <= _GEN_15423;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_61_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_61_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_61_tag <= _GEN_6205;
      end
    end else begin
      btb_61_tag <= _GEN_6205;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_61_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_61_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_61_target_address <= _GEN_10937;
      end
    end else begin
      btb_61_target_address <= _GEN_10937;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_61_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_61_bht <= 2'h1;
        end else begin
          btb_61_bht <= 2'h0;
        end
      end else begin
        btb_61_bht <= _GEN_10939;
      end
    end else begin
      btb_61_bht <= _GEN_10939;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_62_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_62_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_62_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_62_valid <= _GEN_15424;
      end
    end else begin
      btb_62_valid <= _GEN_15424;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_62_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_62_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_62_tag <= _GEN_6206;
      end
    end else begin
      btb_62_tag <= _GEN_6206;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_62_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_62_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_62_target_address <= _GEN_10940;
      end
    end else begin
      btb_62_target_address <= _GEN_10940;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_62_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_62_bht <= 2'h1;
        end else begin
          btb_62_bht <= 2'h0;
        end
      end else begin
        btb_62_bht <= _GEN_10942;
      end
    end else begin
      btb_62_bht <= _GEN_10942;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_63_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_63_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_63_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_63_valid <= _GEN_15425;
      end
    end else begin
      btb_63_valid <= _GEN_15425;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_63_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_63_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_63_tag <= _GEN_6207;
      end
    end else begin
      btb_63_tag <= _GEN_6207;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_63_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_63_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_63_target_address <= _GEN_10943;
      end
    end else begin
      btb_63_target_address <= _GEN_10943;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_63_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h3f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_63_bht <= 2'h1;
        end else begin
          btb_63_bht <= 2'h0;
        end
      end else begin
        btb_63_bht <= _GEN_10945;
      end
    end else begin
      btb_63_bht <= _GEN_10945;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_64_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_64_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_64_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_64_valid <= _GEN_15426;
      end
    end else begin
      btb_64_valid <= _GEN_15426;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_64_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h40 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_64_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_64_tag <= _GEN_6208;
      end
    end else begin
      btb_64_tag <= _GEN_6208;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_64_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h40 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_64_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_64_target_address <= _GEN_10946;
      end
    end else begin
      btb_64_target_address <= _GEN_10946;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_64_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h40 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_64_bht <= 2'h1;
        end else begin
          btb_64_bht <= 2'h0;
        end
      end else begin
        btb_64_bht <= _GEN_10948;
      end
    end else begin
      btb_64_bht <= _GEN_10948;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_65_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_65_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_65_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_65_valid <= _GEN_15427;
      end
    end else begin
      btb_65_valid <= _GEN_15427;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_65_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h41 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_65_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_65_tag <= _GEN_6209;
      end
    end else begin
      btb_65_tag <= _GEN_6209;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_65_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h41 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_65_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_65_target_address <= _GEN_10949;
      end
    end else begin
      btb_65_target_address <= _GEN_10949;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_65_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h41 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_65_bht <= 2'h1;
        end else begin
          btb_65_bht <= 2'h0;
        end
      end else begin
        btb_65_bht <= _GEN_10951;
      end
    end else begin
      btb_65_bht <= _GEN_10951;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_66_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_66_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_66_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_66_valid <= _GEN_15428;
      end
    end else begin
      btb_66_valid <= _GEN_15428;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_66_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h42 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_66_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_66_tag <= _GEN_6210;
      end
    end else begin
      btb_66_tag <= _GEN_6210;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_66_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h42 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_66_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_66_target_address <= _GEN_10952;
      end
    end else begin
      btb_66_target_address <= _GEN_10952;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_66_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h42 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_66_bht <= 2'h1;
        end else begin
          btb_66_bht <= 2'h0;
        end
      end else begin
        btb_66_bht <= _GEN_10954;
      end
    end else begin
      btb_66_bht <= _GEN_10954;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_67_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_67_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_67_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_67_valid <= _GEN_15429;
      end
    end else begin
      btb_67_valid <= _GEN_15429;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_67_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h43 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_67_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_67_tag <= _GEN_6211;
      end
    end else begin
      btb_67_tag <= _GEN_6211;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_67_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h43 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_67_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_67_target_address <= _GEN_10955;
      end
    end else begin
      btb_67_target_address <= _GEN_10955;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_67_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h43 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_67_bht <= 2'h1;
        end else begin
          btb_67_bht <= 2'h0;
        end
      end else begin
        btb_67_bht <= _GEN_10957;
      end
    end else begin
      btb_67_bht <= _GEN_10957;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_68_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_68_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_68_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_68_valid <= _GEN_15430;
      end
    end else begin
      btb_68_valid <= _GEN_15430;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_68_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h44 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_68_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_68_tag <= _GEN_6212;
      end
    end else begin
      btb_68_tag <= _GEN_6212;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_68_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h44 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_68_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_68_target_address <= _GEN_10958;
      end
    end else begin
      btb_68_target_address <= _GEN_10958;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_68_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h44 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_68_bht <= 2'h1;
        end else begin
          btb_68_bht <= 2'h0;
        end
      end else begin
        btb_68_bht <= _GEN_10960;
      end
    end else begin
      btb_68_bht <= _GEN_10960;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_69_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_69_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_69_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_69_valid <= _GEN_15431;
      end
    end else begin
      btb_69_valid <= _GEN_15431;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_69_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h45 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_69_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_69_tag <= _GEN_6213;
      end
    end else begin
      btb_69_tag <= _GEN_6213;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_69_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h45 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_69_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_69_target_address <= _GEN_10961;
      end
    end else begin
      btb_69_target_address <= _GEN_10961;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_69_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h45 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_69_bht <= 2'h1;
        end else begin
          btb_69_bht <= 2'h0;
        end
      end else begin
        btb_69_bht <= _GEN_10963;
      end
    end else begin
      btb_69_bht <= _GEN_10963;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_70_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_70_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_70_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_70_valid <= _GEN_15432;
      end
    end else begin
      btb_70_valid <= _GEN_15432;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_70_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h46 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_70_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_70_tag <= _GEN_6214;
      end
    end else begin
      btb_70_tag <= _GEN_6214;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_70_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h46 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_70_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_70_target_address <= _GEN_10964;
      end
    end else begin
      btb_70_target_address <= _GEN_10964;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_70_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h46 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_70_bht <= 2'h1;
        end else begin
          btb_70_bht <= 2'h0;
        end
      end else begin
        btb_70_bht <= _GEN_10966;
      end
    end else begin
      btb_70_bht <= _GEN_10966;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_71_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_71_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_71_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_71_valid <= _GEN_15433;
      end
    end else begin
      btb_71_valid <= _GEN_15433;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_71_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h47 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_71_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_71_tag <= _GEN_6215;
      end
    end else begin
      btb_71_tag <= _GEN_6215;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_71_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h47 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_71_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_71_target_address <= _GEN_10967;
      end
    end else begin
      btb_71_target_address <= _GEN_10967;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_71_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h47 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_71_bht <= 2'h1;
        end else begin
          btb_71_bht <= 2'h0;
        end
      end else begin
        btb_71_bht <= _GEN_10969;
      end
    end else begin
      btb_71_bht <= _GEN_10969;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_72_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_72_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_72_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_72_valid <= _GEN_15434;
      end
    end else begin
      btb_72_valid <= _GEN_15434;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_72_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h48 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_72_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_72_tag <= _GEN_6216;
      end
    end else begin
      btb_72_tag <= _GEN_6216;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_72_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h48 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_72_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_72_target_address <= _GEN_10970;
      end
    end else begin
      btb_72_target_address <= _GEN_10970;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_72_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h48 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_72_bht <= 2'h1;
        end else begin
          btb_72_bht <= 2'h0;
        end
      end else begin
        btb_72_bht <= _GEN_10972;
      end
    end else begin
      btb_72_bht <= _GEN_10972;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_73_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_73_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_73_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_73_valid <= _GEN_15435;
      end
    end else begin
      btb_73_valid <= _GEN_15435;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_73_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h49 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_73_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_73_tag <= _GEN_6217;
      end
    end else begin
      btb_73_tag <= _GEN_6217;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_73_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h49 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_73_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_73_target_address <= _GEN_10973;
      end
    end else begin
      btb_73_target_address <= _GEN_10973;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_73_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h49 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_73_bht <= 2'h1;
        end else begin
          btb_73_bht <= 2'h0;
        end
      end else begin
        btb_73_bht <= _GEN_10975;
      end
    end else begin
      btb_73_bht <= _GEN_10975;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_74_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_74_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_74_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_74_valid <= _GEN_15436;
      end
    end else begin
      btb_74_valid <= _GEN_15436;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_74_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_74_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_74_tag <= _GEN_6218;
      end
    end else begin
      btb_74_tag <= _GEN_6218;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_74_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_74_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_74_target_address <= _GEN_10976;
      end
    end else begin
      btb_74_target_address <= _GEN_10976;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_74_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_74_bht <= 2'h1;
        end else begin
          btb_74_bht <= 2'h0;
        end
      end else begin
        btb_74_bht <= _GEN_10978;
      end
    end else begin
      btb_74_bht <= _GEN_10978;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_75_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_75_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_75_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_75_valid <= _GEN_15437;
      end
    end else begin
      btb_75_valid <= _GEN_15437;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_75_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_75_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_75_tag <= _GEN_6219;
      end
    end else begin
      btb_75_tag <= _GEN_6219;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_75_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_75_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_75_target_address <= _GEN_10979;
      end
    end else begin
      btb_75_target_address <= _GEN_10979;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_75_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_75_bht <= 2'h1;
        end else begin
          btb_75_bht <= 2'h0;
        end
      end else begin
        btb_75_bht <= _GEN_10981;
      end
    end else begin
      btb_75_bht <= _GEN_10981;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_76_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_76_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_76_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_76_valid <= _GEN_15438;
      end
    end else begin
      btb_76_valid <= _GEN_15438;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_76_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_76_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_76_tag <= _GEN_6220;
      end
    end else begin
      btb_76_tag <= _GEN_6220;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_76_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_76_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_76_target_address <= _GEN_10982;
      end
    end else begin
      btb_76_target_address <= _GEN_10982;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_76_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_76_bht <= 2'h1;
        end else begin
          btb_76_bht <= 2'h0;
        end
      end else begin
        btb_76_bht <= _GEN_10984;
      end
    end else begin
      btb_76_bht <= _GEN_10984;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_77_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_77_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_77_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_77_valid <= _GEN_15439;
      end
    end else begin
      btb_77_valid <= _GEN_15439;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_77_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_77_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_77_tag <= _GEN_6221;
      end
    end else begin
      btb_77_tag <= _GEN_6221;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_77_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_77_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_77_target_address <= _GEN_10985;
      end
    end else begin
      btb_77_target_address <= _GEN_10985;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_77_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_77_bht <= 2'h1;
        end else begin
          btb_77_bht <= 2'h0;
        end
      end else begin
        btb_77_bht <= _GEN_10987;
      end
    end else begin
      btb_77_bht <= _GEN_10987;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_78_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_78_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_78_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_78_valid <= _GEN_15440;
      end
    end else begin
      btb_78_valid <= _GEN_15440;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_78_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_78_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_78_tag <= _GEN_6222;
      end
    end else begin
      btb_78_tag <= _GEN_6222;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_78_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_78_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_78_target_address <= _GEN_10988;
      end
    end else begin
      btb_78_target_address <= _GEN_10988;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_78_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_78_bht <= 2'h1;
        end else begin
          btb_78_bht <= 2'h0;
        end
      end else begin
        btb_78_bht <= _GEN_10990;
      end
    end else begin
      btb_78_bht <= _GEN_10990;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_79_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_79_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_79_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_79_valid <= _GEN_15441;
      end
    end else begin
      btb_79_valid <= _GEN_15441;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_79_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_79_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_79_tag <= _GEN_6223;
      end
    end else begin
      btb_79_tag <= _GEN_6223;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_79_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_79_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_79_target_address <= _GEN_10991;
      end
    end else begin
      btb_79_target_address <= _GEN_10991;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_79_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h4f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_79_bht <= 2'h1;
        end else begin
          btb_79_bht <= 2'h0;
        end
      end else begin
        btb_79_bht <= _GEN_10993;
      end
    end else begin
      btb_79_bht <= _GEN_10993;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_80_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_80_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_80_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_80_valid <= _GEN_15442;
      end
    end else begin
      btb_80_valid <= _GEN_15442;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_80_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h50 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_80_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_80_tag <= _GEN_6224;
      end
    end else begin
      btb_80_tag <= _GEN_6224;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_80_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h50 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_80_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_80_target_address <= _GEN_10994;
      end
    end else begin
      btb_80_target_address <= _GEN_10994;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_80_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h50 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_80_bht <= 2'h1;
        end else begin
          btb_80_bht <= 2'h0;
        end
      end else begin
        btb_80_bht <= _GEN_10996;
      end
    end else begin
      btb_80_bht <= _GEN_10996;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_81_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_81_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_81_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_81_valid <= _GEN_15443;
      end
    end else begin
      btb_81_valid <= _GEN_15443;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_81_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h51 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_81_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_81_tag <= _GEN_6225;
      end
    end else begin
      btb_81_tag <= _GEN_6225;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_81_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h51 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_81_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_81_target_address <= _GEN_10997;
      end
    end else begin
      btb_81_target_address <= _GEN_10997;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_81_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h51 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_81_bht <= 2'h1;
        end else begin
          btb_81_bht <= 2'h0;
        end
      end else begin
        btb_81_bht <= _GEN_10999;
      end
    end else begin
      btb_81_bht <= _GEN_10999;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_82_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_82_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_82_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_82_valid <= _GEN_15444;
      end
    end else begin
      btb_82_valid <= _GEN_15444;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_82_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h52 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_82_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_82_tag <= _GEN_6226;
      end
    end else begin
      btb_82_tag <= _GEN_6226;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_82_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h52 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_82_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_82_target_address <= _GEN_11000;
      end
    end else begin
      btb_82_target_address <= _GEN_11000;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_82_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h52 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_82_bht <= 2'h1;
        end else begin
          btb_82_bht <= 2'h0;
        end
      end else begin
        btb_82_bht <= _GEN_11002;
      end
    end else begin
      btb_82_bht <= _GEN_11002;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_83_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_83_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_83_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_83_valid <= _GEN_15445;
      end
    end else begin
      btb_83_valid <= _GEN_15445;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_83_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h53 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_83_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_83_tag <= _GEN_6227;
      end
    end else begin
      btb_83_tag <= _GEN_6227;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_83_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h53 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_83_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_83_target_address <= _GEN_11003;
      end
    end else begin
      btb_83_target_address <= _GEN_11003;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_83_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h53 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_83_bht <= 2'h1;
        end else begin
          btb_83_bht <= 2'h0;
        end
      end else begin
        btb_83_bht <= _GEN_11005;
      end
    end else begin
      btb_83_bht <= _GEN_11005;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_84_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_84_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_84_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_84_valid <= _GEN_15446;
      end
    end else begin
      btb_84_valid <= _GEN_15446;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_84_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h54 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_84_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_84_tag <= _GEN_6228;
      end
    end else begin
      btb_84_tag <= _GEN_6228;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_84_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h54 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_84_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_84_target_address <= _GEN_11006;
      end
    end else begin
      btb_84_target_address <= _GEN_11006;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_84_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h54 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_84_bht <= 2'h1;
        end else begin
          btb_84_bht <= 2'h0;
        end
      end else begin
        btb_84_bht <= _GEN_11008;
      end
    end else begin
      btb_84_bht <= _GEN_11008;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_85_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_85_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_85_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_85_valid <= _GEN_15447;
      end
    end else begin
      btb_85_valid <= _GEN_15447;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_85_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h55 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_85_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_85_tag <= _GEN_6229;
      end
    end else begin
      btb_85_tag <= _GEN_6229;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_85_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h55 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_85_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_85_target_address <= _GEN_11009;
      end
    end else begin
      btb_85_target_address <= _GEN_11009;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_85_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h55 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_85_bht <= 2'h1;
        end else begin
          btb_85_bht <= 2'h0;
        end
      end else begin
        btb_85_bht <= _GEN_11011;
      end
    end else begin
      btb_85_bht <= _GEN_11011;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_86_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_86_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_86_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_86_valid <= _GEN_15448;
      end
    end else begin
      btb_86_valid <= _GEN_15448;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_86_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h56 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_86_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_86_tag <= _GEN_6230;
      end
    end else begin
      btb_86_tag <= _GEN_6230;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_86_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h56 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_86_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_86_target_address <= _GEN_11012;
      end
    end else begin
      btb_86_target_address <= _GEN_11012;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_86_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h56 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_86_bht <= 2'h1;
        end else begin
          btb_86_bht <= 2'h0;
        end
      end else begin
        btb_86_bht <= _GEN_11014;
      end
    end else begin
      btb_86_bht <= _GEN_11014;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_87_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_87_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_87_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_87_valid <= _GEN_15449;
      end
    end else begin
      btb_87_valid <= _GEN_15449;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_87_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h57 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_87_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_87_tag <= _GEN_6231;
      end
    end else begin
      btb_87_tag <= _GEN_6231;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_87_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h57 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_87_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_87_target_address <= _GEN_11015;
      end
    end else begin
      btb_87_target_address <= _GEN_11015;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_87_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h57 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_87_bht <= 2'h1;
        end else begin
          btb_87_bht <= 2'h0;
        end
      end else begin
        btb_87_bht <= _GEN_11017;
      end
    end else begin
      btb_87_bht <= _GEN_11017;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_88_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_88_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_88_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_88_valid <= _GEN_15450;
      end
    end else begin
      btb_88_valid <= _GEN_15450;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_88_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h58 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_88_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_88_tag <= _GEN_6232;
      end
    end else begin
      btb_88_tag <= _GEN_6232;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_88_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h58 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_88_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_88_target_address <= _GEN_11018;
      end
    end else begin
      btb_88_target_address <= _GEN_11018;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_88_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h58 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_88_bht <= 2'h1;
        end else begin
          btb_88_bht <= 2'h0;
        end
      end else begin
        btb_88_bht <= _GEN_11020;
      end
    end else begin
      btb_88_bht <= _GEN_11020;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_89_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_89_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_89_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_89_valid <= _GEN_15451;
      end
    end else begin
      btb_89_valid <= _GEN_15451;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_89_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h59 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_89_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_89_tag <= _GEN_6233;
      end
    end else begin
      btb_89_tag <= _GEN_6233;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_89_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h59 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_89_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_89_target_address <= _GEN_11021;
      end
    end else begin
      btb_89_target_address <= _GEN_11021;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_89_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h59 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_89_bht <= 2'h1;
        end else begin
          btb_89_bht <= 2'h0;
        end
      end else begin
        btb_89_bht <= _GEN_11023;
      end
    end else begin
      btb_89_bht <= _GEN_11023;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_90_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_90_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_90_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_90_valid <= _GEN_15452;
      end
    end else begin
      btb_90_valid <= _GEN_15452;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_90_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_90_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_90_tag <= _GEN_6234;
      end
    end else begin
      btb_90_tag <= _GEN_6234;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_90_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_90_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_90_target_address <= _GEN_11024;
      end
    end else begin
      btb_90_target_address <= _GEN_11024;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_90_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_90_bht <= 2'h1;
        end else begin
          btb_90_bht <= 2'h0;
        end
      end else begin
        btb_90_bht <= _GEN_11026;
      end
    end else begin
      btb_90_bht <= _GEN_11026;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_91_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_91_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_91_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_91_valid <= _GEN_15453;
      end
    end else begin
      btb_91_valid <= _GEN_15453;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_91_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_91_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_91_tag <= _GEN_6235;
      end
    end else begin
      btb_91_tag <= _GEN_6235;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_91_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_91_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_91_target_address <= _GEN_11027;
      end
    end else begin
      btb_91_target_address <= _GEN_11027;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_91_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_91_bht <= 2'h1;
        end else begin
          btb_91_bht <= 2'h0;
        end
      end else begin
        btb_91_bht <= _GEN_11029;
      end
    end else begin
      btb_91_bht <= _GEN_11029;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_92_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_92_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_92_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_92_valid <= _GEN_15454;
      end
    end else begin
      btb_92_valid <= _GEN_15454;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_92_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_92_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_92_tag <= _GEN_6236;
      end
    end else begin
      btb_92_tag <= _GEN_6236;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_92_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_92_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_92_target_address <= _GEN_11030;
      end
    end else begin
      btb_92_target_address <= _GEN_11030;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_92_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_92_bht <= 2'h1;
        end else begin
          btb_92_bht <= 2'h0;
        end
      end else begin
        btb_92_bht <= _GEN_11032;
      end
    end else begin
      btb_92_bht <= _GEN_11032;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_93_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_93_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_93_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_93_valid <= _GEN_15455;
      end
    end else begin
      btb_93_valid <= _GEN_15455;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_93_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_93_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_93_tag <= _GEN_6237;
      end
    end else begin
      btb_93_tag <= _GEN_6237;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_93_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_93_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_93_target_address <= _GEN_11033;
      end
    end else begin
      btb_93_target_address <= _GEN_11033;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_93_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_93_bht <= 2'h1;
        end else begin
          btb_93_bht <= 2'h0;
        end
      end else begin
        btb_93_bht <= _GEN_11035;
      end
    end else begin
      btb_93_bht <= _GEN_11035;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_94_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_94_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_94_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_94_valid <= _GEN_15456;
      end
    end else begin
      btb_94_valid <= _GEN_15456;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_94_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_94_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_94_tag <= _GEN_6238;
      end
    end else begin
      btb_94_tag <= _GEN_6238;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_94_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_94_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_94_target_address <= _GEN_11036;
      end
    end else begin
      btb_94_target_address <= _GEN_11036;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_94_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_94_bht <= 2'h1;
        end else begin
          btb_94_bht <= 2'h0;
        end
      end else begin
        btb_94_bht <= _GEN_11038;
      end
    end else begin
      btb_94_bht <= _GEN_11038;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_95_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_95_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_95_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_95_valid <= _GEN_15457;
      end
    end else begin
      btb_95_valid <= _GEN_15457;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_95_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_95_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_95_tag <= _GEN_6239;
      end
    end else begin
      btb_95_tag <= _GEN_6239;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_95_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_95_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_95_target_address <= _GEN_11039;
      end
    end else begin
      btb_95_target_address <= _GEN_11039;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_95_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h5f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_95_bht <= 2'h1;
        end else begin
          btb_95_bht <= 2'h0;
        end
      end else begin
        btb_95_bht <= _GEN_11041;
      end
    end else begin
      btb_95_bht <= _GEN_11041;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_96_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_96_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_96_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_96_valid <= _GEN_15458;
      end
    end else begin
      btb_96_valid <= _GEN_15458;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_96_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h60 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_96_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_96_tag <= _GEN_6240;
      end
    end else begin
      btb_96_tag <= _GEN_6240;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_96_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h60 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_96_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_96_target_address <= _GEN_11042;
      end
    end else begin
      btb_96_target_address <= _GEN_11042;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_96_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h60 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_96_bht <= 2'h1;
        end else begin
          btb_96_bht <= 2'h0;
        end
      end else begin
        btb_96_bht <= _GEN_11044;
      end
    end else begin
      btb_96_bht <= _GEN_11044;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_97_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_97_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_97_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_97_valid <= _GEN_15459;
      end
    end else begin
      btb_97_valid <= _GEN_15459;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_97_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h61 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_97_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_97_tag <= _GEN_6241;
      end
    end else begin
      btb_97_tag <= _GEN_6241;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_97_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h61 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_97_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_97_target_address <= _GEN_11045;
      end
    end else begin
      btb_97_target_address <= _GEN_11045;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_97_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h61 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_97_bht <= 2'h1;
        end else begin
          btb_97_bht <= 2'h0;
        end
      end else begin
        btb_97_bht <= _GEN_11047;
      end
    end else begin
      btb_97_bht <= _GEN_11047;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_98_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_98_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_98_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_98_valid <= _GEN_15460;
      end
    end else begin
      btb_98_valid <= _GEN_15460;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_98_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h62 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_98_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_98_tag <= _GEN_6242;
      end
    end else begin
      btb_98_tag <= _GEN_6242;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_98_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h62 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_98_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_98_target_address <= _GEN_11048;
      end
    end else begin
      btb_98_target_address <= _GEN_11048;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_98_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h62 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_98_bht <= 2'h1;
        end else begin
          btb_98_bht <= 2'h0;
        end
      end else begin
        btb_98_bht <= _GEN_11050;
      end
    end else begin
      btb_98_bht <= _GEN_11050;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_99_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_99_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_99_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_99_valid <= _GEN_15461;
      end
    end else begin
      btb_99_valid <= _GEN_15461;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_99_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h63 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_99_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_99_tag <= _GEN_6243;
      end
    end else begin
      btb_99_tag <= _GEN_6243;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_99_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h63 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_99_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_99_target_address <= _GEN_11051;
      end
    end else begin
      btb_99_target_address <= _GEN_11051;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_99_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h63 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_99_bht <= 2'h1;
        end else begin
          btb_99_bht <= 2'h0;
        end
      end else begin
        btb_99_bht <= _GEN_11053;
      end
    end else begin
      btb_99_bht <= _GEN_11053;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_100_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_100_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_100_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_100_valid <= _GEN_15462;
      end
    end else begin
      btb_100_valid <= _GEN_15462;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_100_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h64 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_100_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_100_tag <= _GEN_6244;
      end
    end else begin
      btb_100_tag <= _GEN_6244;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_100_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h64 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_100_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_100_target_address <= _GEN_11054;
      end
    end else begin
      btb_100_target_address <= _GEN_11054;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_100_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h64 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_100_bht <= 2'h1;
        end else begin
          btb_100_bht <= 2'h0;
        end
      end else begin
        btb_100_bht <= _GEN_11056;
      end
    end else begin
      btb_100_bht <= _GEN_11056;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_101_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_101_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_101_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_101_valid <= _GEN_15463;
      end
    end else begin
      btb_101_valid <= _GEN_15463;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_101_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h65 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_101_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_101_tag <= _GEN_6245;
      end
    end else begin
      btb_101_tag <= _GEN_6245;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_101_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h65 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_101_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_101_target_address <= _GEN_11057;
      end
    end else begin
      btb_101_target_address <= _GEN_11057;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_101_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h65 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_101_bht <= 2'h1;
        end else begin
          btb_101_bht <= 2'h0;
        end
      end else begin
        btb_101_bht <= _GEN_11059;
      end
    end else begin
      btb_101_bht <= _GEN_11059;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_102_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_102_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_102_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_102_valid <= _GEN_15464;
      end
    end else begin
      btb_102_valid <= _GEN_15464;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_102_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h66 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_102_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_102_tag <= _GEN_6246;
      end
    end else begin
      btb_102_tag <= _GEN_6246;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_102_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h66 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_102_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_102_target_address <= _GEN_11060;
      end
    end else begin
      btb_102_target_address <= _GEN_11060;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_102_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h66 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_102_bht <= 2'h1;
        end else begin
          btb_102_bht <= 2'h0;
        end
      end else begin
        btb_102_bht <= _GEN_11062;
      end
    end else begin
      btb_102_bht <= _GEN_11062;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_103_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_103_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_103_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_103_valid <= _GEN_15465;
      end
    end else begin
      btb_103_valid <= _GEN_15465;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_103_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h67 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_103_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_103_tag <= _GEN_6247;
      end
    end else begin
      btb_103_tag <= _GEN_6247;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_103_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h67 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_103_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_103_target_address <= _GEN_11063;
      end
    end else begin
      btb_103_target_address <= _GEN_11063;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_103_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h67 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_103_bht <= 2'h1;
        end else begin
          btb_103_bht <= 2'h0;
        end
      end else begin
        btb_103_bht <= _GEN_11065;
      end
    end else begin
      btb_103_bht <= _GEN_11065;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_104_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_104_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_104_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_104_valid <= _GEN_15466;
      end
    end else begin
      btb_104_valid <= _GEN_15466;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_104_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h68 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_104_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_104_tag <= _GEN_6248;
      end
    end else begin
      btb_104_tag <= _GEN_6248;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_104_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h68 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_104_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_104_target_address <= _GEN_11066;
      end
    end else begin
      btb_104_target_address <= _GEN_11066;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_104_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h68 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_104_bht <= 2'h1;
        end else begin
          btb_104_bht <= 2'h0;
        end
      end else begin
        btb_104_bht <= _GEN_11068;
      end
    end else begin
      btb_104_bht <= _GEN_11068;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_105_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_105_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_105_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_105_valid <= _GEN_15467;
      end
    end else begin
      btb_105_valid <= _GEN_15467;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_105_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h69 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_105_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_105_tag <= _GEN_6249;
      end
    end else begin
      btb_105_tag <= _GEN_6249;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_105_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h69 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_105_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_105_target_address <= _GEN_11069;
      end
    end else begin
      btb_105_target_address <= _GEN_11069;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_105_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h69 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_105_bht <= 2'h1;
        end else begin
          btb_105_bht <= 2'h0;
        end
      end else begin
        btb_105_bht <= _GEN_11071;
      end
    end else begin
      btb_105_bht <= _GEN_11071;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_106_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_106_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_106_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_106_valid <= _GEN_15468;
      end
    end else begin
      btb_106_valid <= _GEN_15468;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_106_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_106_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_106_tag <= _GEN_6250;
      end
    end else begin
      btb_106_tag <= _GEN_6250;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_106_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_106_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_106_target_address <= _GEN_11072;
      end
    end else begin
      btb_106_target_address <= _GEN_11072;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_106_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_106_bht <= 2'h1;
        end else begin
          btb_106_bht <= 2'h0;
        end
      end else begin
        btb_106_bht <= _GEN_11074;
      end
    end else begin
      btb_106_bht <= _GEN_11074;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_107_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_107_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_107_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_107_valid <= _GEN_15469;
      end
    end else begin
      btb_107_valid <= _GEN_15469;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_107_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_107_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_107_tag <= _GEN_6251;
      end
    end else begin
      btb_107_tag <= _GEN_6251;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_107_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_107_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_107_target_address <= _GEN_11075;
      end
    end else begin
      btb_107_target_address <= _GEN_11075;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_107_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_107_bht <= 2'h1;
        end else begin
          btb_107_bht <= 2'h0;
        end
      end else begin
        btb_107_bht <= _GEN_11077;
      end
    end else begin
      btb_107_bht <= _GEN_11077;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_108_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_108_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_108_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_108_valid <= _GEN_15470;
      end
    end else begin
      btb_108_valid <= _GEN_15470;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_108_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_108_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_108_tag <= _GEN_6252;
      end
    end else begin
      btb_108_tag <= _GEN_6252;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_108_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_108_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_108_target_address <= _GEN_11078;
      end
    end else begin
      btb_108_target_address <= _GEN_11078;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_108_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_108_bht <= 2'h1;
        end else begin
          btb_108_bht <= 2'h0;
        end
      end else begin
        btb_108_bht <= _GEN_11080;
      end
    end else begin
      btb_108_bht <= _GEN_11080;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_109_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_109_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_109_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_109_valid <= _GEN_15471;
      end
    end else begin
      btb_109_valid <= _GEN_15471;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_109_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_109_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_109_tag <= _GEN_6253;
      end
    end else begin
      btb_109_tag <= _GEN_6253;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_109_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_109_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_109_target_address <= _GEN_11081;
      end
    end else begin
      btb_109_target_address <= _GEN_11081;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_109_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_109_bht <= 2'h1;
        end else begin
          btb_109_bht <= 2'h0;
        end
      end else begin
        btb_109_bht <= _GEN_11083;
      end
    end else begin
      btb_109_bht <= _GEN_11083;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_110_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_110_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_110_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_110_valid <= _GEN_15472;
      end
    end else begin
      btb_110_valid <= _GEN_15472;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_110_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_110_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_110_tag <= _GEN_6254;
      end
    end else begin
      btb_110_tag <= _GEN_6254;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_110_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_110_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_110_target_address <= _GEN_11084;
      end
    end else begin
      btb_110_target_address <= _GEN_11084;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_110_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_110_bht <= 2'h1;
        end else begin
          btb_110_bht <= 2'h0;
        end
      end else begin
        btb_110_bht <= _GEN_11086;
      end
    end else begin
      btb_110_bht <= _GEN_11086;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_111_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_111_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_111_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_111_valid <= _GEN_15473;
      end
    end else begin
      btb_111_valid <= _GEN_15473;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_111_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_111_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_111_tag <= _GEN_6255;
      end
    end else begin
      btb_111_tag <= _GEN_6255;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_111_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_111_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_111_target_address <= _GEN_11087;
      end
    end else begin
      btb_111_target_address <= _GEN_11087;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_111_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h6f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_111_bht <= 2'h1;
        end else begin
          btb_111_bht <= 2'h0;
        end
      end else begin
        btb_111_bht <= _GEN_11089;
      end
    end else begin
      btb_111_bht <= _GEN_11089;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_112_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_112_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_112_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_112_valid <= _GEN_15474;
      end
    end else begin
      btb_112_valid <= _GEN_15474;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_112_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h70 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_112_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_112_tag <= _GEN_6256;
      end
    end else begin
      btb_112_tag <= _GEN_6256;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_112_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h70 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_112_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_112_target_address <= _GEN_11090;
      end
    end else begin
      btb_112_target_address <= _GEN_11090;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_112_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h70 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_112_bht <= 2'h1;
        end else begin
          btb_112_bht <= 2'h0;
        end
      end else begin
        btb_112_bht <= _GEN_11092;
      end
    end else begin
      btb_112_bht <= _GEN_11092;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_113_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_113_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_113_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_113_valid <= _GEN_15475;
      end
    end else begin
      btb_113_valid <= _GEN_15475;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_113_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h71 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_113_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_113_tag <= _GEN_6257;
      end
    end else begin
      btb_113_tag <= _GEN_6257;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_113_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h71 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_113_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_113_target_address <= _GEN_11093;
      end
    end else begin
      btb_113_target_address <= _GEN_11093;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_113_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h71 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_113_bht <= 2'h1;
        end else begin
          btb_113_bht <= 2'h0;
        end
      end else begin
        btb_113_bht <= _GEN_11095;
      end
    end else begin
      btb_113_bht <= _GEN_11095;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_114_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_114_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_114_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_114_valid <= _GEN_15476;
      end
    end else begin
      btb_114_valid <= _GEN_15476;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_114_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h72 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_114_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_114_tag <= _GEN_6258;
      end
    end else begin
      btb_114_tag <= _GEN_6258;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_114_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h72 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_114_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_114_target_address <= _GEN_11096;
      end
    end else begin
      btb_114_target_address <= _GEN_11096;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_114_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h72 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_114_bht <= 2'h1;
        end else begin
          btb_114_bht <= 2'h0;
        end
      end else begin
        btb_114_bht <= _GEN_11098;
      end
    end else begin
      btb_114_bht <= _GEN_11098;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_115_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_115_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_115_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_115_valid <= _GEN_15477;
      end
    end else begin
      btb_115_valid <= _GEN_15477;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_115_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h73 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_115_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_115_tag <= _GEN_6259;
      end
    end else begin
      btb_115_tag <= _GEN_6259;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_115_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h73 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_115_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_115_target_address <= _GEN_11099;
      end
    end else begin
      btb_115_target_address <= _GEN_11099;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_115_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h73 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_115_bht <= 2'h1;
        end else begin
          btb_115_bht <= 2'h0;
        end
      end else begin
        btb_115_bht <= _GEN_11101;
      end
    end else begin
      btb_115_bht <= _GEN_11101;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_116_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_116_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_116_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_116_valid <= _GEN_15478;
      end
    end else begin
      btb_116_valid <= _GEN_15478;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_116_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h74 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_116_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_116_tag <= _GEN_6260;
      end
    end else begin
      btb_116_tag <= _GEN_6260;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_116_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h74 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_116_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_116_target_address <= _GEN_11102;
      end
    end else begin
      btb_116_target_address <= _GEN_11102;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_116_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h74 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_116_bht <= 2'h1;
        end else begin
          btb_116_bht <= 2'h0;
        end
      end else begin
        btb_116_bht <= _GEN_11104;
      end
    end else begin
      btb_116_bht <= _GEN_11104;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_117_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_117_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_117_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_117_valid <= _GEN_15479;
      end
    end else begin
      btb_117_valid <= _GEN_15479;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_117_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h75 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_117_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_117_tag <= _GEN_6261;
      end
    end else begin
      btb_117_tag <= _GEN_6261;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_117_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h75 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_117_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_117_target_address <= _GEN_11105;
      end
    end else begin
      btb_117_target_address <= _GEN_11105;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_117_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h75 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_117_bht <= 2'h1;
        end else begin
          btb_117_bht <= 2'h0;
        end
      end else begin
        btb_117_bht <= _GEN_11107;
      end
    end else begin
      btb_117_bht <= _GEN_11107;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_118_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_118_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_118_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_118_valid <= _GEN_15480;
      end
    end else begin
      btb_118_valid <= _GEN_15480;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_118_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h76 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_118_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_118_tag <= _GEN_6262;
      end
    end else begin
      btb_118_tag <= _GEN_6262;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_118_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h76 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_118_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_118_target_address <= _GEN_11108;
      end
    end else begin
      btb_118_target_address <= _GEN_11108;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_118_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h76 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_118_bht <= 2'h1;
        end else begin
          btb_118_bht <= 2'h0;
        end
      end else begin
        btb_118_bht <= _GEN_11110;
      end
    end else begin
      btb_118_bht <= _GEN_11110;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_119_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_119_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_119_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_119_valid <= _GEN_15481;
      end
    end else begin
      btb_119_valid <= _GEN_15481;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_119_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h77 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_119_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_119_tag <= _GEN_6263;
      end
    end else begin
      btb_119_tag <= _GEN_6263;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_119_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h77 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_119_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_119_target_address <= _GEN_11111;
      end
    end else begin
      btb_119_target_address <= _GEN_11111;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_119_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h77 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_119_bht <= 2'h1;
        end else begin
          btb_119_bht <= 2'h0;
        end
      end else begin
        btb_119_bht <= _GEN_11113;
      end
    end else begin
      btb_119_bht <= _GEN_11113;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_120_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_120_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_120_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_120_valid <= _GEN_15482;
      end
    end else begin
      btb_120_valid <= _GEN_15482;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_120_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h78 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_120_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_120_tag <= _GEN_6264;
      end
    end else begin
      btb_120_tag <= _GEN_6264;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_120_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h78 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_120_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_120_target_address <= _GEN_11114;
      end
    end else begin
      btb_120_target_address <= _GEN_11114;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_120_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h78 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_120_bht <= 2'h1;
        end else begin
          btb_120_bht <= 2'h0;
        end
      end else begin
        btb_120_bht <= _GEN_11116;
      end
    end else begin
      btb_120_bht <= _GEN_11116;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_121_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_121_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_121_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_121_valid <= _GEN_15483;
      end
    end else begin
      btb_121_valid <= _GEN_15483;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_121_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h79 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_121_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_121_tag <= _GEN_6265;
      end
    end else begin
      btb_121_tag <= _GEN_6265;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_121_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h79 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_121_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_121_target_address <= _GEN_11117;
      end
    end else begin
      btb_121_target_address <= _GEN_11117;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_121_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h79 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_121_bht <= 2'h1;
        end else begin
          btb_121_bht <= 2'h0;
        end
      end else begin
        btb_121_bht <= _GEN_11119;
      end
    end else begin
      btb_121_bht <= _GEN_11119;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_122_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_122_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_122_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_122_valid <= _GEN_15484;
      end
    end else begin
      btb_122_valid <= _GEN_15484;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_122_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_122_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_122_tag <= _GEN_6266;
      end
    end else begin
      btb_122_tag <= _GEN_6266;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_122_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_122_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_122_target_address <= _GEN_11120;
      end
    end else begin
      btb_122_target_address <= _GEN_11120;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_122_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_122_bht <= 2'h1;
        end else begin
          btb_122_bht <= 2'h0;
        end
      end else begin
        btb_122_bht <= _GEN_11122;
      end
    end else begin
      btb_122_bht <= _GEN_11122;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_123_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_123_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_123_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_123_valid <= _GEN_15485;
      end
    end else begin
      btb_123_valid <= _GEN_15485;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_123_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_123_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_123_tag <= _GEN_6267;
      end
    end else begin
      btb_123_tag <= _GEN_6267;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_123_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_123_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_123_target_address <= _GEN_11123;
      end
    end else begin
      btb_123_target_address <= _GEN_11123;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_123_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_123_bht <= 2'h1;
        end else begin
          btb_123_bht <= 2'h0;
        end
      end else begin
        btb_123_bht <= _GEN_11125;
      end
    end else begin
      btb_123_bht <= _GEN_11125;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_124_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_124_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_124_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_124_valid <= _GEN_15486;
      end
    end else begin
      btb_124_valid <= _GEN_15486;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_124_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_124_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_124_tag <= _GEN_6268;
      end
    end else begin
      btb_124_tag <= _GEN_6268;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_124_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_124_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_124_target_address <= _GEN_11126;
      end
    end else begin
      btb_124_target_address <= _GEN_11126;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_124_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_124_bht <= 2'h1;
        end else begin
          btb_124_bht <= 2'h0;
        end
      end else begin
        btb_124_bht <= _GEN_11128;
      end
    end else begin
      btb_124_bht <= _GEN_11128;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_125_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_125_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_125_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_125_valid <= _GEN_15487;
      end
    end else begin
      btb_125_valid <= _GEN_15487;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_125_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_125_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_125_tag <= _GEN_6269;
      end
    end else begin
      btb_125_tag <= _GEN_6269;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_125_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_125_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_125_target_address <= _GEN_11129;
      end
    end else begin
      btb_125_target_address <= _GEN_11129;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_125_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_125_bht <= 2'h1;
        end else begin
          btb_125_bht <= 2'h0;
        end
      end else begin
        btb_125_bht <= _GEN_11131;
      end
    end else begin
      btb_125_bht <= _GEN_11131;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_126_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_126_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_126_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_126_valid <= _GEN_15488;
      end
    end else begin
      btb_126_valid <= _GEN_15488;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_126_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_126_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_126_tag <= _GEN_6270;
      end
    end else begin
      btb_126_tag <= _GEN_6270;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_126_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_126_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_126_target_address <= _GEN_11132;
      end
    end else begin
      btb_126_target_address <= _GEN_11132;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_126_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_126_bht <= 2'h1;
        end else begin
          btb_126_bht <= 2'h0;
        end
      end else begin
        btb_126_bht <= _GEN_11134;
      end
    end else begin
      btb_126_bht <= _GEN_11134;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_127_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_127_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_127_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_127_valid <= _GEN_15489;
      end
    end else begin
      btb_127_valid <= _GEN_15489;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_127_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_127_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_127_tag <= _GEN_6271;
      end
    end else begin
      btb_127_tag <= _GEN_6271;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_127_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_127_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_127_target_address <= _GEN_11135;
      end
    end else begin
      btb_127_target_address <= _GEN_11135;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_127_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h7f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_127_bht <= 2'h1;
        end else begin
          btb_127_bht <= 2'h0;
        end
      end else begin
        btb_127_bht <= _GEN_11137;
      end
    end else begin
      btb_127_bht <= _GEN_11137;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_128_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_128_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_128_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_128_valid <= _GEN_15490;
      end
    end else begin
      btb_128_valid <= _GEN_15490;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_128_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h80 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_128_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_128_tag <= _GEN_6272;
      end
    end else begin
      btb_128_tag <= _GEN_6272;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_128_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h80 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_128_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_128_target_address <= _GEN_11138;
      end
    end else begin
      btb_128_target_address <= _GEN_11138;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_128_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h80 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_128_bht <= 2'h1;
        end else begin
          btb_128_bht <= 2'h0;
        end
      end else begin
        btb_128_bht <= _GEN_11140;
      end
    end else begin
      btb_128_bht <= _GEN_11140;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_129_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_129_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_129_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_129_valid <= _GEN_15491;
      end
    end else begin
      btb_129_valid <= _GEN_15491;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_129_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h81 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_129_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_129_tag <= _GEN_6273;
      end
    end else begin
      btb_129_tag <= _GEN_6273;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_129_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h81 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_129_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_129_target_address <= _GEN_11141;
      end
    end else begin
      btb_129_target_address <= _GEN_11141;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_129_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h81 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_129_bht <= 2'h1;
        end else begin
          btb_129_bht <= 2'h0;
        end
      end else begin
        btb_129_bht <= _GEN_11143;
      end
    end else begin
      btb_129_bht <= _GEN_11143;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_130_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_130_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_130_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_130_valid <= _GEN_15492;
      end
    end else begin
      btb_130_valid <= _GEN_15492;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_130_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h82 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_130_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_130_tag <= _GEN_6274;
      end
    end else begin
      btb_130_tag <= _GEN_6274;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_130_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h82 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_130_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_130_target_address <= _GEN_11144;
      end
    end else begin
      btb_130_target_address <= _GEN_11144;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_130_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h82 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_130_bht <= 2'h1;
        end else begin
          btb_130_bht <= 2'h0;
        end
      end else begin
        btb_130_bht <= _GEN_11146;
      end
    end else begin
      btb_130_bht <= _GEN_11146;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_131_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_131_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_131_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_131_valid <= _GEN_15493;
      end
    end else begin
      btb_131_valid <= _GEN_15493;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_131_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h83 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_131_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_131_tag <= _GEN_6275;
      end
    end else begin
      btb_131_tag <= _GEN_6275;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_131_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h83 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_131_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_131_target_address <= _GEN_11147;
      end
    end else begin
      btb_131_target_address <= _GEN_11147;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_131_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h83 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_131_bht <= 2'h1;
        end else begin
          btb_131_bht <= 2'h0;
        end
      end else begin
        btb_131_bht <= _GEN_11149;
      end
    end else begin
      btb_131_bht <= _GEN_11149;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_132_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_132_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_132_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_132_valid <= _GEN_15494;
      end
    end else begin
      btb_132_valid <= _GEN_15494;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_132_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h84 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_132_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_132_tag <= _GEN_6276;
      end
    end else begin
      btb_132_tag <= _GEN_6276;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_132_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h84 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_132_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_132_target_address <= _GEN_11150;
      end
    end else begin
      btb_132_target_address <= _GEN_11150;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_132_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h84 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_132_bht <= 2'h1;
        end else begin
          btb_132_bht <= 2'h0;
        end
      end else begin
        btb_132_bht <= _GEN_11152;
      end
    end else begin
      btb_132_bht <= _GEN_11152;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_133_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_133_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_133_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_133_valid <= _GEN_15495;
      end
    end else begin
      btb_133_valid <= _GEN_15495;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_133_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h85 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_133_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_133_tag <= _GEN_6277;
      end
    end else begin
      btb_133_tag <= _GEN_6277;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_133_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h85 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_133_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_133_target_address <= _GEN_11153;
      end
    end else begin
      btb_133_target_address <= _GEN_11153;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_133_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h85 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_133_bht <= 2'h1;
        end else begin
          btb_133_bht <= 2'h0;
        end
      end else begin
        btb_133_bht <= _GEN_11155;
      end
    end else begin
      btb_133_bht <= _GEN_11155;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_134_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_134_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_134_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_134_valid <= _GEN_15496;
      end
    end else begin
      btb_134_valid <= _GEN_15496;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_134_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h86 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_134_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_134_tag <= _GEN_6278;
      end
    end else begin
      btb_134_tag <= _GEN_6278;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_134_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h86 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_134_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_134_target_address <= _GEN_11156;
      end
    end else begin
      btb_134_target_address <= _GEN_11156;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_134_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h86 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_134_bht <= 2'h1;
        end else begin
          btb_134_bht <= 2'h0;
        end
      end else begin
        btb_134_bht <= _GEN_11158;
      end
    end else begin
      btb_134_bht <= _GEN_11158;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_135_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_135_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_135_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_135_valid <= _GEN_15497;
      end
    end else begin
      btb_135_valid <= _GEN_15497;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_135_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h87 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_135_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_135_tag <= _GEN_6279;
      end
    end else begin
      btb_135_tag <= _GEN_6279;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_135_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h87 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_135_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_135_target_address <= _GEN_11159;
      end
    end else begin
      btb_135_target_address <= _GEN_11159;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_135_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h87 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_135_bht <= 2'h1;
        end else begin
          btb_135_bht <= 2'h0;
        end
      end else begin
        btb_135_bht <= _GEN_11161;
      end
    end else begin
      btb_135_bht <= _GEN_11161;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_136_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_136_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_136_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_136_valid <= _GEN_15498;
      end
    end else begin
      btb_136_valid <= _GEN_15498;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_136_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h88 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_136_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_136_tag <= _GEN_6280;
      end
    end else begin
      btb_136_tag <= _GEN_6280;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_136_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h88 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_136_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_136_target_address <= _GEN_11162;
      end
    end else begin
      btb_136_target_address <= _GEN_11162;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_136_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h88 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_136_bht <= 2'h1;
        end else begin
          btb_136_bht <= 2'h0;
        end
      end else begin
        btb_136_bht <= _GEN_11164;
      end
    end else begin
      btb_136_bht <= _GEN_11164;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_137_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_137_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_137_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_137_valid <= _GEN_15499;
      end
    end else begin
      btb_137_valid <= _GEN_15499;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_137_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h89 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_137_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_137_tag <= _GEN_6281;
      end
    end else begin
      btb_137_tag <= _GEN_6281;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_137_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h89 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_137_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_137_target_address <= _GEN_11165;
      end
    end else begin
      btb_137_target_address <= _GEN_11165;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_137_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h89 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_137_bht <= 2'h1;
        end else begin
          btb_137_bht <= 2'h0;
        end
      end else begin
        btb_137_bht <= _GEN_11167;
      end
    end else begin
      btb_137_bht <= _GEN_11167;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_138_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_138_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_138_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_138_valid <= _GEN_15500;
      end
    end else begin
      btb_138_valid <= _GEN_15500;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_138_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_138_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_138_tag <= _GEN_6282;
      end
    end else begin
      btb_138_tag <= _GEN_6282;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_138_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_138_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_138_target_address <= _GEN_11168;
      end
    end else begin
      btb_138_target_address <= _GEN_11168;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_138_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_138_bht <= 2'h1;
        end else begin
          btb_138_bht <= 2'h0;
        end
      end else begin
        btb_138_bht <= _GEN_11170;
      end
    end else begin
      btb_138_bht <= _GEN_11170;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_139_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_139_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_139_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_139_valid <= _GEN_15501;
      end
    end else begin
      btb_139_valid <= _GEN_15501;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_139_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_139_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_139_tag <= _GEN_6283;
      end
    end else begin
      btb_139_tag <= _GEN_6283;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_139_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_139_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_139_target_address <= _GEN_11171;
      end
    end else begin
      btb_139_target_address <= _GEN_11171;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_139_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_139_bht <= 2'h1;
        end else begin
          btb_139_bht <= 2'h0;
        end
      end else begin
        btb_139_bht <= _GEN_11173;
      end
    end else begin
      btb_139_bht <= _GEN_11173;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_140_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_140_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_140_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_140_valid <= _GEN_15502;
      end
    end else begin
      btb_140_valid <= _GEN_15502;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_140_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_140_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_140_tag <= _GEN_6284;
      end
    end else begin
      btb_140_tag <= _GEN_6284;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_140_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_140_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_140_target_address <= _GEN_11174;
      end
    end else begin
      btb_140_target_address <= _GEN_11174;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_140_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_140_bht <= 2'h1;
        end else begin
          btb_140_bht <= 2'h0;
        end
      end else begin
        btb_140_bht <= _GEN_11176;
      end
    end else begin
      btb_140_bht <= _GEN_11176;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_141_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_141_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_141_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_141_valid <= _GEN_15503;
      end
    end else begin
      btb_141_valid <= _GEN_15503;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_141_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_141_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_141_tag <= _GEN_6285;
      end
    end else begin
      btb_141_tag <= _GEN_6285;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_141_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_141_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_141_target_address <= _GEN_11177;
      end
    end else begin
      btb_141_target_address <= _GEN_11177;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_141_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_141_bht <= 2'h1;
        end else begin
          btb_141_bht <= 2'h0;
        end
      end else begin
        btb_141_bht <= _GEN_11179;
      end
    end else begin
      btb_141_bht <= _GEN_11179;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_142_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_142_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_142_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_142_valid <= _GEN_15504;
      end
    end else begin
      btb_142_valid <= _GEN_15504;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_142_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_142_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_142_tag <= _GEN_6286;
      end
    end else begin
      btb_142_tag <= _GEN_6286;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_142_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_142_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_142_target_address <= _GEN_11180;
      end
    end else begin
      btb_142_target_address <= _GEN_11180;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_142_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_142_bht <= 2'h1;
        end else begin
          btb_142_bht <= 2'h0;
        end
      end else begin
        btb_142_bht <= _GEN_11182;
      end
    end else begin
      btb_142_bht <= _GEN_11182;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_143_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_143_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_143_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_143_valid <= _GEN_15505;
      end
    end else begin
      btb_143_valid <= _GEN_15505;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_143_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_143_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_143_tag <= _GEN_6287;
      end
    end else begin
      btb_143_tag <= _GEN_6287;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_143_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_143_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_143_target_address <= _GEN_11183;
      end
    end else begin
      btb_143_target_address <= _GEN_11183;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_143_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h8f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_143_bht <= 2'h1;
        end else begin
          btb_143_bht <= 2'h0;
        end
      end else begin
        btb_143_bht <= _GEN_11185;
      end
    end else begin
      btb_143_bht <= _GEN_11185;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_144_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_144_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_144_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_144_valid <= _GEN_15506;
      end
    end else begin
      btb_144_valid <= _GEN_15506;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_144_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h90 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_144_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_144_tag <= _GEN_6288;
      end
    end else begin
      btb_144_tag <= _GEN_6288;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_144_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h90 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_144_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_144_target_address <= _GEN_11186;
      end
    end else begin
      btb_144_target_address <= _GEN_11186;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_144_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h90 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_144_bht <= 2'h1;
        end else begin
          btb_144_bht <= 2'h0;
        end
      end else begin
        btb_144_bht <= _GEN_11188;
      end
    end else begin
      btb_144_bht <= _GEN_11188;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_145_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_145_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_145_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_145_valid <= _GEN_15507;
      end
    end else begin
      btb_145_valid <= _GEN_15507;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_145_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h91 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_145_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_145_tag <= _GEN_6289;
      end
    end else begin
      btb_145_tag <= _GEN_6289;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_145_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h91 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_145_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_145_target_address <= _GEN_11189;
      end
    end else begin
      btb_145_target_address <= _GEN_11189;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_145_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h91 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_145_bht <= 2'h1;
        end else begin
          btb_145_bht <= 2'h0;
        end
      end else begin
        btb_145_bht <= _GEN_11191;
      end
    end else begin
      btb_145_bht <= _GEN_11191;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_146_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_146_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_146_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_146_valid <= _GEN_15508;
      end
    end else begin
      btb_146_valid <= _GEN_15508;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_146_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h92 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_146_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_146_tag <= _GEN_6290;
      end
    end else begin
      btb_146_tag <= _GEN_6290;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_146_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h92 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_146_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_146_target_address <= _GEN_11192;
      end
    end else begin
      btb_146_target_address <= _GEN_11192;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_146_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h92 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_146_bht <= 2'h1;
        end else begin
          btb_146_bht <= 2'h0;
        end
      end else begin
        btb_146_bht <= _GEN_11194;
      end
    end else begin
      btb_146_bht <= _GEN_11194;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_147_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_147_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_147_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_147_valid <= _GEN_15509;
      end
    end else begin
      btb_147_valid <= _GEN_15509;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_147_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h93 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_147_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_147_tag <= _GEN_6291;
      end
    end else begin
      btb_147_tag <= _GEN_6291;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_147_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h93 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_147_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_147_target_address <= _GEN_11195;
      end
    end else begin
      btb_147_target_address <= _GEN_11195;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_147_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h93 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_147_bht <= 2'h1;
        end else begin
          btb_147_bht <= 2'h0;
        end
      end else begin
        btb_147_bht <= _GEN_11197;
      end
    end else begin
      btb_147_bht <= _GEN_11197;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_148_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_148_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_148_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_148_valid <= _GEN_15510;
      end
    end else begin
      btb_148_valid <= _GEN_15510;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_148_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h94 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_148_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_148_tag <= _GEN_6292;
      end
    end else begin
      btb_148_tag <= _GEN_6292;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_148_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h94 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_148_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_148_target_address <= _GEN_11198;
      end
    end else begin
      btb_148_target_address <= _GEN_11198;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_148_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h94 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_148_bht <= 2'h1;
        end else begin
          btb_148_bht <= 2'h0;
        end
      end else begin
        btb_148_bht <= _GEN_11200;
      end
    end else begin
      btb_148_bht <= _GEN_11200;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_149_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_149_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_149_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_149_valid <= _GEN_15511;
      end
    end else begin
      btb_149_valid <= _GEN_15511;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_149_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h95 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_149_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_149_tag <= _GEN_6293;
      end
    end else begin
      btb_149_tag <= _GEN_6293;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_149_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h95 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_149_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_149_target_address <= _GEN_11201;
      end
    end else begin
      btb_149_target_address <= _GEN_11201;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_149_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h95 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_149_bht <= 2'h1;
        end else begin
          btb_149_bht <= 2'h0;
        end
      end else begin
        btb_149_bht <= _GEN_11203;
      end
    end else begin
      btb_149_bht <= _GEN_11203;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_150_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_150_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_150_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_150_valid <= _GEN_15512;
      end
    end else begin
      btb_150_valid <= _GEN_15512;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_150_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h96 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_150_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_150_tag <= _GEN_6294;
      end
    end else begin
      btb_150_tag <= _GEN_6294;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_150_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h96 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_150_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_150_target_address <= _GEN_11204;
      end
    end else begin
      btb_150_target_address <= _GEN_11204;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_150_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h96 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_150_bht <= 2'h1;
        end else begin
          btb_150_bht <= 2'h0;
        end
      end else begin
        btb_150_bht <= _GEN_11206;
      end
    end else begin
      btb_150_bht <= _GEN_11206;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_151_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_151_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_151_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_151_valid <= _GEN_15513;
      end
    end else begin
      btb_151_valid <= _GEN_15513;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_151_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h97 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_151_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_151_tag <= _GEN_6295;
      end
    end else begin
      btb_151_tag <= _GEN_6295;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_151_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h97 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_151_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_151_target_address <= _GEN_11207;
      end
    end else begin
      btb_151_target_address <= _GEN_11207;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_151_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h97 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_151_bht <= 2'h1;
        end else begin
          btb_151_bht <= 2'h0;
        end
      end else begin
        btb_151_bht <= _GEN_11209;
      end
    end else begin
      btb_151_bht <= _GEN_11209;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_152_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_152_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_152_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_152_valid <= _GEN_15514;
      end
    end else begin
      btb_152_valid <= _GEN_15514;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_152_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h98 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_152_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_152_tag <= _GEN_6296;
      end
    end else begin
      btb_152_tag <= _GEN_6296;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_152_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h98 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_152_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_152_target_address <= _GEN_11210;
      end
    end else begin
      btb_152_target_address <= _GEN_11210;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_152_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h98 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_152_bht <= 2'h1;
        end else begin
          btb_152_bht <= 2'h0;
        end
      end else begin
        btb_152_bht <= _GEN_11212;
      end
    end else begin
      btb_152_bht <= _GEN_11212;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_153_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_153_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_153_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_153_valid <= _GEN_15515;
      end
    end else begin
      btb_153_valid <= _GEN_15515;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_153_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h99 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_153_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_153_tag <= _GEN_6297;
      end
    end else begin
      btb_153_tag <= _GEN_6297;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_153_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h99 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_153_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_153_target_address <= _GEN_11213;
      end
    end else begin
      btb_153_target_address <= _GEN_11213;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_153_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h99 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_153_bht <= 2'h1;
        end else begin
          btb_153_bht <= 2'h0;
        end
      end else begin
        btb_153_bht <= _GEN_11215;
      end
    end else begin
      btb_153_bht <= _GEN_11215;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_154_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_154_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_154_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_154_valid <= _GEN_15516;
      end
    end else begin
      btb_154_valid <= _GEN_15516;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_154_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_154_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_154_tag <= _GEN_6298;
      end
    end else begin
      btb_154_tag <= _GEN_6298;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_154_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_154_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_154_target_address <= _GEN_11216;
      end
    end else begin
      btb_154_target_address <= _GEN_11216;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_154_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_154_bht <= 2'h1;
        end else begin
          btb_154_bht <= 2'h0;
        end
      end else begin
        btb_154_bht <= _GEN_11218;
      end
    end else begin
      btb_154_bht <= _GEN_11218;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_155_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_155_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_155_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_155_valid <= _GEN_15517;
      end
    end else begin
      btb_155_valid <= _GEN_15517;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_155_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_155_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_155_tag <= _GEN_6299;
      end
    end else begin
      btb_155_tag <= _GEN_6299;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_155_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_155_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_155_target_address <= _GEN_11219;
      end
    end else begin
      btb_155_target_address <= _GEN_11219;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_155_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_155_bht <= 2'h1;
        end else begin
          btb_155_bht <= 2'h0;
        end
      end else begin
        btb_155_bht <= _GEN_11221;
      end
    end else begin
      btb_155_bht <= _GEN_11221;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_156_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_156_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_156_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_156_valid <= _GEN_15518;
      end
    end else begin
      btb_156_valid <= _GEN_15518;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_156_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_156_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_156_tag <= _GEN_6300;
      end
    end else begin
      btb_156_tag <= _GEN_6300;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_156_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_156_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_156_target_address <= _GEN_11222;
      end
    end else begin
      btb_156_target_address <= _GEN_11222;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_156_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_156_bht <= 2'h1;
        end else begin
          btb_156_bht <= 2'h0;
        end
      end else begin
        btb_156_bht <= _GEN_11224;
      end
    end else begin
      btb_156_bht <= _GEN_11224;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_157_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_157_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_157_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_157_valid <= _GEN_15519;
      end
    end else begin
      btb_157_valid <= _GEN_15519;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_157_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_157_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_157_tag <= _GEN_6301;
      end
    end else begin
      btb_157_tag <= _GEN_6301;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_157_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_157_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_157_target_address <= _GEN_11225;
      end
    end else begin
      btb_157_target_address <= _GEN_11225;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_157_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_157_bht <= 2'h1;
        end else begin
          btb_157_bht <= 2'h0;
        end
      end else begin
        btb_157_bht <= _GEN_11227;
      end
    end else begin
      btb_157_bht <= _GEN_11227;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_158_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_158_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_158_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_158_valid <= _GEN_15520;
      end
    end else begin
      btb_158_valid <= _GEN_15520;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_158_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_158_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_158_tag <= _GEN_6302;
      end
    end else begin
      btb_158_tag <= _GEN_6302;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_158_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_158_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_158_target_address <= _GEN_11228;
      end
    end else begin
      btb_158_target_address <= _GEN_11228;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_158_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_158_bht <= 2'h1;
        end else begin
          btb_158_bht <= 2'h0;
        end
      end else begin
        btb_158_bht <= _GEN_11230;
      end
    end else begin
      btb_158_bht <= _GEN_11230;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_159_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_159_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_159_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_159_valid <= _GEN_15521;
      end
    end else begin
      btb_159_valid <= _GEN_15521;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_159_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_159_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_159_tag <= _GEN_6303;
      end
    end else begin
      btb_159_tag <= _GEN_6303;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_159_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_159_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_159_target_address <= _GEN_11231;
      end
    end else begin
      btb_159_target_address <= _GEN_11231;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_159_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h9f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_159_bht <= 2'h1;
        end else begin
          btb_159_bht <= 2'h0;
        end
      end else begin
        btb_159_bht <= _GEN_11233;
      end
    end else begin
      btb_159_bht <= _GEN_11233;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_160_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_160_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_160_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_160_valid <= _GEN_15522;
      end
    end else begin
      btb_160_valid <= _GEN_15522;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_160_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_160_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_160_tag <= _GEN_6304;
      end
    end else begin
      btb_160_tag <= _GEN_6304;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_160_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_160_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_160_target_address <= _GEN_11234;
      end
    end else begin
      btb_160_target_address <= _GEN_11234;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_160_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_160_bht <= 2'h1;
        end else begin
          btb_160_bht <= 2'h0;
        end
      end else begin
        btb_160_bht <= _GEN_11236;
      end
    end else begin
      btb_160_bht <= _GEN_11236;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_161_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_161_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_161_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_161_valid <= _GEN_15523;
      end
    end else begin
      btb_161_valid <= _GEN_15523;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_161_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_161_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_161_tag <= _GEN_6305;
      end
    end else begin
      btb_161_tag <= _GEN_6305;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_161_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_161_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_161_target_address <= _GEN_11237;
      end
    end else begin
      btb_161_target_address <= _GEN_11237;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_161_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_161_bht <= 2'h1;
        end else begin
          btb_161_bht <= 2'h0;
        end
      end else begin
        btb_161_bht <= _GEN_11239;
      end
    end else begin
      btb_161_bht <= _GEN_11239;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_162_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_162_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_162_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_162_valid <= _GEN_15524;
      end
    end else begin
      btb_162_valid <= _GEN_15524;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_162_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_162_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_162_tag <= _GEN_6306;
      end
    end else begin
      btb_162_tag <= _GEN_6306;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_162_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_162_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_162_target_address <= _GEN_11240;
      end
    end else begin
      btb_162_target_address <= _GEN_11240;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_162_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_162_bht <= 2'h1;
        end else begin
          btb_162_bht <= 2'h0;
        end
      end else begin
        btb_162_bht <= _GEN_11242;
      end
    end else begin
      btb_162_bht <= _GEN_11242;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_163_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_163_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_163_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_163_valid <= _GEN_15525;
      end
    end else begin
      btb_163_valid <= _GEN_15525;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_163_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_163_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_163_tag <= _GEN_6307;
      end
    end else begin
      btb_163_tag <= _GEN_6307;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_163_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_163_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_163_target_address <= _GEN_11243;
      end
    end else begin
      btb_163_target_address <= _GEN_11243;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_163_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_163_bht <= 2'h1;
        end else begin
          btb_163_bht <= 2'h0;
        end
      end else begin
        btb_163_bht <= _GEN_11245;
      end
    end else begin
      btb_163_bht <= _GEN_11245;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_164_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_164_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_164_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_164_valid <= _GEN_15526;
      end
    end else begin
      btb_164_valid <= _GEN_15526;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_164_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_164_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_164_tag <= _GEN_6308;
      end
    end else begin
      btb_164_tag <= _GEN_6308;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_164_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_164_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_164_target_address <= _GEN_11246;
      end
    end else begin
      btb_164_target_address <= _GEN_11246;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_164_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_164_bht <= 2'h1;
        end else begin
          btb_164_bht <= 2'h0;
        end
      end else begin
        btb_164_bht <= _GEN_11248;
      end
    end else begin
      btb_164_bht <= _GEN_11248;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_165_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_165_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_165_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_165_valid <= _GEN_15527;
      end
    end else begin
      btb_165_valid <= _GEN_15527;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_165_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_165_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_165_tag <= _GEN_6309;
      end
    end else begin
      btb_165_tag <= _GEN_6309;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_165_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_165_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_165_target_address <= _GEN_11249;
      end
    end else begin
      btb_165_target_address <= _GEN_11249;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_165_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_165_bht <= 2'h1;
        end else begin
          btb_165_bht <= 2'h0;
        end
      end else begin
        btb_165_bht <= _GEN_11251;
      end
    end else begin
      btb_165_bht <= _GEN_11251;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_166_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_166_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_166_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_166_valid <= _GEN_15528;
      end
    end else begin
      btb_166_valid <= _GEN_15528;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_166_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_166_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_166_tag <= _GEN_6310;
      end
    end else begin
      btb_166_tag <= _GEN_6310;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_166_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_166_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_166_target_address <= _GEN_11252;
      end
    end else begin
      btb_166_target_address <= _GEN_11252;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_166_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_166_bht <= 2'h1;
        end else begin
          btb_166_bht <= 2'h0;
        end
      end else begin
        btb_166_bht <= _GEN_11254;
      end
    end else begin
      btb_166_bht <= _GEN_11254;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_167_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_167_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_167_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_167_valid <= _GEN_15529;
      end
    end else begin
      btb_167_valid <= _GEN_15529;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_167_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_167_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_167_tag <= _GEN_6311;
      end
    end else begin
      btb_167_tag <= _GEN_6311;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_167_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_167_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_167_target_address <= _GEN_11255;
      end
    end else begin
      btb_167_target_address <= _GEN_11255;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_167_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_167_bht <= 2'h1;
        end else begin
          btb_167_bht <= 2'h0;
        end
      end else begin
        btb_167_bht <= _GEN_11257;
      end
    end else begin
      btb_167_bht <= _GEN_11257;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_168_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_168_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_168_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_168_valid <= _GEN_15530;
      end
    end else begin
      btb_168_valid <= _GEN_15530;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_168_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_168_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_168_tag <= _GEN_6312;
      end
    end else begin
      btb_168_tag <= _GEN_6312;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_168_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_168_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_168_target_address <= _GEN_11258;
      end
    end else begin
      btb_168_target_address <= _GEN_11258;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_168_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_168_bht <= 2'h1;
        end else begin
          btb_168_bht <= 2'h0;
        end
      end else begin
        btb_168_bht <= _GEN_11260;
      end
    end else begin
      btb_168_bht <= _GEN_11260;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_169_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_169_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_169_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_169_valid <= _GEN_15531;
      end
    end else begin
      btb_169_valid <= _GEN_15531;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_169_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_169_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_169_tag <= _GEN_6313;
      end
    end else begin
      btb_169_tag <= _GEN_6313;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_169_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_169_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_169_target_address <= _GEN_11261;
      end
    end else begin
      btb_169_target_address <= _GEN_11261;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_169_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'ha9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_169_bht <= 2'h1;
        end else begin
          btb_169_bht <= 2'h0;
        end
      end else begin
        btb_169_bht <= _GEN_11263;
      end
    end else begin
      btb_169_bht <= _GEN_11263;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_170_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_170_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_170_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_170_valid <= _GEN_15532;
      end
    end else begin
      btb_170_valid <= _GEN_15532;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_170_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'haa == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_170_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_170_tag <= _GEN_6314;
      end
    end else begin
      btb_170_tag <= _GEN_6314;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_170_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'haa == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_170_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_170_target_address <= _GEN_11264;
      end
    end else begin
      btb_170_target_address <= _GEN_11264;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_170_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'haa == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_170_bht <= 2'h1;
        end else begin
          btb_170_bht <= 2'h0;
        end
      end else begin
        btb_170_bht <= _GEN_11266;
      end
    end else begin
      btb_170_bht <= _GEN_11266;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_171_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_171_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_171_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_171_valid <= _GEN_15533;
      end
    end else begin
      btb_171_valid <= _GEN_15533;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_171_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hab == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_171_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_171_tag <= _GEN_6315;
      end
    end else begin
      btb_171_tag <= _GEN_6315;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_171_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hab == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_171_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_171_target_address <= _GEN_11267;
      end
    end else begin
      btb_171_target_address <= _GEN_11267;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_171_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hab == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_171_bht <= 2'h1;
        end else begin
          btb_171_bht <= 2'h0;
        end
      end else begin
        btb_171_bht <= _GEN_11269;
      end
    end else begin
      btb_171_bht <= _GEN_11269;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_172_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_172_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_172_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_172_valid <= _GEN_15534;
      end
    end else begin
      btb_172_valid <= _GEN_15534;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_172_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hac == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_172_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_172_tag <= _GEN_6316;
      end
    end else begin
      btb_172_tag <= _GEN_6316;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_172_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hac == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_172_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_172_target_address <= _GEN_11270;
      end
    end else begin
      btb_172_target_address <= _GEN_11270;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_172_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hac == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_172_bht <= 2'h1;
        end else begin
          btb_172_bht <= 2'h0;
        end
      end else begin
        btb_172_bht <= _GEN_11272;
      end
    end else begin
      btb_172_bht <= _GEN_11272;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_173_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_173_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_173_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_173_valid <= _GEN_15535;
      end
    end else begin
      btb_173_valid <= _GEN_15535;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_173_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'had == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_173_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_173_tag <= _GEN_6317;
      end
    end else begin
      btb_173_tag <= _GEN_6317;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_173_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'had == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_173_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_173_target_address <= _GEN_11273;
      end
    end else begin
      btb_173_target_address <= _GEN_11273;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_173_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'had == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_173_bht <= 2'h1;
        end else begin
          btb_173_bht <= 2'h0;
        end
      end else begin
        btb_173_bht <= _GEN_11275;
      end
    end else begin
      btb_173_bht <= _GEN_11275;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_174_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_174_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_174_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_174_valid <= _GEN_15536;
      end
    end else begin
      btb_174_valid <= _GEN_15536;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_174_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hae == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_174_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_174_tag <= _GEN_6318;
      end
    end else begin
      btb_174_tag <= _GEN_6318;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_174_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hae == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_174_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_174_target_address <= _GEN_11276;
      end
    end else begin
      btb_174_target_address <= _GEN_11276;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_174_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hae == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_174_bht <= 2'h1;
        end else begin
          btb_174_bht <= 2'h0;
        end
      end else begin
        btb_174_bht <= _GEN_11278;
      end
    end else begin
      btb_174_bht <= _GEN_11278;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_175_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_175_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_175_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_175_valid <= _GEN_15537;
      end
    end else begin
      btb_175_valid <= _GEN_15537;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_175_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'haf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_175_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_175_tag <= _GEN_6319;
      end
    end else begin
      btb_175_tag <= _GEN_6319;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_175_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'haf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_175_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_175_target_address <= _GEN_11279;
      end
    end else begin
      btb_175_target_address <= _GEN_11279;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_175_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'haf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_175_bht <= 2'h1;
        end else begin
          btb_175_bht <= 2'h0;
        end
      end else begin
        btb_175_bht <= _GEN_11281;
      end
    end else begin
      btb_175_bht <= _GEN_11281;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_176_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_176_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_176_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_176_valid <= _GEN_15538;
      end
    end else begin
      btb_176_valid <= _GEN_15538;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_176_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_176_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_176_tag <= _GEN_6320;
      end
    end else begin
      btb_176_tag <= _GEN_6320;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_176_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_176_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_176_target_address <= _GEN_11282;
      end
    end else begin
      btb_176_target_address <= _GEN_11282;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_176_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_176_bht <= 2'h1;
        end else begin
          btb_176_bht <= 2'h0;
        end
      end else begin
        btb_176_bht <= _GEN_11284;
      end
    end else begin
      btb_176_bht <= _GEN_11284;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_177_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_177_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_177_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_177_valid <= _GEN_15539;
      end
    end else begin
      btb_177_valid <= _GEN_15539;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_177_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_177_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_177_tag <= _GEN_6321;
      end
    end else begin
      btb_177_tag <= _GEN_6321;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_177_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_177_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_177_target_address <= _GEN_11285;
      end
    end else begin
      btb_177_target_address <= _GEN_11285;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_177_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_177_bht <= 2'h1;
        end else begin
          btb_177_bht <= 2'h0;
        end
      end else begin
        btb_177_bht <= _GEN_11287;
      end
    end else begin
      btb_177_bht <= _GEN_11287;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_178_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_178_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_178_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_178_valid <= _GEN_15540;
      end
    end else begin
      btb_178_valid <= _GEN_15540;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_178_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_178_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_178_tag <= _GEN_6322;
      end
    end else begin
      btb_178_tag <= _GEN_6322;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_178_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_178_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_178_target_address <= _GEN_11288;
      end
    end else begin
      btb_178_target_address <= _GEN_11288;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_178_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_178_bht <= 2'h1;
        end else begin
          btb_178_bht <= 2'h0;
        end
      end else begin
        btb_178_bht <= _GEN_11290;
      end
    end else begin
      btb_178_bht <= _GEN_11290;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_179_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_179_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_179_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_179_valid <= _GEN_15541;
      end
    end else begin
      btb_179_valid <= _GEN_15541;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_179_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_179_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_179_tag <= _GEN_6323;
      end
    end else begin
      btb_179_tag <= _GEN_6323;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_179_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_179_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_179_target_address <= _GEN_11291;
      end
    end else begin
      btb_179_target_address <= _GEN_11291;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_179_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_179_bht <= 2'h1;
        end else begin
          btb_179_bht <= 2'h0;
        end
      end else begin
        btb_179_bht <= _GEN_11293;
      end
    end else begin
      btb_179_bht <= _GEN_11293;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_180_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_180_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_180_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_180_valid <= _GEN_15542;
      end
    end else begin
      btb_180_valid <= _GEN_15542;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_180_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_180_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_180_tag <= _GEN_6324;
      end
    end else begin
      btb_180_tag <= _GEN_6324;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_180_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_180_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_180_target_address <= _GEN_11294;
      end
    end else begin
      btb_180_target_address <= _GEN_11294;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_180_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_180_bht <= 2'h1;
        end else begin
          btb_180_bht <= 2'h0;
        end
      end else begin
        btb_180_bht <= _GEN_11296;
      end
    end else begin
      btb_180_bht <= _GEN_11296;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_181_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_181_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_181_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_181_valid <= _GEN_15543;
      end
    end else begin
      btb_181_valid <= _GEN_15543;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_181_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_181_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_181_tag <= _GEN_6325;
      end
    end else begin
      btb_181_tag <= _GEN_6325;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_181_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_181_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_181_target_address <= _GEN_11297;
      end
    end else begin
      btb_181_target_address <= _GEN_11297;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_181_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_181_bht <= 2'h1;
        end else begin
          btb_181_bht <= 2'h0;
        end
      end else begin
        btb_181_bht <= _GEN_11299;
      end
    end else begin
      btb_181_bht <= _GEN_11299;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_182_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_182_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_182_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_182_valid <= _GEN_15544;
      end
    end else begin
      btb_182_valid <= _GEN_15544;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_182_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_182_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_182_tag <= _GEN_6326;
      end
    end else begin
      btb_182_tag <= _GEN_6326;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_182_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_182_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_182_target_address <= _GEN_11300;
      end
    end else begin
      btb_182_target_address <= _GEN_11300;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_182_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_182_bht <= 2'h1;
        end else begin
          btb_182_bht <= 2'h0;
        end
      end else begin
        btb_182_bht <= _GEN_11302;
      end
    end else begin
      btb_182_bht <= _GEN_11302;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_183_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_183_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_183_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_183_valid <= _GEN_15545;
      end
    end else begin
      btb_183_valid <= _GEN_15545;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_183_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_183_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_183_tag <= _GEN_6327;
      end
    end else begin
      btb_183_tag <= _GEN_6327;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_183_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_183_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_183_target_address <= _GEN_11303;
      end
    end else begin
      btb_183_target_address <= _GEN_11303;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_183_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_183_bht <= 2'h1;
        end else begin
          btb_183_bht <= 2'h0;
        end
      end else begin
        btb_183_bht <= _GEN_11305;
      end
    end else begin
      btb_183_bht <= _GEN_11305;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_184_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_184_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_184_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_184_valid <= _GEN_15546;
      end
    end else begin
      btb_184_valid <= _GEN_15546;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_184_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_184_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_184_tag <= _GEN_6328;
      end
    end else begin
      btb_184_tag <= _GEN_6328;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_184_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_184_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_184_target_address <= _GEN_11306;
      end
    end else begin
      btb_184_target_address <= _GEN_11306;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_184_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_184_bht <= 2'h1;
        end else begin
          btb_184_bht <= 2'h0;
        end
      end else begin
        btb_184_bht <= _GEN_11308;
      end
    end else begin
      btb_184_bht <= _GEN_11308;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_185_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_185_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_185_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_185_valid <= _GEN_15547;
      end
    end else begin
      btb_185_valid <= _GEN_15547;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_185_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_185_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_185_tag <= _GEN_6329;
      end
    end else begin
      btb_185_tag <= _GEN_6329;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_185_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_185_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_185_target_address <= _GEN_11309;
      end
    end else begin
      btb_185_target_address <= _GEN_11309;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_185_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hb9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_185_bht <= 2'h1;
        end else begin
          btb_185_bht <= 2'h0;
        end
      end else begin
        btb_185_bht <= _GEN_11311;
      end
    end else begin
      btb_185_bht <= _GEN_11311;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_186_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_186_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_186_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_186_valid <= _GEN_15548;
      end
    end else begin
      btb_186_valid <= _GEN_15548;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_186_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hba == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_186_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_186_tag <= _GEN_6330;
      end
    end else begin
      btb_186_tag <= _GEN_6330;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_186_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hba == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_186_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_186_target_address <= _GEN_11312;
      end
    end else begin
      btb_186_target_address <= _GEN_11312;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_186_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hba == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_186_bht <= 2'h1;
        end else begin
          btb_186_bht <= 2'h0;
        end
      end else begin
        btb_186_bht <= _GEN_11314;
      end
    end else begin
      btb_186_bht <= _GEN_11314;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_187_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_187_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_187_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_187_valid <= _GEN_15549;
      end
    end else begin
      btb_187_valid <= _GEN_15549;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_187_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_187_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_187_tag <= _GEN_6331;
      end
    end else begin
      btb_187_tag <= _GEN_6331;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_187_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_187_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_187_target_address <= _GEN_11315;
      end
    end else begin
      btb_187_target_address <= _GEN_11315;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_187_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_187_bht <= 2'h1;
        end else begin
          btb_187_bht <= 2'h0;
        end
      end else begin
        btb_187_bht <= _GEN_11317;
      end
    end else begin
      btb_187_bht <= _GEN_11317;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_188_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_188_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_188_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_188_valid <= _GEN_15550;
      end
    end else begin
      btb_188_valid <= _GEN_15550;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_188_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_188_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_188_tag <= _GEN_6332;
      end
    end else begin
      btb_188_tag <= _GEN_6332;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_188_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_188_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_188_target_address <= _GEN_11318;
      end
    end else begin
      btb_188_target_address <= _GEN_11318;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_188_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_188_bht <= 2'h1;
        end else begin
          btb_188_bht <= 2'h0;
        end
      end else begin
        btb_188_bht <= _GEN_11320;
      end
    end else begin
      btb_188_bht <= _GEN_11320;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_189_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_189_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_189_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_189_valid <= _GEN_15551;
      end
    end else begin
      btb_189_valid <= _GEN_15551;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_189_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_189_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_189_tag <= _GEN_6333;
      end
    end else begin
      btb_189_tag <= _GEN_6333;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_189_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_189_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_189_target_address <= _GEN_11321;
      end
    end else begin
      btb_189_target_address <= _GEN_11321;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_189_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_189_bht <= 2'h1;
        end else begin
          btb_189_bht <= 2'h0;
        end
      end else begin
        btb_189_bht <= _GEN_11323;
      end
    end else begin
      btb_189_bht <= _GEN_11323;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_190_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_190_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_190_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_190_valid <= _GEN_15552;
      end
    end else begin
      btb_190_valid <= _GEN_15552;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_190_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbe == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_190_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_190_tag <= _GEN_6334;
      end
    end else begin
      btb_190_tag <= _GEN_6334;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_190_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbe == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_190_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_190_target_address <= _GEN_11324;
      end
    end else begin
      btb_190_target_address <= _GEN_11324;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_190_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbe == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_190_bht <= 2'h1;
        end else begin
          btb_190_bht <= 2'h0;
        end
      end else begin
        btb_190_bht <= _GEN_11326;
      end
    end else begin
      btb_190_bht <= _GEN_11326;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_191_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_191_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_191_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_191_valid <= _GEN_15553;
      end
    end else begin
      btb_191_valid <= _GEN_15553;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_191_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_191_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_191_tag <= _GEN_6335;
      end
    end else begin
      btb_191_tag <= _GEN_6335;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_191_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_191_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_191_target_address <= _GEN_11327;
      end
    end else begin
      btb_191_target_address <= _GEN_11327;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_191_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hbf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_191_bht <= 2'h1;
        end else begin
          btb_191_bht <= 2'h0;
        end
      end else begin
        btb_191_bht <= _GEN_11329;
      end
    end else begin
      btb_191_bht <= _GEN_11329;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_192_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_192_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_192_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_192_valid <= _GEN_15554;
      end
    end else begin
      btb_192_valid <= _GEN_15554;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_192_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_192_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_192_tag <= _GEN_6336;
      end
    end else begin
      btb_192_tag <= _GEN_6336;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_192_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_192_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_192_target_address <= _GEN_11330;
      end
    end else begin
      btb_192_target_address <= _GEN_11330;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_192_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_192_bht <= 2'h1;
        end else begin
          btb_192_bht <= 2'h0;
        end
      end else begin
        btb_192_bht <= _GEN_11332;
      end
    end else begin
      btb_192_bht <= _GEN_11332;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_193_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_193_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_193_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_193_valid <= _GEN_15555;
      end
    end else begin
      btb_193_valid <= _GEN_15555;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_193_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_193_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_193_tag <= _GEN_6337;
      end
    end else begin
      btb_193_tag <= _GEN_6337;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_193_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_193_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_193_target_address <= _GEN_11333;
      end
    end else begin
      btb_193_target_address <= _GEN_11333;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_193_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_193_bht <= 2'h1;
        end else begin
          btb_193_bht <= 2'h0;
        end
      end else begin
        btb_193_bht <= _GEN_11335;
      end
    end else begin
      btb_193_bht <= _GEN_11335;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_194_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_194_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_194_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_194_valid <= _GEN_15556;
      end
    end else begin
      btb_194_valid <= _GEN_15556;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_194_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_194_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_194_tag <= _GEN_6338;
      end
    end else begin
      btb_194_tag <= _GEN_6338;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_194_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_194_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_194_target_address <= _GEN_11336;
      end
    end else begin
      btb_194_target_address <= _GEN_11336;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_194_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_194_bht <= 2'h1;
        end else begin
          btb_194_bht <= 2'h0;
        end
      end else begin
        btb_194_bht <= _GEN_11338;
      end
    end else begin
      btb_194_bht <= _GEN_11338;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_195_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_195_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_195_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_195_valid <= _GEN_15557;
      end
    end else begin
      btb_195_valid <= _GEN_15557;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_195_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_195_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_195_tag <= _GEN_6339;
      end
    end else begin
      btb_195_tag <= _GEN_6339;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_195_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_195_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_195_target_address <= _GEN_11339;
      end
    end else begin
      btb_195_target_address <= _GEN_11339;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_195_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_195_bht <= 2'h1;
        end else begin
          btb_195_bht <= 2'h0;
        end
      end else begin
        btb_195_bht <= _GEN_11341;
      end
    end else begin
      btb_195_bht <= _GEN_11341;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_196_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_196_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_196_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_196_valid <= _GEN_15558;
      end
    end else begin
      btb_196_valid <= _GEN_15558;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_196_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_196_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_196_tag <= _GEN_6340;
      end
    end else begin
      btb_196_tag <= _GEN_6340;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_196_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_196_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_196_target_address <= _GEN_11342;
      end
    end else begin
      btb_196_target_address <= _GEN_11342;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_196_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_196_bht <= 2'h1;
        end else begin
          btb_196_bht <= 2'h0;
        end
      end else begin
        btb_196_bht <= _GEN_11344;
      end
    end else begin
      btb_196_bht <= _GEN_11344;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_197_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_197_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_197_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_197_valid <= _GEN_15559;
      end
    end else begin
      btb_197_valid <= _GEN_15559;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_197_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_197_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_197_tag <= _GEN_6341;
      end
    end else begin
      btb_197_tag <= _GEN_6341;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_197_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_197_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_197_target_address <= _GEN_11345;
      end
    end else begin
      btb_197_target_address <= _GEN_11345;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_197_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_197_bht <= 2'h1;
        end else begin
          btb_197_bht <= 2'h0;
        end
      end else begin
        btb_197_bht <= _GEN_11347;
      end
    end else begin
      btb_197_bht <= _GEN_11347;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_198_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_198_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_198_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_198_valid <= _GEN_15560;
      end
    end else begin
      btb_198_valid <= _GEN_15560;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_198_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_198_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_198_tag <= _GEN_6342;
      end
    end else begin
      btb_198_tag <= _GEN_6342;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_198_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_198_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_198_target_address <= _GEN_11348;
      end
    end else begin
      btb_198_target_address <= _GEN_11348;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_198_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_198_bht <= 2'h1;
        end else begin
          btb_198_bht <= 2'h0;
        end
      end else begin
        btb_198_bht <= _GEN_11350;
      end
    end else begin
      btb_198_bht <= _GEN_11350;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_199_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_199_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_199_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_199_valid <= _GEN_15561;
      end
    end else begin
      btb_199_valid <= _GEN_15561;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_199_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_199_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_199_tag <= _GEN_6343;
      end
    end else begin
      btb_199_tag <= _GEN_6343;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_199_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_199_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_199_target_address <= _GEN_11351;
      end
    end else begin
      btb_199_target_address <= _GEN_11351;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_199_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_199_bht <= 2'h1;
        end else begin
          btb_199_bht <= 2'h0;
        end
      end else begin
        btb_199_bht <= _GEN_11353;
      end
    end else begin
      btb_199_bht <= _GEN_11353;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_200_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_200_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_200_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_200_valid <= _GEN_15562;
      end
    end else begin
      btb_200_valid <= _GEN_15562;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_200_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_200_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_200_tag <= _GEN_6344;
      end
    end else begin
      btb_200_tag <= _GEN_6344;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_200_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_200_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_200_target_address <= _GEN_11354;
      end
    end else begin
      btb_200_target_address <= _GEN_11354;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_200_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_200_bht <= 2'h1;
        end else begin
          btb_200_bht <= 2'h0;
        end
      end else begin
        btb_200_bht <= _GEN_11356;
      end
    end else begin
      btb_200_bht <= _GEN_11356;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_201_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_201_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_201_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_201_valid <= _GEN_15563;
      end
    end else begin
      btb_201_valid <= _GEN_15563;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_201_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_201_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_201_tag <= _GEN_6345;
      end
    end else begin
      btb_201_tag <= _GEN_6345;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_201_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_201_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_201_target_address <= _GEN_11357;
      end
    end else begin
      btb_201_target_address <= _GEN_11357;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_201_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hc9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_201_bht <= 2'h1;
        end else begin
          btb_201_bht <= 2'h0;
        end
      end else begin
        btb_201_bht <= _GEN_11359;
      end
    end else begin
      btb_201_bht <= _GEN_11359;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_202_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_202_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_202_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_202_valid <= _GEN_15564;
      end
    end else begin
      btb_202_valid <= _GEN_15564;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_202_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hca == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_202_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_202_tag <= _GEN_6346;
      end
    end else begin
      btb_202_tag <= _GEN_6346;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_202_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hca == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_202_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_202_target_address <= _GEN_11360;
      end
    end else begin
      btb_202_target_address <= _GEN_11360;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_202_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hca == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_202_bht <= 2'h1;
        end else begin
          btb_202_bht <= 2'h0;
        end
      end else begin
        btb_202_bht <= _GEN_11362;
      end
    end else begin
      btb_202_bht <= _GEN_11362;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_203_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_203_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_203_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_203_valid <= _GEN_15565;
      end
    end else begin
      btb_203_valid <= _GEN_15565;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_203_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_203_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_203_tag <= _GEN_6347;
      end
    end else begin
      btb_203_tag <= _GEN_6347;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_203_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_203_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_203_target_address <= _GEN_11363;
      end
    end else begin
      btb_203_target_address <= _GEN_11363;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_203_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_203_bht <= 2'h1;
        end else begin
          btb_203_bht <= 2'h0;
        end
      end else begin
        btb_203_bht <= _GEN_11365;
      end
    end else begin
      btb_203_bht <= _GEN_11365;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_204_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_204_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_204_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_204_valid <= _GEN_15566;
      end
    end else begin
      btb_204_valid <= _GEN_15566;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_204_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_204_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_204_tag <= _GEN_6348;
      end
    end else begin
      btb_204_tag <= _GEN_6348;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_204_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_204_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_204_target_address <= _GEN_11366;
      end
    end else begin
      btb_204_target_address <= _GEN_11366;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_204_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_204_bht <= 2'h1;
        end else begin
          btb_204_bht <= 2'h0;
        end
      end else begin
        btb_204_bht <= _GEN_11368;
      end
    end else begin
      btb_204_bht <= _GEN_11368;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_205_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_205_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_205_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_205_valid <= _GEN_15567;
      end
    end else begin
      btb_205_valid <= _GEN_15567;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_205_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_205_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_205_tag <= _GEN_6349;
      end
    end else begin
      btb_205_tag <= _GEN_6349;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_205_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_205_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_205_target_address <= _GEN_11369;
      end
    end else begin
      btb_205_target_address <= _GEN_11369;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_205_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_205_bht <= 2'h1;
        end else begin
          btb_205_bht <= 2'h0;
        end
      end else begin
        btb_205_bht <= _GEN_11371;
      end
    end else begin
      btb_205_bht <= _GEN_11371;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_206_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_206_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_206_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_206_valid <= _GEN_15568;
      end
    end else begin
      btb_206_valid <= _GEN_15568;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_206_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hce == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_206_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_206_tag <= _GEN_6350;
      end
    end else begin
      btb_206_tag <= _GEN_6350;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_206_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hce == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_206_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_206_target_address <= _GEN_11372;
      end
    end else begin
      btb_206_target_address <= _GEN_11372;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_206_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hce == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_206_bht <= 2'h1;
        end else begin
          btb_206_bht <= 2'h0;
        end
      end else begin
        btb_206_bht <= _GEN_11374;
      end
    end else begin
      btb_206_bht <= _GEN_11374;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_207_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_207_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_207_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_207_valid <= _GEN_15569;
      end
    end else begin
      btb_207_valid <= _GEN_15569;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_207_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_207_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_207_tag <= _GEN_6351;
      end
    end else begin
      btb_207_tag <= _GEN_6351;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_207_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_207_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_207_target_address <= _GEN_11375;
      end
    end else begin
      btb_207_target_address <= _GEN_11375;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_207_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hcf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_207_bht <= 2'h1;
        end else begin
          btb_207_bht <= 2'h0;
        end
      end else begin
        btb_207_bht <= _GEN_11377;
      end
    end else begin
      btb_207_bht <= _GEN_11377;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_208_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_208_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_208_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_208_valid <= _GEN_15570;
      end
    end else begin
      btb_208_valid <= _GEN_15570;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_208_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_208_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_208_tag <= _GEN_6352;
      end
    end else begin
      btb_208_tag <= _GEN_6352;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_208_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_208_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_208_target_address <= _GEN_11378;
      end
    end else begin
      btb_208_target_address <= _GEN_11378;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_208_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_208_bht <= 2'h1;
        end else begin
          btb_208_bht <= 2'h0;
        end
      end else begin
        btb_208_bht <= _GEN_11380;
      end
    end else begin
      btb_208_bht <= _GEN_11380;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_209_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_209_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_209_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_209_valid <= _GEN_15571;
      end
    end else begin
      btb_209_valid <= _GEN_15571;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_209_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_209_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_209_tag <= _GEN_6353;
      end
    end else begin
      btb_209_tag <= _GEN_6353;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_209_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_209_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_209_target_address <= _GEN_11381;
      end
    end else begin
      btb_209_target_address <= _GEN_11381;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_209_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_209_bht <= 2'h1;
        end else begin
          btb_209_bht <= 2'h0;
        end
      end else begin
        btb_209_bht <= _GEN_11383;
      end
    end else begin
      btb_209_bht <= _GEN_11383;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_210_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_210_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_210_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_210_valid <= _GEN_15572;
      end
    end else begin
      btb_210_valid <= _GEN_15572;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_210_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_210_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_210_tag <= _GEN_6354;
      end
    end else begin
      btb_210_tag <= _GEN_6354;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_210_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_210_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_210_target_address <= _GEN_11384;
      end
    end else begin
      btb_210_target_address <= _GEN_11384;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_210_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_210_bht <= 2'h1;
        end else begin
          btb_210_bht <= 2'h0;
        end
      end else begin
        btb_210_bht <= _GEN_11386;
      end
    end else begin
      btb_210_bht <= _GEN_11386;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_211_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_211_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_211_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_211_valid <= _GEN_15573;
      end
    end else begin
      btb_211_valid <= _GEN_15573;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_211_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_211_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_211_tag <= _GEN_6355;
      end
    end else begin
      btb_211_tag <= _GEN_6355;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_211_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_211_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_211_target_address <= _GEN_11387;
      end
    end else begin
      btb_211_target_address <= _GEN_11387;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_211_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_211_bht <= 2'h1;
        end else begin
          btb_211_bht <= 2'h0;
        end
      end else begin
        btb_211_bht <= _GEN_11389;
      end
    end else begin
      btb_211_bht <= _GEN_11389;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_212_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_212_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_212_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_212_valid <= _GEN_15574;
      end
    end else begin
      btb_212_valid <= _GEN_15574;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_212_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_212_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_212_tag <= _GEN_6356;
      end
    end else begin
      btb_212_tag <= _GEN_6356;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_212_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_212_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_212_target_address <= _GEN_11390;
      end
    end else begin
      btb_212_target_address <= _GEN_11390;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_212_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_212_bht <= 2'h1;
        end else begin
          btb_212_bht <= 2'h0;
        end
      end else begin
        btb_212_bht <= _GEN_11392;
      end
    end else begin
      btb_212_bht <= _GEN_11392;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_213_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_213_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_213_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_213_valid <= _GEN_15575;
      end
    end else begin
      btb_213_valid <= _GEN_15575;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_213_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_213_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_213_tag <= _GEN_6357;
      end
    end else begin
      btb_213_tag <= _GEN_6357;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_213_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_213_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_213_target_address <= _GEN_11393;
      end
    end else begin
      btb_213_target_address <= _GEN_11393;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_213_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_213_bht <= 2'h1;
        end else begin
          btb_213_bht <= 2'h0;
        end
      end else begin
        btb_213_bht <= _GEN_11395;
      end
    end else begin
      btb_213_bht <= _GEN_11395;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_214_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_214_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_214_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_214_valid <= _GEN_15576;
      end
    end else begin
      btb_214_valid <= _GEN_15576;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_214_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_214_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_214_tag <= _GEN_6358;
      end
    end else begin
      btb_214_tag <= _GEN_6358;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_214_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_214_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_214_target_address <= _GEN_11396;
      end
    end else begin
      btb_214_target_address <= _GEN_11396;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_214_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_214_bht <= 2'h1;
        end else begin
          btb_214_bht <= 2'h0;
        end
      end else begin
        btb_214_bht <= _GEN_11398;
      end
    end else begin
      btb_214_bht <= _GEN_11398;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_215_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_215_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_215_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_215_valid <= _GEN_15577;
      end
    end else begin
      btb_215_valid <= _GEN_15577;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_215_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_215_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_215_tag <= _GEN_6359;
      end
    end else begin
      btb_215_tag <= _GEN_6359;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_215_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_215_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_215_target_address <= _GEN_11399;
      end
    end else begin
      btb_215_target_address <= _GEN_11399;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_215_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_215_bht <= 2'h1;
        end else begin
          btb_215_bht <= 2'h0;
        end
      end else begin
        btb_215_bht <= _GEN_11401;
      end
    end else begin
      btb_215_bht <= _GEN_11401;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_216_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_216_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_216_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_216_valid <= _GEN_15578;
      end
    end else begin
      btb_216_valid <= _GEN_15578;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_216_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_216_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_216_tag <= _GEN_6360;
      end
    end else begin
      btb_216_tag <= _GEN_6360;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_216_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_216_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_216_target_address <= _GEN_11402;
      end
    end else begin
      btb_216_target_address <= _GEN_11402;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_216_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_216_bht <= 2'h1;
        end else begin
          btb_216_bht <= 2'h0;
        end
      end else begin
        btb_216_bht <= _GEN_11404;
      end
    end else begin
      btb_216_bht <= _GEN_11404;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_217_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_217_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_217_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_217_valid <= _GEN_15579;
      end
    end else begin
      btb_217_valid <= _GEN_15579;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_217_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_217_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_217_tag <= _GEN_6361;
      end
    end else begin
      btb_217_tag <= _GEN_6361;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_217_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_217_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_217_target_address <= _GEN_11405;
      end
    end else begin
      btb_217_target_address <= _GEN_11405;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_217_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hd9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_217_bht <= 2'h1;
        end else begin
          btb_217_bht <= 2'h0;
        end
      end else begin
        btb_217_bht <= _GEN_11407;
      end
    end else begin
      btb_217_bht <= _GEN_11407;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_218_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_218_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_218_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_218_valid <= _GEN_15580;
      end
    end else begin
      btb_218_valid <= _GEN_15580;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_218_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hda == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_218_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_218_tag <= _GEN_6362;
      end
    end else begin
      btb_218_tag <= _GEN_6362;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_218_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hda == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_218_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_218_target_address <= _GEN_11408;
      end
    end else begin
      btb_218_target_address <= _GEN_11408;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_218_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hda == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_218_bht <= 2'h1;
        end else begin
          btb_218_bht <= 2'h0;
        end
      end else begin
        btb_218_bht <= _GEN_11410;
      end
    end else begin
      btb_218_bht <= _GEN_11410;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_219_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_219_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_219_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_219_valid <= _GEN_15581;
      end
    end else begin
      btb_219_valid <= _GEN_15581;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_219_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_219_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_219_tag <= _GEN_6363;
      end
    end else begin
      btb_219_tag <= _GEN_6363;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_219_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_219_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_219_target_address <= _GEN_11411;
      end
    end else begin
      btb_219_target_address <= _GEN_11411;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_219_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_219_bht <= 2'h1;
        end else begin
          btb_219_bht <= 2'h0;
        end
      end else begin
        btb_219_bht <= _GEN_11413;
      end
    end else begin
      btb_219_bht <= _GEN_11413;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_220_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_220_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_220_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_220_valid <= _GEN_15582;
      end
    end else begin
      btb_220_valid <= _GEN_15582;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_220_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_220_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_220_tag <= _GEN_6364;
      end
    end else begin
      btb_220_tag <= _GEN_6364;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_220_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_220_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_220_target_address <= _GEN_11414;
      end
    end else begin
      btb_220_target_address <= _GEN_11414;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_220_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_220_bht <= 2'h1;
        end else begin
          btb_220_bht <= 2'h0;
        end
      end else begin
        btb_220_bht <= _GEN_11416;
      end
    end else begin
      btb_220_bht <= _GEN_11416;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_221_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_221_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_221_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_221_valid <= _GEN_15583;
      end
    end else begin
      btb_221_valid <= _GEN_15583;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_221_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_221_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_221_tag <= _GEN_6365;
      end
    end else begin
      btb_221_tag <= _GEN_6365;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_221_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_221_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_221_target_address <= _GEN_11417;
      end
    end else begin
      btb_221_target_address <= _GEN_11417;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_221_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_221_bht <= 2'h1;
        end else begin
          btb_221_bht <= 2'h0;
        end
      end else begin
        btb_221_bht <= _GEN_11419;
      end
    end else begin
      btb_221_bht <= _GEN_11419;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_222_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_222_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_222_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_222_valid <= _GEN_15584;
      end
    end else begin
      btb_222_valid <= _GEN_15584;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_222_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hde == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_222_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_222_tag <= _GEN_6366;
      end
    end else begin
      btb_222_tag <= _GEN_6366;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_222_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hde == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_222_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_222_target_address <= _GEN_11420;
      end
    end else begin
      btb_222_target_address <= _GEN_11420;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_222_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hde == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_222_bht <= 2'h1;
        end else begin
          btb_222_bht <= 2'h0;
        end
      end else begin
        btb_222_bht <= _GEN_11422;
      end
    end else begin
      btb_222_bht <= _GEN_11422;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_223_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_223_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_223_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_223_valid <= _GEN_15585;
      end
    end else begin
      btb_223_valid <= _GEN_15585;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_223_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_223_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_223_tag <= _GEN_6367;
      end
    end else begin
      btb_223_tag <= _GEN_6367;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_223_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_223_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_223_target_address <= _GEN_11423;
      end
    end else begin
      btb_223_target_address <= _GEN_11423;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_223_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hdf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_223_bht <= 2'h1;
        end else begin
          btb_223_bht <= 2'h0;
        end
      end else begin
        btb_223_bht <= _GEN_11425;
      end
    end else begin
      btb_223_bht <= _GEN_11425;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_224_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_224_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_224_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_224_valid <= _GEN_15586;
      end
    end else begin
      btb_224_valid <= _GEN_15586;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_224_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_224_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_224_tag <= _GEN_6368;
      end
    end else begin
      btb_224_tag <= _GEN_6368;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_224_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_224_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_224_target_address <= _GEN_11426;
      end
    end else begin
      btb_224_target_address <= _GEN_11426;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_224_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_224_bht <= 2'h1;
        end else begin
          btb_224_bht <= 2'h0;
        end
      end else begin
        btb_224_bht <= _GEN_11428;
      end
    end else begin
      btb_224_bht <= _GEN_11428;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_225_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_225_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_225_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_225_valid <= _GEN_15587;
      end
    end else begin
      btb_225_valid <= _GEN_15587;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_225_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_225_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_225_tag <= _GEN_6369;
      end
    end else begin
      btb_225_tag <= _GEN_6369;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_225_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_225_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_225_target_address <= _GEN_11429;
      end
    end else begin
      btb_225_target_address <= _GEN_11429;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_225_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_225_bht <= 2'h1;
        end else begin
          btb_225_bht <= 2'h0;
        end
      end else begin
        btb_225_bht <= _GEN_11431;
      end
    end else begin
      btb_225_bht <= _GEN_11431;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_226_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_226_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_226_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_226_valid <= _GEN_15588;
      end
    end else begin
      btb_226_valid <= _GEN_15588;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_226_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_226_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_226_tag <= _GEN_6370;
      end
    end else begin
      btb_226_tag <= _GEN_6370;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_226_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_226_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_226_target_address <= _GEN_11432;
      end
    end else begin
      btb_226_target_address <= _GEN_11432;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_226_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_226_bht <= 2'h1;
        end else begin
          btb_226_bht <= 2'h0;
        end
      end else begin
        btb_226_bht <= _GEN_11434;
      end
    end else begin
      btb_226_bht <= _GEN_11434;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_227_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_227_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_227_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_227_valid <= _GEN_15589;
      end
    end else begin
      btb_227_valid <= _GEN_15589;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_227_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_227_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_227_tag <= _GEN_6371;
      end
    end else begin
      btb_227_tag <= _GEN_6371;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_227_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_227_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_227_target_address <= _GEN_11435;
      end
    end else begin
      btb_227_target_address <= _GEN_11435;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_227_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_227_bht <= 2'h1;
        end else begin
          btb_227_bht <= 2'h0;
        end
      end else begin
        btb_227_bht <= _GEN_11437;
      end
    end else begin
      btb_227_bht <= _GEN_11437;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_228_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_228_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_228_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_228_valid <= _GEN_15590;
      end
    end else begin
      btb_228_valid <= _GEN_15590;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_228_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_228_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_228_tag <= _GEN_6372;
      end
    end else begin
      btb_228_tag <= _GEN_6372;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_228_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_228_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_228_target_address <= _GEN_11438;
      end
    end else begin
      btb_228_target_address <= _GEN_11438;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_228_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_228_bht <= 2'h1;
        end else begin
          btb_228_bht <= 2'h0;
        end
      end else begin
        btb_228_bht <= _GEN_11440;
      end
    end else begin
      btb_228_bht <= _GEN_11440;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_229_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_229_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_229_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_229_valid <= _GEN_15591;
      end
    end else begin
      btb_229_valid <= _GEN_15591;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_229_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_229_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_229_tag <= _GEN_6373;
      end
    end else begin
      btb_229_tag <= _GEN_6373;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_229_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_229_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_229_target_address <= _GEN_11441;
      end
    end else begin
      btb_229_target_address <= _GEN_11441;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_229_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_229_bht <= 2'h1;
        end else begin
          btb_229_bht <= 2'h0;
        end
      end else begin
        btb_229_bht <= _GEN_11443;
      end
    end else begin
      btb_229_bht <= _GEN_11443;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_230_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_230_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_230_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_230_valid <= _GEN_15592;
      end
    end else begin
      btb_230_valid <= _GEN_15592;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_230_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_230_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_230_tag <= _GEN_6374;
      end
    end else begin
      btb_230_tag <= _GEN_6374;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_230_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_230_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_230_target_address <= _GEN_11444;
      end
    end else begin
      btb_230_target_address <= _GEN_11444;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_230_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_230_bht <= 2'h1;
        end else begin
          btb_230_bht <= 2'h0;
        end
      end else begin
        btb_230_bht <= _GEN_11446;
      end
    end else begin
      btb_230_bht <= _GEN_11446;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_231_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_231_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_231_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_231_valid <= _GEN_15593;
      end
    end else begin
      btb_231_valid <= _GEN_15593;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_231_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_231_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_231_tag <= _GEN_6375;
      end
    end else begin
      btb_231_tag <= _GEN_6375;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_231_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_231_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_231_target_address <= _GEN_11447;
      end
    end else begin
      btb_231_target_address <= _GEN_11447;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_231_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_231_bht <= 2'h1;
        end else begin
          btb_231_bht <= 2'h0;
        end
      end else begin
        btb_231_bht <= _GEN_11449;
      end
    end else begin
      btb_231_bht <= _GEN_11449;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_232_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_232_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_232_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_232_valid <= _GEN_15594;
      end
    end else begin
      btb_232_valid <= _GEN_15594;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_232_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_232_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_232_tag <= _GEN_6376;
      end
    end else begin
      btb_232_tag <= _GEN_6376;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_232_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_232_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_232_target_address <= _GEN_11450;
      end
    end else begin
      btb_232_target_address <= _GEN_11450;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_232_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_232_bht <= 2'h1;
        end else begin
          btb_232_bht <= 2'h0;
        end
      end else begin
        btb_232_bht <= _GEN_11452;
      end
    end else begin
      btb_232_bht <= _GEN_11452;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_233_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_233_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_233_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_233_valid <= _GEN_15595;
      end
    end else begin
      btb_233_valid <= _GEN_15595;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_233_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_233_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_233_tag <= _GEN_6377;
      end
    end else begin
      btb_233_tag <= _GEN_6377;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_233_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_233_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_233_target_address <= _GEN_11453;
      end
    end else begin
      btb_233_target_address <= _GEN_11453;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_233_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'he9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_233_bht <= 2'h1;
        end else begin
          btb_233_bht <= 2'h0;
        end
      end else begin
        btb_233_bht <= _GEN_11455;
      end
    end else begin
      btb_233_bht <= _GEN_11455;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_234_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_234_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_234_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_234_valid <= _GEN_15596;
      end
    end else begin
      btb_234_valid <= _GEN_15596;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_234_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hea == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_234_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_234_tag <= _GEN_6378;
      end
    end else begin
      btb_234_tag <= _GEN_6378;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_234_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hea == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_234_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_234_target_address <= _GEN_11456;
      end
    end else begin
      btb_234_target_address <= _GEN_11456;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_234_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hea == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_234_bht <= 2'h1;
        end else begin
          btb_234_bht <= 2'h0;
        end
      end else begin
        btb_234_bht <= _GEN_11458;
      end
    end else begin
      btb_234_bht <= _GEN_11458;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_235_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_235_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_235_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_235_valid <= _GEN_15597;
      end
    end else begin
      btb_235_valid <= _GEN_15597;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_235_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'heb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_235_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_235_tag <= _GEN_6379;
      end
    end else begin
      btb_235_tag <= _GEN_6379;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_235_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'heb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_235_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_235_target_address <= _GEN_11459;
      end
    end else begin
      btb_235_target_address <= _GEN_11459;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_235_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'heb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_235_bht <= 2'h1;
        end else begin
          btb_235_bht <= 2'h0;
        end
      end else begin
        btb_235_bht <= _GEN_11461;
      end
    end else begin
      btb_235_bht <= _GEN_11461;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_236_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_236_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_236_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_236_valid <= _GEN_15598;
      end
    end else begin
      btb_236_valid <= _GEN_15598;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_236_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hec == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_236_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_236_tag <= _GEN_6380;
      end
    end else begin
      btb_236_tag <= _GEN_6380;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_236_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hec == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_236_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_236_target_address <= _GEN_11462;
      end
    end else begin
      btb_236_target_address <= _GEN_11462;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_236_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hec == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_236_bht <= 2'h1;
        end else begin
          btb_236_bht <= 2'h0;
        end
      end else begin
        btb_236_bht <= _GEN_11464;
      end
    end else begin
      btb_236_bht <= _GEN_11464;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_237_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_237_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_237_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_237_valid <= _GEN_15599;
      end
    end else begin
      btb_237_valid <= _GEN_15599;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_237_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hed == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_237_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_237_tag <= _GEN_6381;
      end
    end else begin
      btb_237_tag <= _GEN_6381;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_237_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hed == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_237_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_237_target_address <= _GEN_11465;
      end
    end else begin
      btb_237_target_address <= _GEN_11465;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_237_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hed == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_237_bht <= 2'h1;
        end else begin
          btb_237_bht <= 2'h0;
        end
      end else begin
        btb_237_bht <= _GEN_11467;
      end
    end else begin
      btb_237_bht <= _GEN_11467;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_238_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_238_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_238_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_238_valid <= _GEN_15600;
      end
    end else begin
      btb_238_valid <= _GEN_15600;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_238_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hee == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_238_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_238_tag <= _GEN_6382;
      end
    end else begin
      btb_238_tag <= _GEN_6382;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_238_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hee == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_238_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_238_target_address <= _GEN_11468;
      end
    end else begin
      btb_238_target_address <= _GEN_11468;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_238_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hee == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_238_bht <= 2'h1;
        end else begin
          btb_238_bht <= 2'h0;
        end
      end else begin
        btb_238_bht <= _GEN_11470;
      end
    end else begin
      btb_238_bht <= _GEN_11470;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_239_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_239_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_239_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_239_valid <= _GEN_15601;
      end
    end else begin
      btb_239_valid <= _GEN_15601;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_239_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hef == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_239_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_239_tag <= _GEN_6383;
      end
    end else begin
      btb_239_tag <= _GEN_6383;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_239_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hef == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_239_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_239_target_address <= _GEN_11471;
      end
    end else begin
      btb_239_target_address <= _GEN_11471;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_239_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hef == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_239_bht <= 2'h1;
        end else begin
          btb_239_bht <= 2'h0;
        end
      end else begin
        btb_239_bht <= _GEN_11473;
      end
    end else begin
      btb_239_bht <= _GEN_11473;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_240_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_240_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_240_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_240_valid <= _GEN_15602;
      end
    end else begin
      btb_240_valid <= _GEN_15602;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_240_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_240_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_240_tag <= _GEN_6384;
      end
    end else begin
      btb_240_tag <= _GEN_6384;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_240_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_240_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_240_target_address <= _GEN_11474;
      end
    end else begin
      btb_240_target_address <= _GEN_11474;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_240_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_240_bht <= 2'h1;
        end else begin
          btb_240_bht <= 2'h0;
        end
      end else begin
        btb_240_bht <= _GEN_11476;
      end
    end else begin
      btb_240_bht <= _GEN_11476;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_241_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_241_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_241_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_241_valid <= _GEN_15603;
      end
    end else begin
      btb_241_valid <= _GEN_15603;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_241_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_241_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_241_tag <= _GEN_6385;
      end
    end else begin
      btb_241_tag <= _GEN_6385;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_241_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_241_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_241_target_address <= _GEN_11477;
      end
    end else begin
      btb_241_target_address <= _GEN_11477;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_241_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_241_bht <= 2'h1;
        end else begin
          btb_241_bht <= 2'h0;
        end
      end else begin
        btb_241_bht <= _GEN_11479;
      end
    end else begin
      btb_241_bht <= _GEN_11479;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_242_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_242_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_242_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_242_valid <= _GEN_15604;
      end
    end else begin
      btb_242_valid <= _GEN_15604;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_242_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_242_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_242_tag <= _GEN_6386;
      end
    end else begin
      btb_242_tag <= _GEN_6386;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_242_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_242_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_242_target_address <= _GEN_11480;
      end
    end else begin
      btb_242_target_address <= _GEN_11480;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_242_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_242_bht <= 2'h1;
        end else begin
          btb_242_bht <= 2'h0;
        end
      end else begin
        btb_242_bht <= _GEN_11482;
      end
    end else begin
      btb_242_bht <= _GEN_11482;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_243_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_243_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_243_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_243_valid <= _GEN_15605;
      end
    end else begin
      btb_243_valid <= _GEN_15605;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_243_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_243_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_243_tag <= _GEN_6387;
      end
    end else begin
      btb_243_tag <= _GEN_6387;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_243_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_243_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_243_target_address <= _GEN_11483;
      end
    end else begin
      btb_243_target_address <= _GEN_11483;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_243_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_243_bht <= 2'h1;
        end else begin
          btb_243_bht <= 2'h0;
        end
      end else begin
        btb_243_bht <= _GEN_11485;
      end
    end else begin
      btb_243_bht <= _GEN_11485;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_244_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_244_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_244_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_244_valid <= _GEN_15606;
      end
    end else begin
      btb_244_valid <= _GEN_15606;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_244_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_244_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_244_tag <= _GEN_6388;
      end
    end else begin
      btb_244_tag <= _GEN_6388;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_244_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_244_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_244_target_address <= _GEN_11486;
      end
    end else begin
      btb_244_target_address <= _GEN_11486;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_244_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_244_bht <= 2'h1;
        end else begin
          btb_244_bht <= 2'h0;
        end
      end else begin
        btb_244_bht <= _GEN_11488;
      end
    end else begin
      btb_244_bht <= _GEN_11488;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_245_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_245_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_245_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_245_valid <= _GEN_15607;
      end
    end else begin
      btb_245_valid <= _GEN_15607;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_245_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_245_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_245_tag <= _GEN_6389;
      end
    end else begin
      btb_245_tag <= _GEN_6389;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_245_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_245_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_245_target_address <= _GEN_11489;
      end
    end else begin
      btb_245_target_address <= _GEN_11489;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_245_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_245_bht <= 2'h1;
        end else begin
          btb_245_bht <= 2'h0;
        end
      end else begin
        btb_245_bht <= _GEN_11491;
      end
    end else begin
      btb_245_bht <= _GEN_11491;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_246_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_246_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_246_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_246_valid <= _GEN_15608;
      end
    end else begin
      btb_246_valid <= _GEN_15608;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_246_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_246_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_246_tag <= _GEN_6390;
      end
    end else begin
      btb_246_tag <= _GEN_6390;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_246_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_246_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_246_target_address <= _GEN_11492;
      end
    end else begin
      btb_246_target_address <= _GEN_11492;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_246_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_246_bht <= 2'h1;
        end else begin
          btb_246_bht <= 2'h0;
        end
      end else begin
        btb_246_bht <= _GEN_11494;
      end
    end else begin
      btb_246_bht <= _GEN_11494;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_247_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_247_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_247_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_247_valid <= _GEN_15609;
      end
    end else begin
      btb_247_valid <= _GEN_15609;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_247_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_247_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_247_tag <= _GEN_6391;
      end
    end else begin
      btb_247_tag <= _GEN_6391;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_247_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_247_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_247_target_address <= _GEN_11495;
      end
    end else begin
      btb_247_target_address <= _GEN_11495;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_247_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_247_bht <= 2'h1;
        end else begin
          btb_247_bht <= 2'h0;
        end
      end else begin
        btb_247_bht <= _GEN_11497;
      end
    end else begin
      btb_247_bht <= _GEN_11497;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_248_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_248_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_248_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_248_valid <= _GEN_15610;
      end
    end else begin
      btb_248_valid <= _GEN_15610;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_248_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_248_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_248_tag <= _GEN_6392;
      end
    end else begin
      btb_248_tag <= _GEN_6392;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_248_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_248_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_248_target_address <= _GEN_11498;
      end
    end else begin
      btb_248_target_address <= _GEN_11498;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_248_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_248_bht <= 2'h1;
        end else begin
          btb_248_bht <= 2'h0;
        end
      end else begin
        btb_248_bht <= _GEN_11500;
      end
    end else begin
      btb_248_bht <= _GEN_11500;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_249_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_249_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_249_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_249_valid <= _GEN_15611;
      end
    end else begin
      btb_249_valid <= _GEN_15611;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_249_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_249_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_249_tag <= _GEN_6393;
      end
    end else begin
      btb_249_tag <= _GEN_6393;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_249_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_249_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_249_target_address <= _GEN_11501;
      end
    end else begin
      btb_249_target_address <= _GEN_11501;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_249_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hf9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_249_bht <= 2'h1;
        end else begin
          btb_249_bht <= 2'h0;
        end
      end else begin
        btb_249_bht <= _GEN_11503;
      end
    end else begin
      btb_249_bht <= _GEN_11503;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_250_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_250_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_250_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_250_valid <= _GEN_15612;
      end
    end else begin
      btb_250_valid <= _GEN_15612;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_250_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfa == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_250_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_250_tag <= _GEN_6394;
      end
    end else begin
      btb_250_tag <= _GEN_6394;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_250_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfa == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_250_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_250_target_address <= _GEN_11504;
      end
    end else begin
      btb_250_target_address <= _GEN_11504;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_250_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfa == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_250_bht <= 2'h1;
        end else begin
          btb_250_bht <= 2'h0;
        end
      end else begin
        btb_250_bht <= _GEN_11506;
      end
    end else begin
      btb_250_bht <= _GEN_11506;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_251_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_251_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_251_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_251_valid <= _GEN_15613;
      end
    end else begin
      btb_251_valid <= _GEN_15613;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_251_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_251_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_251_tag <= _GEN_6395;
      end
    end else begin
      btb_251_tag <= _GEN_6395;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_251_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_251_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_251_target_address <= _GEN_11507;
      end
    end else begin
      btb_251_target_address <= _GEN_11507;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_251_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_251_bht <= 2'h1;
        end else begin
          btb_251_bht <= 2'h0;
        end
      end else begin
        btb_251_bht <= _GEN_11509;
      end
    end else begin
      btb_251_bht <= _GEN_11509;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_252_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_252_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_252_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_252_valid <= _GEN_15614;
      end
    end else begin
      btb_252_valid <= _GEN_15614;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_252_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_252_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_252_tag <= _GEN_6396;
      end
    end else begin
      btb_252_tag <= _GEN_6396;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_252_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_252_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_252_target_address <= _GEN_11510;
      end
    end else begin
      btb_252_target_address <= _GEN_11510;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_252_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_252_bht <= 2'h1;
        end else begin
          btb_252_bht <= 2'h0;
        end
      end else begin
        btb_252_bht <= _GEN_11512;
      end
    end else begin
      btb_252_bht <= _GEN_11512;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_253_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_253_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_253_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_253_valid <= _GEN_15615;
      end
    end else begin
      btb_253_valid <= _GEN_15615;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_253_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_253_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_253_tag <= _GEN_6397;
      end
    end else begin
      btb_253_tag <= _GEN_6397;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_253_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_253_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_253_target_address <= _GEN_11513;
      end
    end else begin
      btb_253_target_address <= _GEN_11513;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_253_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_253_bht <= 2'h1;
        end else begin
          btb_253_bht <= 2'h0;
        end
      end else begin
        btb_253_bht <= _GEN_11515;
      end
    end else begin
      btb_253_bht <= _GEN_11515;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_254_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_254_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_254_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_254_valid <= _GEN_15616;
      end
    end else begin
      btb_254_valid <= _GEN_15616;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_254_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfe == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_254_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_254_tag <= _GEN_6398;
      end
    end else begin
      btb_254_tag <= _GEN_6398;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_254_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfe == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_254_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_254_target_address <= _GEN_11516;
      end
    end else begin
      btb_254_target_address <= _GEN_11516;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_254_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hfe == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_254_bht <= 2'h1;
        end else begin
          btb_254_bht <= 2'h0;
        end
      end else begin
        btb_254_bht <= _GEN_11518;
      end
    end else begin
      btb_254_bht <= _GEN_11518;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_255_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_255_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_255_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_255_valid <= _GEN_15617;
      end
    end else begin
      btb_255_valid <= _GEN_15617;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_255_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hff == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_255_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_255_tag <= _GEN_6399;
      end
    end else begin
      btb_255_tag <= _GEN_6399;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_255_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hff == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_255_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_255_target_address <= _GEN_11519;
      end
    end else begin
      btb_255_target_address <= _GEN_11519;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_255_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'hff == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_255_bht <= 2'h1;
        end else begin
          btb_255_bht <= 2'h0;
        end
      end else begin
        btb_255_bht <= _GEN_11521;
      end
    end else begin
      btb_255_bht <= _GEN_11521;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_256_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_256_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_256_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_256_valid <= _GEN_15618;
      end
    end else begin
      btb_256_valid <= _GEN_15618;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_256_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h100 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_256_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_256_tag <= _GEN_6400;
      end
    end else begin
      btb_256_tag <= _GEN_6400;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_256_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h100 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_256_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_256_target_address <= _GEN_11522;
      end
    end else begin
      btb_256_target_address <= _GEN_11522;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_256_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h100 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_256_bht <= 2'h1;
        end else begin
          btb_256_bht <= 2'h0;
        end
      end else begin
        btb_256_bht <= _GEN_11524;
      end
    end else begin
      btb_256_bht <= _GEN_11524;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_257_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_257_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_257_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_257_valid <= _GEN_15619;
      end
    end else begin
      btb_257_valid <= _GEN_15619;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_257_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h101 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_257_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_257_tag <= _GEN_6401;
      end
    end else begin
      btb_257_tag <= _GEN_6401;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_257_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h101 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_257_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_257_target_address <= _GEN_11525;
      end
    end else begin
      btb_257_target_address <= _GEN_11525;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_257_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h101 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_257_bht <= 2'h1;
        end else begin
          btb_257_bht <= 2'h0;
        end
      end else begin
        btb_257_bht <= _GEN_11527;
      end
    end else begin
      btb_257_bht <= _GEN_11527;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_258_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_258_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_258_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_258_valid <= _GEN_15620;
      end
    end else begin
      btb_258_valid <= _GEN_15620;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_258_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h102 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_258_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_258_tag <= _GEN_6402;
      end
    end else begin
      btb_258_tag <= _GEN_6402;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_258_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h102 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_258_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_258_target_address <= _GEN_11528;
      end
    end else begin
      btb_258_target_address <= _GEN_11528;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_258_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h102 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_258_bht <= 2'h1;
        end else begin
          btb_258_bht <= 2'h0;
        end
      end else begin
        btb_258_bht <= _GEN_11530;
      end
    end else begin
      btb_258_bht <= _GEN_11530;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_259_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_259_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_259_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_259_valid <= _GEN_15621;
      end
    end else begin
      btb_259_valid <= _GEN_15621;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_259_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h103 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_259_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_259_tag <= _GEN_6403;
      end
    end else begin
      btb_259_tag <= _GEN_6403;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_259_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h103 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_259_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_259_target_address <= _GEN_11531;
      end
    end else begin
      btb_259_target_address <= _GEN_11531;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_259_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h103 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_259_bht <= 2'h1;
        end else begin
          btb_259_bht <= 2'h0;
        end
      end else begin
        btb_259_bht <= _GEN_11533;
      end
    end else begin
      btb_259_bht <= _GEN_11533;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_260_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_260_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_260_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_260_valid <= _GEN_15622;
      end
    end else begin
      btb_260_valid <= _GEN_15622;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_260_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h104 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_260_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_260_tag <= _GEN_6404;
      end
    end else begin
      btb_260_tag <= _GEN_6404;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_260_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h104 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_260_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_260_target_address <= _GEN_11534;
      end
    end else begin
      btb_260_target_address <= _GEN_11534;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_260_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h104 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_260_bht <= 2'h1;
        end else begin
          btb_260_bht <= 2'h0;
        end
      end else begin
        btb_260_bht <= _GEN_11536;
      end
    end else begin
      btb_260_bht <= _GEN_11536;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_261_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_261_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_261_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_261_valid <= _GEN_15623;
      end
    end else begin
      btb_261_valid <= _GEN_15623;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_261_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h105 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_261_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_261_tag <= _GEN_6405;
      end
    end else begin
      btb_261_tag <= _GEN_6405;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_261_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h105 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_261_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_261_target_address <= _GEN_11537;
      end
    end else begin
      btb_261_target_address <= _GEN_11537;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_261_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h105 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_261_bht <= 2'h1;
        end else begin
          btb_261_bht <= 2'h0;
        end
      end else begin
        btb_261_bht <= _GEN_11539;
      end
    end else begin
      btb_261_bht <= _GEN_11539;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_262_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_262_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_262_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_262_valid <= _GEN_15624;
      end
    end else begin
      btb_262_valid <= _GEN_15624;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_262_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h106 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_262_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_262_tag <= _GEN_6406;
      end
    end else begin
      btb_262_tag <= _GEN_6406;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_262_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h106 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_262_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_262_target_address <= _GEN_11540;
      end
    end else begin
      btb_262_target_address <= _GEN_11540;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_262_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h106 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_262_bht <= 2'h1;
        end else begin
          btb_262_bht <= 2'h0;
        end
      end else begin
        btb_262_bht <= _GEN_11542;
      end
    end else begin
      btb_262_bht <= _GEN_11542;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_263_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_263_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_263_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_263_valid <= _GEN_15625;
      end
    end else begin
      btb_263_valid <= _GEN_15625;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_263_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h107 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_263_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_263_tag <= _GEN_6407;
      end
    end else begin
      btb_263_tag <= _GEN_6407;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_263_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h107 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_263_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_263_target_address <= _GEN_11543;
      end
    end else begin
      btb_263_target_address <= _GEN_11543;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_263_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h107 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_263_bht <= 2'h1;
        end else begin
          btb_263_bht <= 2'h0;
        end
      end else begin
        btb_263_bht <= _GEN_11545;
      end
    end else begin
      btb_263_bht <= _GEN_11545;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_264_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_264_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_264_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_264_valid <= _GEN_15626;
      end
    end else begin
      btb_264_valid <= _GEN_15626;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_264_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h108 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_264_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_264_tag <= _GEN_6408;
      end
    end else begin
      btb_264_tag <= _GEN_6408;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_264_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h108 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_264_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_264_target_address <= _GEN_11546;
      end
    end else begin
      btb_264_target_address <= _GEN_11546;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_264_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h108 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_264_bht <= 2'h1;
        end else begin
          btb_264_bht <= 2'h0;
        end
      end else begin
        btb_264_bht <= _GEN_11548;
      end
    end else begin
      btb_264_bht <= _GEN_11548;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_265_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_265_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_265_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_265_valid <= _GEN_15627;
      end
    end else begin
      btb_265_valid <= _GEN_15627;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_265_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h109 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_265_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_265_tag <= _GEN_6409;
      end
    end else begin
      btb_265_tag <= _GEN_6409;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_265_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h109 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_265_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_265_target_address <= _GEN_11549;
      end
    end else begin
      btb_265_target_address <= _GEN_11549;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_265_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h109 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_265_bht <= 2'h1;
        end else begin
          btb_265_bht <= 2'h0;
        end
      end else begin
        btb_265_bht <= _GEN_11551;
      end
    end else begin
      btb_265_bht <= _GEN_11551;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_266_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_266_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_266_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_266_valid <= _GEN_15628;
      end
    end else begin
      btb_266_valid <= _GEN_15628;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_266_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_266_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_266_tag <= _GEN_6410;
      end
    end else begin
      btb_266_tag <= _GEN_6410;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_266_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_266_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_266_target_address <= _GEN_11552;
      end
    end else begin
      btb_266_target_address <= _GEN_11552;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_266_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_266_bht <= 2'h1;
        end else begin
          btb_266_bht <= 2'h0;
        end
      end else begin
        btb_266_bht <= _GEN_11554;
      end
    end else begin
      btb_266_bht <= _GEN_11554;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_267_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_267_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_267_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_267_valid <= _GEN_15629;
      end
    end else begin
      btb_267_valid <= _GEN_15629;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_267_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_267_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_267_tag <= _GEN_6411;
      end
    end else begin
      btb_267_tag <= _GEN_6411;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_267_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_267_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_267_target_address <= _GEN_11555;
      end
    end else begin
      btb_267_target_address <= _GEN_11555;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_267_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_267_bht <= 2'h1;
        end else begin
          btb_267_bht <= 2'h0;
        end
      end else begin
        btb_267_bht <= _GEN_11557;
      end
    end else begin
      btb_267_bht <= _GEN_11557;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_268_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_268_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_268_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_268_valid <= _GEN_15630;
      end
    end else begin
      btb_268_valid <= _GEN_15630;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_268_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_268_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_268_tag <= _GEN_6412;
      end
    end else begin
      btb_268_tag <= _GEN_6412;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_268_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_268_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_268_target_address <= _GEN_11558;
      end
    end else begin
      btb_268_target_address <= _GEN_11558;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_268_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_268_bht <= 2'h1;
        end else begin
          btb_268_bht <= 2'h0;
        end
      end else begin
        btb_268_bht <= _GEN_11560;
      end
    end else begin
      btb_268_bht <= _GEN_11560;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_269_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_269_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_269_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_269_valid <= _GEN_15631;
      end
    end else begin
      btb_269_valid <= _GEN_15631;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_269_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_269_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_269_tag <= _GEN_6413;
      end
    end else begin
      btb_269_tag <= _GEN_6413;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_269_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_269_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_269_target_address <= _GEN_11561;
      end
    end else begin
      btb_269_target_address <= _GEN_11561;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_269_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_269_bht <= 2'h1;
        end else begin
          btb_269_bht <= 2'h0;
        end
      end else begin
        btb_269_bht <= _GEN_11563;
      end
    end else begin
      btb_269_bht <= _GEN_11563;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_270_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_270_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_270_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_270_valid <= _GEN_15632;
      end
    end else begin
      btb_270_valid <= _GEN_15632;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_270_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_270_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_270_tag <= _GEN_6414;
      end
    end else begin
      btb_270_tag <= _GEN_6414;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_270_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_270_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_270_target_address <= _GEN_11564;
      end
    end else begin
      btb_270_target_address <= _GEN_11564;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_270_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_270_bht <= 2'h1;
        end else begin
          btb_270_bht <= 2'h0;
        end
      end else begin
        btb_270_bht <= _GEN_11566;
      end
    end else begin
      btb_270_bht <= _GEN_11566;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_271_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_271_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_271_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_271_valid <= _GEN_15633;
      end
    end else begin
      btb_271_valid <= _GEN_15633;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_271_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_271_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_271_tag <= _GEN_6415;
      end
    end else begin
      btb_271_tag <= _GEN_6415;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_271_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_271_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_271_target_address <= _GEN_11567;
      end
    end else begin
      btb_271_target_address <= _GEN_11567;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_271_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h10f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_271_bht <= 2'h1;
        end else begin
          btb_271_bht <= 2'h0;
        end
      end else begin
        btb_271_bht <= _GEN_11569;
      end
    end else begin
      btb_271_bht <= _GEN_11569;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_272_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_272_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_272_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_272_valid <= _GEN_15634;
      end
    end else begin
      btb_272_valid <= _GEN_15634;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_272_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h110 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_272_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_272_tag <= _GEN_6416;
      end
    end else begin
      btb_272_tag <= _GEN_6416;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_272_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h110 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_272_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_272_target_address <= _GEN_11570;
      end
    end else begin
      btb_272_target_address <= _GEN_11570;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_272_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h110 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_272_bht <= 2'h1;
        end else begin
          btb_272_bht <= 2'h0;
        end
      end else begin
        btb_272_bht <= _GEN_11572;
      end
    end else begin
      btb_272_bht <= _GEN_11572;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_273_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_273_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_273_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_273_valid <= _GEN_15635;
      end
    end else begin
      btb_273_valid <= _GEN_15635;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_273_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h111 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_273_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_273_tag <= _GEN_6417;
      end
    end else begin
      btb_273_tag <= _GEN_6417;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_273_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h111 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_273_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_273_target_address <= _GEN_11573;
      end
    end else begin
      btb_273_target_address <= _GEN_11573;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_273_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h111 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_273_bht <= 2'h1;
        end else begin
          btb_273_bht <= 2'h0;
        end
      end else begin
        btb_273_bht <= _GEN_11575;
      end
    end else begin
      btb_273_bht <= _GEN_11575;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_274_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_274_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_274_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_274_valid <= _GEN_15636;
      end
    end else begin
      btb_274_valid <= _GEN_15636;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_274_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h112 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_274_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_274_tag <= _GEN_6418;
      end
    end else begin
      btb_274_tag <= _GEN_6418;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_274_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h112 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_274_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_274_target_address <= _GEN_11576;
      end
    end else begin
      btb_274_target_address <= _GEN_11576;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_274_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h112 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_274_bht <= 2'h1;
        end else begin
          btb_274_bht <= 2'h0;
        end
      end else begin
        btb_274_bht <= _GEN_11578;
      end
    end else begin
      btb_274_bht <= _GEN_11578;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_275_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_275_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_275_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_275_valid <= _GEN_15637;
      end
    end else begin
      btb_275_valid <= _GEN_15637;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_275_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h113 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_275_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_275_tag <= _GEN_6419;
      end
    end else begin
      btb_275_tag <= _GEN_6419;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_275_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h113 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_275_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_275_target_address <= _GEN_11579;
      end
    end else begin
      btb_275_target_address <= _GEN_11579;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_275_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h113 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_275_bht <= 2'h1;
        end else begin
          btb_275_bht <= 2'h0;
        end
      end else begin
        btb_275_bht <= _GEN_11581;
      end
    end else begin
      btb_275_bht <= _GEN_11581;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_276_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_276_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_276_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_276_valid <= _GEN_15638;
      end
    end else begin
      btb_276_valid <= _GEN_15638;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_276_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h114 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_276_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_276_tag <= _GEN_6420;
      end
    end else begin
      btb_276_tag <= _GEN_6420;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_276_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h114 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_276_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_276_target_address <= _GEN_11582;
      end
    end else begin
      btb_276_target_address <= _GEN_11582;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_276_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h114 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_276_bht <= 2'h1;
        end else begin
          btb_276_bht <= 2'h0;
        end
      end else begin
        btb_276_bht <= _GEN_11584;
      end
    end else begin
      btb_276_bht <= _GEN_11584;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_277_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_277_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_277_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_277_valid <= _GEN_15639;
      end
    end else begin
      btb_277_valid <= _GEN_15639;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_277_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h115 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_277_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_277_tag <= _GEN_6421;
      end
    end else begin
      btb_277_tag <= _GEN_6421;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_277_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h115 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_277_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_277_target_address <= _GEN_11585;
      end
    end else begin
      btb_277_target_address <= _GEN_11585;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_277_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h115 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_277_bht <= 2'h1;
        end else begin
          btb_277_bht <= 2'h0;
        end
      end else begin
        btb_277_bht <= _GEN_11587;
      end
    end else begin
      btb_277_bht <= _GEN_11587;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_278_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_278_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_278_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_278_valid <= _GEN_15640;
      end
    end else begin
      btb_278_valid <= _GEN_15640;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_278_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h116 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_278_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_278_tag <= _GEN_6422;
      end
    end else begin
      btb_278_tag <= _GEN_6422;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_278_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h116 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_278_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_278_target_address <= _GEN_11588;
      end
    end else begin
      btb_278_target_address <= _GEN_11588;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_278_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h116 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_278_bht <= 2'h1;
        end else begin
          btb_278_bht <= 2'h0;
        end
      end else begin
        btb_278_bht <= _GEN_11590;
      end
    end else begin
      btb_278_bht <= _GEN_11590;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_279_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_279_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_279_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_279_valid <= _GEN_15641;
      end
    end else begin
      btb_279_valid <= _GEN_15641;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_279_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h117 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_279_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_279_tag <= _GEN_6423;
      end
    end else begin
      btb_279_tag <= _GEN_6423;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_279_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h117 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_279_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_279_target_address <= _GEN_11591;
      end
    end else begin
      btb_279_target_address <= _GEN_11591;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_279_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h117 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_279_bht <= 2'h1;
        end else begin
          btb_279_bht <= 2'h0;
        end
      end else begin
        btb_279_bht <= _GEN_11593;
      end
    end else begin
      btb_279_bht <= _GEN_11593;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_280_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_280_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_280_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_280_valid <= _GEN_15642;
      end
    end else begin
      btb_280_valid <= _GEN_15642;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_280_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h118 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_280_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_280_tag <= _GEN_6424;
      end
    end else begin
      btb_280_tag <= _GEN_6424;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_280_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h118 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_280_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_280_target_address <= _GEN_11594;
      end
    end else begin
      btb_280_target_address <= _GEN_11594;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_280_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h118 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_280_bht <= 2'h1;
        end else begin
          btb_280_bht <= 2'h0;
        end
      end else begin
        btb_280_bht <= _GEN_11596;
      end
    end else begin
      btb_280_bht <= _GEN_11596;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_281_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_281_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_281_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_281_valid <= _GEN_15643;
      end
    end else begin
      btb_281_valid <= _GEN_15643;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_281_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h119 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_281_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_281_tag <= _GEN_6425;
      end
    end else begin
      btb_281_tag <= _GEN_6425;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_281_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h119 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_281_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_281_target_address <= _GEN_11597;
      end
    end else begin
      btb_281_target_address <= _GEN_11597;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_281_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h119 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_281_bht <= 2'h1;
        end else begin
          btb_281_bht <= 2'h0;
        end
      end else begin
        btb_281_bht <= _GEN_11599;
      end
    end else begin
      btb_281_bht <= _GEN_11599;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_282_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_282_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_282_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_282_valid <= _GEN_15644;
      end
    end else begin
      btb_282_valid <= _GEN_15644;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_282_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_282_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_282_tag <= _GEN_6426;
      end
    end else begin
      btb_282_tag <= _GEN_6426;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_282_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_282_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_282_target_address <= _GEN_11600;
      end
    end else begin
      btb_282_target_address <= _GEN_11600;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_282_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_282_bht <= 2'h1;
        end else begin
          btb_282_bht <= 2'h0;
        end
      end else begin
        btb_282_bht <= _GEN_11602;
      end
    end else begin
      btb_282_bht <= _GEN_11602;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_283_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_283_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_283_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_283_valid <= _GEN_15645;
      end
    end else begin
      btb_283_valid <= _GEN_15645;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_283_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_283_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_283_tag <= _GEN_6427;
      end
    end else begin
      btb_283_tag <= _GEN_6427;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_283_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_283_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_283_target_address <= _GEN_11603;
      end
    end else begin
      btb_283_target_address <= _GEN_11603;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_283_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_283_bht <= 2'h1;
        end else begin
          btb_283_bht <= 2'h0;
        end
      end else begin
        btb_283_bht <= _GEN_11605;
      end
    end else begin
      btb_283_bht <= _GEN_11605;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_284_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_284_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_284_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_284_valid <= _GEN_15646;
      end
    end else begin
      btb_284_valid <= _GEN_15646;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_284_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_284_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_284_tag <= _GEN_6428;
      end
    end else begin
      btb_284_tag <= _GEN_6428;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_284_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_284_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_284_target_address <= _GEN_11606;
      end
    end else begin
      btb_284_target_address <= _GEN_11606;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_284_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_284_bht <= 2'h1;
        end else begin
          btb_284_bht <= 2'h0;
        end
      end else begin
        btb_284_bht <= _GEN_11608;
      end
    end else begin
      btb_284_bht <= _GEN_11608;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_285_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_285_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_285_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_285_valid <= _GEN_15647;
      end
    end else begin
      btb_285_valid <= _GEN_15647;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_285_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_285_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_285_tag <= _GEN_6429;
      end
    end else begin
      btb_285_tag <= _GEN_6429;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_285_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_285_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_285_target_address <= _GEN_11609;
      end
    end else begin
      btb_285_target_address <= _GEN_11609;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_285_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_285_bht <= 2'h1;
        end else begin
          btb_285_bht <= 2'h0;
        end
      end else begin
        btb_285_bht <= _GEN_11611;
      end
    end else begin
      btb_285_bht <= _GEN_11611;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_286_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_286_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_286_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_286_valid <= _GEN_15648;
      end
    end else begin
      btb_286_valid <= _GEN_15648;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_286_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_286_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_286_tag <= _GEN_6430;
      end
    end else begin
      btb_286_tag <= _GEN_6430;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_286_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_286_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_286_target_address <= _GEN_11612;
      end
    end else begin
      btb_286_target_address <= _GEN_11612;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_286_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_286_bht <= 2'h1;
        end else begin
          btb_286_bht <= 2'h0;
        end
      end else begin
        btb_286_bht <= _GEN_11614;
      end
    end else begin
      btb_286_bht <= _GEN_11614;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_287_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_287_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_287_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_287_valid <= _GEN_15649;
      end
    end else begin
      btb_287_valid <= _GEN_15649;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_287_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_287_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_287_tag <= _GEN_6431;
      end
    end else begin
      btb_287_tag <= _GEN_6431;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_287_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_287_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_287_target_address <= _GEN_11615;
      end
    end else begin
      btb_287_target_address <= _GEN_11615;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_287_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h11f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_287_bht <= 2'h1;
        end else begin
          btb_287_bht <= 2'h0;
        end
      end else begin
        btb_287_bht <= _GEN_11617;
      end
    end else begin
      btb_287_bht <= _GEN_11617;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_288_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_288_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_288_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_288_valid <= _GEN_15650;
      end
    end else begin
      btb_288_valid <= _GEN_15650;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_288_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h120 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_288_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_288_tag <= _GEN_6432;
      end
    end else begin
      btb_288_tag <= _GEN_6432;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_288_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h120 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_288_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_288_target_address <= _GEN_11618;
      end
    end else begin
      btb_288_target_address <= _GEN_11618;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_288_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h120 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_288_bht <= 2'h1;
        end else begin
          btb_288_bht <= 2'h0;
        end
      end else begin
        btb_288_bht <= _GEN_11620;
      end
    end else begin
      btb_288_bht <= _GEN_11620;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_289_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_289_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_289_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_289_valid <= _GEN_15651;
      end
    end else begin
      btb_289_valid <= _GEN_15651;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_289_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h121 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_289_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_289_tag <= _GEN_6433;
      end
    end else begin
      btb_289_tag <= _GEN_6433;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_289_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h121 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_289_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_289_target_address <= _GEN_11621;
      end
    end else begin
      btb_289_target_address <= _GEN_11621;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_289_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h121 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_289_bht <= 2'h1;
        end else begin
          btb_289_bht <= 2'h0;
        end
      end else begin
        btb_289_bht <= _GEN_11623;
      end
    end else begin
      btb_289_bht <= _GEN_11623;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_290_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_290_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_290_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_290_valid <= _GEN_15652;
      end
    end else begin
      btb_290_valid <= _GEN_15652;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_290_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h122 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_290_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_290_tag <= _GEN_6434;
      end
    end else begin
      btb_290_tag <= _GEN_6434;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_290_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h122 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_290_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_290_target_address <= _GEN_11624;
      end
    end else begin
      btb_290_target_address <= _GEN_11624;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_290_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h122 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_290_bht <= 2'h1;
        end else begin
          btb_290_bht <= 2'h0;
        end
      end else begin
        btb_290_bht <= _GEN_11626;
      end
    end else begin
      btb_290_bht <= _GEN_11626;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_291_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_291_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_291_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_291_valid <= _GEN_15653;
      end
    end else begin
      btb_291_valid <= _GEN_15653;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_291_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h123 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_291_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_291_tag <= _GEN_6435;
      end
    end else begin
      btb_291_tag <= _GEN_6435;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_291_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h123 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_291_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_291_target_address <= _GEN_11627;
      end
    end else begin
      btb_291_target_address <= _GEN_11627;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_291_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h123 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_291_bht <= 2'h1;
        end else begin
          btb_291_bht <= 2'h0;
        end
      end else begin
        btb_291_bht <= _GEN_11629;
      end
    end else begin
      btb_291_bht <= _GEN_11629;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_292_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_292_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_292_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_292_valid <= _GEN_15654;
      end
    end else begin
      btb_292_valid <= _GEN_15654;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_292_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h124 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_292_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_292_tag <= _GEN_6436;
      end
    end else begin
      btb_292_tag <= _GEN_6436;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_292_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h124 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_292_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_292_target_address <= _GEN_11630;
      end
    end else begin
      btb_292_target_address <= _GEN_11630;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_292_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h124 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_292_bht <= 2'h1;
        end else begin
          btb_292_bht <= 2'h0;
        end
      end else begin
        btb_292_bht <= _GEN_11632;
      end
    end else begin
      btb_292_bht <= _GEN_11632;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_293_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_293_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_293_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_293_valid <= _GEN_15655;
      end
    end else begin
      btb_293_valid <= _GEN_15655;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_293_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h125 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_293_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_293_tag <= _GEN_6437;
      end
    end else begin
      btb_293_tag <= _GEN_6437;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_293_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h125 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_293_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_293_target_address <= _GEN_11633;
      end
    end else begin
      btb_293_target_address <= _GEN_11633;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_293_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h125 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_293_bht <= 2'h1;
        end else begin
          btb_293_bht <= 2'h0;
        end
      end else begin
        btb_293_bht <= _GEN_11635;
      end
    end else begin
      btb_293_bht <= _GEN_11635;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_294_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_294_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_294_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_294_valid <= _GEN_15656;
      end
    end else begin
      btb_294_valid <= _GEN_15656;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_294_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h126 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_294_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_294_tag <= _GEN_6438;
      end
    end else begin
      btb_294_tag <= _GEN_6438;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_294_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h126 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_294_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_294_target_address <= _GEN_11636;
      end
    end else begin
      btb_294_target_address <= _GEN_11636;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_294_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h126 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_294_bht <= 2'h1;
        end else begin
          btb_294_bht <= 2'h0;
        end
      end else begin
        btb_294_bht <= _GEN_11638;
      end
    end else begin
      btb_294_bht <= _GEN_11638;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_295_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_295_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_295_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_295_valid <= _GEN_15657;
      end
    end else begin
      btb_295_valid <= _GEN_15657;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_295_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h127 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_295_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_295_tag <= _GEN_6439;
      end
    end else begin
      btb_295_tag <= _GEN_6439;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_295_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h127 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_295_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_295_target_address <= _GEN_11639;
      end
    end else begin
      btb_295_target_address <= _GEN_11639;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_295_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h127 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_295_bht <= 2'h1;
        end else begin
          btb_295_bht <= 2'h0;
        end
      end else begin
        btb_295_bht <= _GEN_11641;
      end
    end else begin
      btb_295_bht <= _GEN_11641;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_296_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_296_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_296_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_296_valid <= _GEN_15658;
      end
    end else begin
      btb_296_valid <= _GEN_15658;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_296_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h128 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_296_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_296_tag <= _GEN_6440;
      end
    end else begin
      btb_296_tag <= _GEN_6440;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_296_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h128 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_296_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_296_target_address <= _GEN_11642;
      end
    end else begin
      btb_296_target_address <= _GEN_11642;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_296_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h128 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_296_bht <= 2'h1;
        end else begin
          btb_296_bht <= 2'h0;
        end
      end else begin
        btb_296_bht <= _GEN_11644;
      end
    end else begin
      btb_296_bht <= _GEN_11644;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_297_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_297_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_297_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_297_valid <= _GEN_15659;
      end
    end else begin
      btb_297_valid <= _GEN_15659;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_297_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h129 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_297_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_297_tag <= _GEN_6441;
      end
    end else begin
      btb_297_tag <= _GEN_6441;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_297_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h129 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_297_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_297_target_address <= _GEN_11645;
      end
    end else begin
      btb_297_target_address <= _GEN_11645;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_297_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h129 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_297_bht <= 2'h1;
        end else begin
          btb_297_bht <= 2'h0;
        end
      end else begin
        btb_297_bht <= _GEN_11647;
      end
    end else begin
      btb_297_bht <= _GEN_11647;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_298_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_298_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_298_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_298_valid <= _GEN_15660;
      end
    end else begin
      btb_298_valid <= _GEN_15660;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_298_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_298_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_298_tag <= _GEN_6442;
      end
    end else begin
      btb_298_tag <= _GEN_6442;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_298_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_298_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_298_target_address <= _GEN_11648;
      end
    end else begin
      btb_298_target_address <= _GEN_11648;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_298_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_298_bht <= 2'h1;
        end else begin
          btb_298_bht <= 2'h0;
        end
      end else begin
        btb_298_bht <= _GEN_11650;
      end
    end else begin
      btb_298_bht <= _GEN_11650;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_299_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_299_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_299_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_299_valid <= _GEN_15661;
      end
    end else begin
      btb_299_valid <= _GEN_15661;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_299_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_299_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_299_tag <= _GEN_6443;
      end
    end else begin
      btb_299_tag <= _GEN_6443;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_299_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_299_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_299_target_address <= _GEN_11651;
      end
    end else begin
      btb_299_target_address <= _GEN_11651;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_299_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_299_bht <= 2'h1;
        end else begin
          btb_299_bht <= 2'h0;
        end
      end else begin
        btb_299_bht <= _GEN_11653;
      end
    end else begin
      btb_299_bht <= _GEN_11653;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_300_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_300_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_300_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_300_valid <= _GEN_15662;
      end
    end else begin
      btb_300_valid <= _GEN_15662;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_300_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_300_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_300_tag <= _GEN_6444;
      end
    end else begin
      btb_300_tag <= _GEN_6444;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_300_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_300_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_300_target_address <= _GEN_11654;
      end
    end else begin
      btb_300_target_address <= _GEN_11654;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_300_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_300_bht <= 2'h1;
        end else begin
          btb_300_bht <= 2'h0;
        end
      end else begin
        btb_300_bht <= _GEN_11656;
      end
    end else begin
      btb_300_bht <= _GEN_11656;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_301_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_301_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_301_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_301_valid <= _GEN_15663;
      end
    end else begin
      btb_301_valid <= _GEN_15663;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_301_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_301_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_301_tag <= _GEN_6445;
      end
    end else begin
      btb_301_tag <= _GEN_6445;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_301_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_301_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_301_target_address <= _GEN_11657;
      end
    end else begin
      btb_301_target_address <= _GEN_11657;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_301_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_301_bht <= 2'h1;
        end else begin
          btb_301_bht <= 2'h0;
        end
      end else begin
        btb_301_bht <= _GEN_11659;
      end
    end else begin
      btb_301_bht <= _GEN_11659;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_302_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_302_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_302_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_302_valid <= _GEN_15664;
      end
    end else begin
      btb_302_valid <= _GEN_15664;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_302_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_302_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_302_tag <= _GEN_6446;
      end
    end else begin
      btb_302_tag <= _GEN_6446;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_302_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_302_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_302_target_address <= _GEN_11660;
      end
    end else begin
      btb_302_target_address <= _GEN_11660;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_302_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_302_bht <= 2'h1;
        end else begin
          btb_302_bht <= 2'h0;
        end
      end else begin
        btb_302_bht <= _GEN_11662;
      end
    end else begin
      btb_302_bht <= _GEN_11662;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_303_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_303_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_303_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_303_valid <= _GEN_15665;
      end
    end else begin
      btb_303_valid <= _GEN_15665;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_303_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_303_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_303_tag <= _GEN_6447;
      end
    end else begin
      btb_303_tag <= _GEN_6447;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_303_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_303_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_303_target_address <= _GEN_11663;
      end
    end else begin
      btb_303_target_address <= _GEN_11663;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_303_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h12f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_303_bht <= 2'h1;
        end else begin
          btb_303_bht <= 2'h0;
        end
      end else begin
        btb_303_bht <= _GEN_11665;
      end
    end else begin
      btb_303_bht <= _GEN_11665;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_304_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_304_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_304_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_304_valid <= _GEN_15666;
      end
    end else begin
      btb_304_valid <= _GEN_15666;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_304_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h130 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_304_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_304_tag <= _GEN_6448;
      end
    end else begin
      btb_304_tag <= _GEN_6448;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_304_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h130 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_304_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_304_target_address <= _GEN_11666;
      end
    end else begin
      btb_304_target_address <= _GEN_11666;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_304_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h130 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_304_bht <= 2'h1;
        end else begin
          btb_304_bht <= 2'h0;
        end
      end else begin
        btb_304_bht <= _GEN_11668;
      end
    end else begin
      btb_304_bht <= _GEN_11668;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_305_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_305_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_305_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_305_valid <= _GEN_15667;
      end
    end else begin
      btb_305_valid <= _GEN_15667;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_305_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h131 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_305_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_305_tag <= _GEN_6449;
      end
    end else begin
      btb_305_tag <= _GEN_6449;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_305_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h131 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_305_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_305_target_address <= _GEN_11669;
      end
    end else begin
      btb_305_target_address <= _GEN_11669;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_305_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h131 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_305_bht <= 2'h1;
        end else begin
          btb_305_bht <= 2'h0;
        end
      end else begin
        btb_305_bht <= _GEN_11671;
      end
    end else begin
      btb_305_bht <= _GEN_11671;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_306_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_306_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_306_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_306_valid <= _GEN_15668;
      end
    end else begin
      btb_306_valid <= _GEN_15668;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_306_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h132 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_306_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_306_tag <= _GEN_6450;
      end
    end else begin
      btb_306_tag <= _GEN_6450;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_306_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h132 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_306_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_306_target_address <= _GEN_11672;
      end
    end else begin
      btb_306_target_address <= _GEN_11672;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_306_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h132 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_306_bht <= 2'h1;
        end else begin
          btb_306_bht <= 2'h0;
        end
      end else begin
        btb_306_bht <= _GEN_11674;
      end
    end else begin
      btb_306_bht <= _GEN_11674;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_307_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_307_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_307_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_307_valid <= _GEN_15669;
      end
    end else begin
      btb_307_valid <= _GEN_15669;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_307_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h133 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_307_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_307_tag <= _GEN_6451;
      end
    end else begin
      btb_307_tag <= _GEN_6451;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_307_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h133 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_307_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_307_target_address <= _GEN_11675;
      end
    end else begin
      btb_307_target_address <= _GEN_11675;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_307_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h133 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_307_bht <= 2'h1;
        end else begin
          btb_307_bht <= 2'h0;
        end
      end else begin
        btb_307_bht <= _GEN_11677;
      end
    end else begin
      btb_307_bht <= _GEN_11677;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_308_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_308_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_308_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_308_valid <= _GEN_15670;
      end
    end else begin
      btb_308_valid <= _GEN_15670;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_308_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h134 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_308_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_308_tag <= _GEN_6452;
      end
    end else begin
      btb_308_tag <= _GEN_6452;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_308_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h134 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_308_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_308_target_address <= _GEN_11678;
      end
    end else begin
      btb_308_target_address <= _GEN_11678;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_308_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h134 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_308_bht <= 2'h1;
        end else begin
          btb_308_bht <= 2'h0;
        end
      end else begin
        btb_308_bht <= _GEN_11680;
      end
    end else begin
      btb_308_bht <= _GEN_11680;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_309_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_309_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_309_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_309_valid <= _GEN_15671;
      end
    end else begin
      btb_309_valid <= _GEN_15671;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_309_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h135 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_309_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_309_tag <= _GEN_6453;
      end
    end else begin
      btb_309_tag <= _GEN_6453;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_309_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h135 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_309_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_309_target_address <= _GEN_11681;
      end
    end else begin
      btb_309_target_address <= _GEN_11681;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_309_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h135 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_309_bht <= 2'h1;
        end else begin
          btb_309_bht <= 2'h0;
        end
      end else begin
        btb_309_bht <= _GEN_11683;
      end
    end else begin
      btb_309_bht <= _GEN_11683;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_310_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_310_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_310_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_310_valid <= _GEN_15672;
      end
    end else begin
      btb_310_valid <= _GEN_15672;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_310_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h136 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_310_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_310_tag <= _GEN_6454;
      end
    end else begin
      btb_310_tag <= _GEN_6454;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_310_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h136 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_310_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_310_target_address <= _GEN_11684;
      end
    end else begin
      btb_310_target_address <= _GEN_11684;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_310_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h136 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_310_bht <= 2'h1;
        end else begin
          btb_310_bht <= 2'h0;
        end
      end else begin
        btb_310_bht <= _GEN_11686;
      end
    end else begin
      btb_310_bht <= _GEN_11686;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_311_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_311_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_311_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_311_valid <= _GEN_15673;
      end
    end else begin
      btb_311_valid <= _GEN_15673;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_311_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h137 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_311_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_311_tag <= _GEN_6455;
      end
    end else begin
      btb_311_tag <= _GEN_6455;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_311_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h137 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_311_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_311_target_address <= _GEN_11687;
      end
    end else begin
      btb_311_target_address <= _GEN_11687;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_311_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h137 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_311_bht <= 2'h1;
        end else begin
          btb_311_bht <= 2'h0;
        end
      end else begin
        btb_311_bht <= _GEN_11689;
      end
    end else begin
      btb_311_bht <= _GEN_11689;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_312_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_312_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_312_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_312_valid <= _GEN_15674;
      end
    end else begin
      btb_312_valid <= _GEN_15674;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_312_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h138 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_312_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_312_tag <= _GEN_6456;
      end
    end else begin
      btb_312_tag <= _GEN_6456;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_312_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h138 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_312_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_312_target_address <= _GEN_11690;
      end
    end else begin
      btb_312_target_address <= _GEN_11690;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_312_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h138 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_312_bht <= 2'h1;
        end else begin
          btb_312_bht <= 2'h0;
        end
      end else begin
        btb_312_bht <= _GEN_11692;
      end
    end else begin
      btb_312_bht <= _GEN_11692;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_313_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_313_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_313_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_313_valid <= _GEN_15675;
      end
    end else begin
      btb_313_valid <= _GEN_15675;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_313_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h139 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_313_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_313_tag <= _GEN_6457;
      end
    end else begin
      btb_313_tag <= _GEN_6457;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_313_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h139 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_313_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_313_target_address <= _GEN_11693;
      end
    end else begin
      btb_313_target_address <= _GEN_11693;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_313_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h139 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_313_bht <= 2'h1;
        end else begin
          btb_313_bht <= 2'h0;
        end
      end else begin
        btb_313_bht <= _GEN_11695;
      end
    end else begin
      btb_313_bht <= _GEN_11695;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_314_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_314_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_314_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_314_valid <= _GEN_15676;
      end
    end else begin
      btb_314_valid <= _GEN_15676;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_314_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_314_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_314_tag <= _GEN_6458;
      end
    end else begin
      btb_314_tag <= _GEN_6458;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_314_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_314_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_314_target_address <= _GEN_11696;
      end
    end else begin
      btb_314_target_address <= _GEN_11696;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_314_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_314_bht <= 2'h1;
        end else begin
          btb_314_bht <= 2'h0;
        end
      end else begin
        btb_314_bht <= _GEN_11698;
      end
    end else begin
      btb_314_bht <= _GEN_11698;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_315_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_315_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_315_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_315_valid <= _GEN_15677;
      end
    end else begin
      btb_315_valid <= _GEN_15677;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_315_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_315_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_315_tag <= _GEN_6459;
      end
    end else begin
      btb_315_tag <= _GEN_6459;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_315_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_315_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_315_target_address <= _GEN_11699;
      end
    end else begin
      btb_315_target_address <= _GEN_11699;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_315_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_315_bht <= 2'h1;
        end else begin
          btb_315_bht <= 2'h0;
        end
      end else begin
        btb_315_bht <= _GEN_11701;
      end
    end else begin
      btb_315_bht <= _GEN_11701;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_316_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_316_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_316_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_316_valid <= _GEN_15678;
      end
    end else begin
      btb_316_valid <= _GEN_15678;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_316_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_316_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_316_tag <= _GEN_6460;
      end
    end else begin
      btb_316_tag <= _GEN_6460;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_316_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_316_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_316_target_address <= _GEN_11702;
      end
    end else begin
      btb_316_target_address <= _GEN_11702;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_316_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_316_bht <= 2'h1;
        end else begin
          btb_316_bht <= 2'h0;
        end
      end else begin
        btb_316_bht <= _GEN_11704;
      end
    end else begin
      btb_316_bht <= _GEN_11704;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_317_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_317_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_317_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_317_valid <= _GEN_15679;
      end
    end else begin
      btb_317_valid <= _GEN_15679;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_317_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_317_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_317_tag <= _GEN_6461;
      end
    end else begin
      btb_317_tag <= _GEN_6461;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_317_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_317_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_317_target_address <= _GEN_11705;
      end
    end else begin
      btb_317_target_address <= _GEN_11705;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_317_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_317_bht <= 2'h1;
        end else begin
          btb_317_bht <= 2'h0;
        end
      end else begin
        btb_317_bht <= _GEN_11707;
      end
    end else begin
      btb_317_bht <= _GEN_11707;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_318_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_318_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_318_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_318_valid <= _GEN_15680;
      end
    end else begin
      btb_318_valid <= _GEN_15680;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_318_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_318_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_318_tag <= _GEN_6462;
      end
    end else begin
      btb_318_tag <= _GEN_6462;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_318_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_318_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_318_target_address <= _GEN_11708;
      end
    end else begin
      btb_318_target_address <= _GEN_11708;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_318_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_318_bht <= 2'h1;
        end else begin
          btb_318_bht <= 2'h0;
        end
      end else begin
        btb_318_bht <= _GEN_11710;
      end
    end else begin
      btb_318_bht <= _GEN_11710;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_319_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_319_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_319_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_319_valid <= _GEN_15681;
      end
    end else begin
      btb_319_valid <= _GEN_15681;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_319_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_319_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_319_tag <= _GEN_6463;
      end
    end else begin
      btb_319_tag <= _GEN_6463;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_319_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_319_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_319_target_address <= _GEN_11711;
      end
    end else begin
      btb_319_target_address <= _GEN_11711;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_319_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h13f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_319_bht <= 2'h1;
        end else begin
          btb_319_bht <= 2'h0;
        end
      end else begin
        btb_319_bht <= _GEN_11713;
      end
    end else begin
      btb_319_bht <= _GEN_11713;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_320_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_320_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_320_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_320_valid <= _GEN_15682;
      end
    end else begin
      btb_320_valid <= _GEN_15682;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_320_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h140 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_320_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_320_tag <= _GEN_6464;
      end
    end else begin
      btb_320_tag <= _GEN_6464;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_320_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h140 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_320_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_320_target_address <= _GEN_11714;
      end
    end else begin
      btb_320_target_address <= _GEN_11714;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_320_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h140 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_320_bht <= 2'h1;
        end else begin
          btb_320_bht <= 2'h0;
        end
      end else begin
        btb_320_bht <= _GEN_11716;
      end
    end else begin
      btb_320_bht <= _GEN_11716;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_321_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_321_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_321_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_321_valid <= _GEN_15683;
      end
    end else begin
      btb_321_valid <= _GEN_15683;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_321_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h141 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_321_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_321_tag <= _GEN_6465;
      end
    end else begin
      btb_321_tag <= _GEN_6465;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_321_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h141 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_321_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_321_target_address <= _GEN_11717;
      end
    end else begin
      btb_321_target_address <= _GEN_11717;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_321_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h141 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_321_bht <= 2'h1;
        end else begin
          btb_321_bht <= 2'h0;
        end
      end else begin
        btb_321_bht <= _GEN_11719;
      end
    end else begin
      btb_321_bht <= _GEN_11719;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_322_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_322_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_322_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_322_valid <= _GEN_15684;
      end
    end else begin
      btb_322_valid <= _GEN_15684;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_322_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h142 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_322_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_322_tag <= _GEN_6466;
      end
    end else begin
      btb_322_tag <= _GEN_6466;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_322_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h142 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_322_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_322_target_address <= _GEN_11720;
      end
    end else begin
      btb_322_target_address <= _GEN_11720;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_322_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h142 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_322_bht <= 2'h1;
        end else begin
          btb_322_bht <= 2'h0;
        end
      end else begin
        btb_322_bht <= _GEN_11722;
      end
    end else begin
      btb_322_bht <= _GEN_11722;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_323_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_323_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_323_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_323_valid <= _GEN_15685;
      end
    end else begin
      btb_323_valid <= _GEN_15685;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_323_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h143 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_323_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_323_tag <= _GEN_6467;
      end
    end else begin
      btb_323_tag <= _GEN_6467;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_323_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h143 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_323_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_323_target_address <= _GEN_11723;
      end
    end else begin
      btb_323_target_address <= _GEN_11723;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_323_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h143 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_323_bht <= 2'h1;
        end else begin
          btb_323_bht <= 2'h0;
        end
      end else begin
        btb_323_bht <= _GEN_11725;
      end
    end else begin
      btb_323_bht <= _GEN_11725;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_324_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_324_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_324_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_324_valid <= _GEN_15686;
      end
    end else begin
      btb_324_valid <= _GEN_15686;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_324_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h144 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_324_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_324_tag <= _GEN_6468;
      end
    end else begin
      btb_324_tag <= _GEN_6468;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_324_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h144 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_324_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_324_target_address <= _GEN_11726;
      end
    end else begin
      btb_324_target_address <= _GEN_11726;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_324_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h144 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_324_bht <= 2'h1;
        end else begin
          btb_324_bht <= 2'h0;
        end
      end else begin
        btb_324_bht <= _GEN_11728;
      end
    end else begin
      btb_324_bht <= _GEN_11728;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_325_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_325_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_325_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_325_valid <= _GEN_15687;
      end
    end else begin
      btb_325_valid <= _GEN_15687;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_325_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h145 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_325_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_325_tag <= _GEN_6469;
      end
    end else begin
      btb_325_tag <= _GEN_6469;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_325_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h145 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_325_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_325_target_address <= _GEN_11729;
      end
    end else begin
      btb_325_target_address <= _GEN_11729;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_325_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h145 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_325_bht <= 2'h1;
        end else begin
          btb_325_bht <= 2'h0;
        end
      end else begin
        btb_325_bht <= _GEN_11731;
      end
    end else begin
      btb_325_bht <= _GEN_11731;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_326_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_326_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_326_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_326_valid <= _GEN_15688;
      end
    end else begin
      btb_326_valid <= _GEN_15688;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_326_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h146 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_326_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_326_tag <= _GEN_6470;
      end
    end else begin
      btb_326_tag <= _GEN_6470;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_326_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h146 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_326_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_326_target_address <= _GEN_11732;
      end
    end else begin
      btb_326_target_address <= _GEN_11732;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_326_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h146 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_326_bht <= 2'h1;
        end else begin
          btb_326_bht <= 2'h0;
        end
      end else begin
        btb_326_bht <= _GEN_11734;
      end
    end else begin
      btb_326_bht <= _GEN_11734;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_327_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_327_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_327_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_327_valid <= _GEN_15689;
      end
    end else begin
      btb_327_valid <= _GEN_15689;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_327_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h147 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_327_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_327_tag <= _GEN_6471;
      end
    end else begin
      btb_327_tag <= _GEN_6471;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_327_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h147 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_327_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_327_target_address <= _GEN_11735;
      end
    end else begin
      btb_327_target_address <= _GEN_11735;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_327_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h147 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_327_bht <= 2'h1;
        end else begin
          btb_327_bht <= 2'h0;
        end
      end else begin
        btb_327_bht <= _GEN_11737;
      end
    end else begin
      btb_327_bht <= _GEN_11737;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_328_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_328_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_328_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_328_valid <= _GEN_15690;
      end
    end else begin
      btb_328_valid <= _GEN_15690;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_328_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h148 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_328_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_328_tag <= _GEN_6472;
      end
    end else begin
      btb_328_tag <= _GEN_6472;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_328_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h148 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_328_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_328_target_address <= _GEN_11738;
      end
    end else begin
      btb_328_target_address <= _GEN_11738;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_328_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h148 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_328_bht <= 2'h1;
        end else begin
          btb_328_bht <= 2'h0;
        end
      end else begin
        btb_328_bht <= _GEN_11740;
      end
    end else begin
      btb_328_bht <= _GEN_11740;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_329_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_329_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_329_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_329_valid <= _GEN_15691;
      end
    end else begin
      btb_329_valid <= _GEN_15691;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_329_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h149 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_329_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_329_tag <= _GEN_6473;
      end
    end else begin
      btb_329_tag <= _GEN_6473;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_329_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h149 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_329_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_329_target_address <= _GEN_11741;
      end
    end else begin
      btb_329_target_address <= _GEN_11741;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_329_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h149 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_329_bht <= 2'h1;
        end else begin
          btb_329_bht <= 2'h0;
        end
      end else begin
        btb_329_bht <= _GEN_11743;
      end
    end else begin
      btb_329_bht <= _GEN_11743;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_330_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_330_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_330_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_330_valid <= _GEN_15692;
      end
    end else begin
      btb_330_valid <= _GEN_15692;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_330_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_330_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_330_tag <= _GEN_6474;
      end
    end else begin
      btb_330_tag <= _GEN_6474;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_330_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_330_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_330_target_address <= _GEN_11744;
      end
    end else begin
      btb_330_target_address <= _GEN_11744;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_330_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_330_bht <= 2'h1;
        end else begin
          btb_330_bht <= 2'h0;
        end
      end else begin
        btb_330_bht <= _GEN_11746;
      end
    end else begin
      btb_330_bht <= _GEN_11746;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_331_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_331_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_331_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_331_valid <= _GEN_15693;
      end
    end else begin
      btb_331_valid <= _GEN_15693;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_331_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_331_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_331_tag <= _GEN_6475;
      end
    end else begin
      btb_331_tag <= _GEN_6475;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_331_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_331_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_331_target_address <= _GEN_11747;
      end
    end else begin
      btb_331_target_address <= _GEN_11747;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_331_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_331_bht <= 2'h1;
        end else begin
          btb_331_bht <= 2'h0;
        end
      end else begin
        btb_331_bht <= _GEN_11749;
      end
    end else begin
      btb_331_bht <= _GEN_11749;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_332_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_332_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_332_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_332_valid <= _GEN_15694;
      end
    end else begin
      btb_332_valid <= _GEN_15694;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_332_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_332_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_332_tag <= _GEN_6476;
      end
    end else begin
      btb_332_tag <= _GEN_6476;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_332_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_332_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_332_target_address <= _GEN_11750;
      end
    end else begin
      btb_332_target_address <= _GEN_11750;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_332_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_332_bht <= 2'h1;
        end else begin
          btb_332_bht <= 2'h0;
        end
      end else begin
        btb_332_bht <= _GEN_11752;
      end
    end else begin
      btb_332_bht <= _GEN_11752;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_333_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_333_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_333_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_333_valid <= _GEN_15695;
      end
    end else begin
      btb_333_valid <= _GEN_15695;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_333_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_333_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_333_tag <= _GEN_6477;
      end
    end else begin
      btb_333_tag <= _GEN_6477;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_333_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_333_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_333_target_address <= _GEN_11753;
      end
    end else begin
      btb_333_target_address <= _GEN_11753;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_333_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_333_bht <= 2'h1;
        end else begin
          btb_333_bht <= 2'h0;
        end
      end else begin
        btb_333_bht <= _GEN_11755;
      end
    end else begin
      btb_333_bht <= _GEN_11755;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_334_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_334_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_334_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_334_valid <= _GEN_15696;
      end
    end else begin
      btb_334_valid <= _GEN_15696;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_334_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_334_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_334_tag <= _GEN_6478;
      end
    end else begin
      btb_334_tag <= _GEN_6478;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_334_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_334_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_334_target_address <= _GEN_11756;
      end
    end else begin
      btb_334_target_address <= _GEN_11756;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_334_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_334_bht <= 2'h1;
        end else begin
          btb_334_bht <= 2'h0;
        end
      end else begin
        btb_334_bht <= _GEN_11758;
      end
    end else begin
      btb_334_bht <= _GEN_11758;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_335_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_335_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_335_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_335_valid <= _GEN_15697;
      end
    end else begin
      btb_335_valid <= _GEN_15697;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_335_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_335_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_335_tag <= _GEN_6479;
      end
    end else begin
      btb_335_tag <= _GEN_6479;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_335_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_335_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_335_target_address <= _GEN_11759;
      end
    end else begin
      btb_335_target_address <= _GEN_11759;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_335_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h14f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_335_bht <= 2'h1;
        end else begin
          btb_335_bht <= 2'h0;
        end
      end else begin
        btb_335_bht <= _GEN_11761;
      end
    end else begin
      btb_335_bht <= _GEN_11761;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_336_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_336_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_336_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_336_valid <= _GEN_15698;
      end
    end else begin
      btb_336_valid <= _GEN_15698;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_336_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h150 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_336_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_336_tag <= _GEN_6480;
      end
    end else begin
      btb_336_tag <= _GEN_6480;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_336_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h150 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_336_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_336_target_address <= _GEN_11762;
      end
    end else begin
      btb_336_target_address <= _GEN_11762;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_336_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h150 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_336_bht <= 2'h1;
        end else begin
          btb_336_bht <= 2'h0;
        end
      end else begin
        btb_336_bht <= _GEN_11764;
      end
    end else begin
      btb_336_bht <= _GEN_11764;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_337_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_337_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_337_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_337_valid <= _GEN_15699;
      end
    end else begin
      btb_337_valid <= _GEN_15699;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_337_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h151 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_337_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_337_tag <= _GEN_6481;
      end
    end else begin
      btb_337_tag <= _GEN_6481;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_337_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h151 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_337_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_337_target_address <= _GEN_11765;
      end
    end else begin
      btb_337_target_address <= _GEN_11765;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_337_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h151 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_337_bht <= 2'h1;
        end else begin
          btb_337_bht <= 2'h0;
        end
      end else begin
        btb_337_bht <= _GEN_11767;
      end
    end else begin
      btb_337_bht <= _GEN_11767;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_338_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_338_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_338_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_338_valid <= _GEN_15700;
      end
    end else begin
      btb_338_valid <= _GEN_15700;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_338_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h152 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_338_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_338_tag <= _GEN_6482;
      end
    end else begin
      btb_338_tag <= _GEN_6482;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_338_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h152 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_338_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_338_target_address <= _GEN_11768;
      end
    end else begin
      btb_338_target_address <= _GEN_11768;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_338_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h152 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_338_bht <= 2'h1;
        end else begin
          btb_338_bht <= 2'h0;
        end
      end else begin
        btb_338_bht <= _GEN_11770;
      end
    end else begin
      btb_338_bht <= _GEN_11770;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_339_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_339_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_339_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_339_valid <= _GEN_15701;
      end
    end else begin
      btb_339_valid <= _GEN_15701;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_339_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h153 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_339_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_339_tag <= _GEN_6483;
      end
    end else begin
      btb_339_tag <= _GEN_6483;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_339_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h153 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_339_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_339_target_address <= _GEN_11771;
      end
    end else begin
      btb_339_target_address <= _GEN_11771;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_339_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h153 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_339_bht <= 2'h1;
        end else begin
          btb_339_bht <= 2'h0;
        end
      end else begin
        btb_339_bht <= _GEN_11773;
      end
    end else begin
      btb_339_bht <= _GEN_11773;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_340_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_340_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_340_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_340_valid <= _GEN_15702;
      end
    end else begin
      btb_340_valid <= _GEN_15702;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_340_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h154 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_340_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_340_tag <= _GEN_6484;
      end
    end else begin
      btb_340_tag <= _GEN_6484;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_340_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h154 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_340_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_340_target_address <= _GEN_11774;
      end
    end else begin
      btb_340_target_address <= _GEN_11774;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_340_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h154 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_340_bht <= 2'h1;
        end else begin
          btb_340_bht <= 2'h0;
        end
      end else begin
        btb_340_bht <= _GEN_11776;
      end
    end else begin
      btb_340_bht <= _GEN_11776;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_341_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_341_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_341_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_341_valid <= _GEN_15703;
      end
    end else begin
      btb_341_valid <= _GEN_15703;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_341_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h155 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_341_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_341_tag <= _GEN_6485;
      end
    end else begin
      btb_341_tag <= _GEN_6485;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_341_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h155 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_341_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_341_target_address <= _GEN_11777;
      end
    end else begin
      btb_341_target_address <= _GEN_11777;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_341_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h155 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_341_bht <= 2'h1;
        end else begin
          btb_341_bht <= 2'h0;
        end
      end else begin
        btb_341_bht <= _GEN_11779;
      end
    end else begin
      btb_341_bht <= _GEN_11779;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_342_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_342_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_342_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_342_valid <= _GEN_15704;
      end
    end else begin
      btb_342_valid <= _GEN_15704;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_342_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h156 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_342_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_342_tag <= _GEN_6486;
      end
    end else begin
      btb_342_tag <= _GEN_6486;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_342_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h156 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_342_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_342_target_address <= _GEN_11780;
      end
    end else begin
      btb_342_target_address <= _GEN_11780;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_342_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h156 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_342_bht <= 2'h1;
        end else begin
          btb_342_bht <= 2'h0;
        end
      end else begin
        btb_342_bht <= _GEN_11782;
      end
    end else begin
      btb_342_bht <= _GEN_11782;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_343_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_343_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_343_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_343_valid <= _GEN_15705;
      end
    end else begin
      btb_343_valid <= _GEN_15705;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_343_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h157 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_343_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_343_tag <= _GEN_6487;
      end
    end else begin
      btb_343_tag <= _GEN_6487;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_343_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h157 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_343_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_343_target_address <= _GEN_11783;
      end
    end else begin
      btb_343_target_address <= _GEN_11783;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_343_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h157 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_343_bht <= 2'h1;
        end else begin
          btb_343_bht <= 2'h0;
        end
      end else begin
        btb_343_bht <= _GEN_11785;
      end
    end else begin
      btb_343_bht <= _GEN_11785;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_344_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_344_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_344_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_344_valid <= _GEN_15706;
      end
    end else begin
      btb_344_valid <= _GEN_15706;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_344_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h158 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_344_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_344_tag <= _GEN_6488;
      end
    end else begin
      btb_344_tag <= _GEN_6488;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_344_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h158 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_344_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_344_target_address <= _GEN_11786;
      end
    end else begin
      btb_344_target_address <= _GEN_11786;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_344_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h158 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_344_bht <= 2'h1;
        end else begin
          btb_344_bht <= 2'h0;
        end
      end else begin
        btb_344_bht <= _GEN_11788;
      end
    end else begin
      btb_344_bht <= _GEN_11788;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_345_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_345_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_345_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_345_valid <= _GEN_15707;
      end
    end else begin
      btb_345_valid <= _GEN_15707;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_345_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h159 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_345_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_345_tag <= _GEN_6489;
      end
    end else begin
      btb_345_tag <= _GEN_6489;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_345_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h159 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_345_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_345_target_address <= _GEN_11789;
      end
    end else begin
      btb_345_target_address <= _GEN_11789;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_345_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h159 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_345_bht <= 2'h1;
        end else begin
          btb_345_bht <= 2'h0;
        end
      end else begin
        btb_345_bht <= _GEN_11791;
      end
    end else begin
      btb_345_bht <= _GEN_11791;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_346_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_346_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_346_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_346_valid <= _GEN_15708;
      end
    end else begin
      btb_346_valid <= _GEN_15708;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_346_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_346_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_346_tag <= _GEN_6490;
      end
    end else begin
      btb_346_tag <= _GEN_6490;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_346_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_346_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_346_target_address <= _GEN_11792;
      end
    end else begin
      btb_346_target_address <= _GEN_11792;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_346_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_346_bht <= 2'h1;
        end else begin
          btb_346_bht <= 2'h0;
        end
      end else begin
        btb_346_bht <= _GEN_11794;
      end
    end else begin
      btb_346_bht <= _GEN_11794;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_347_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_347_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_347_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_347_valid <= _GEN_15709;
      end
    end else begin
      btb_347_valid <= _GEN_15709;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_347_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_347_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_347_tag <= _GEN_6491;
      end
    end else begin
      btb_347_tag <= _GEN_6491;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_347_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_347_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_347_target_address <= _GEN_11795;
      end
    end else begin
      btb_347_target_address <= _GEN_11795;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_347_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_347_bht <= 2'h1;
        end else begin
          btb_347_bht <= 2'h0;
        end
      end else begin
        btb_347_bht <= _GEN_11797;
      end
    end else begin
      btb_347_bht <= _GEN_11797;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_348_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_348_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_348_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_348_valid <= _GEN_15710;
      end
    end else begin
      btb_348_valid <= _GEN_15710;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_348_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_348_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_348_tag <= _GEN_6492;
      end
    end else begin
      btb_348_tag <= _GEN_6492;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_348_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_348_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_348_target_address <= _GEN_11798;
      end
    end else begin
      btb_348_target_address <= _GEN_11798;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_348_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_348_bht <= 2'h1;
        end else begin
          btb_348_bht <= 2'h0;
        end
      end else begin
        btb_348_bht <= _GEN_11800;
      end
    end else begin
      btb_348_bht <= _GEN_11800;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_349_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_349_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_349_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_349_valid <= _GEN_15711;
      end
    end else begin
      btb_349_valid <= _GEN_15711;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_349_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_349_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_349_tag <= _GEN_6493;
      end
    end else begin
      btb_349_tag <= _GEN_6493;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_349_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_349_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_349_target_address <= _GEN_11801;
      end
    end else begin
      btb_349_target_address <= _GEN_11801;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_349_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_349_bht <= 2'h1;
        end else begin
          btb_349_bht <= 2'h0;
        end
      end else begin
        btb_349_bht <= _GEN_11803;
      end
    end else begin
      btb_349_bht <= _GEN_11803;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_350_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_350_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_350_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_350_valid <= _GEN_15712;
      end
    end else begin
      btb_350_valid <= _GEN_15712;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_350_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_350_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_350_tag <= _GEN_6494;
      end
    end else begin
      btb_350_tag <= _GEN_6494;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_350_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_350_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_350_target_address <= _GEN_11804;
      end
    end else begin
      btb_350_target_address <= _GEN_11804;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_350_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_350_bht <= 2'h1;
        end else begin
          btb_350_bht <= 2'h0;
        end
      end else begin
        btb_350_bht <= _GEN_11806;
      end
    end else begin
      btb_350_bht <= _GEN_11806;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_351_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_351_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_351_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_351_valid <= _GEN_15713;
      end
    end else begin
      btb_351_valid <= _GEN_15713;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_351_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_351_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_351_tag <= _GEN_6495;
      end
    end else begin
      btb_351_tag <= _GEN_6495;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_351_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_351_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_351_target_address <= _GEN_11807;
      end
    end else begin
      btb_351_target_address <= _GEN_11807;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_351_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h15f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_351_bht <= 2'h1;
        end else begin
          btb_351_bht <= 2'h0;
        end
      end else begin
        btb_351_bht <= _GEN_11809;
      end
    end else begin
      btb_351_bht <= _GEN_11809;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_352_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_352_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_352_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_352_valid <= _GEN_15714;
      end
    end else begin
      btb_352_valid <= _GEN_15714;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_352_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h160 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_352_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_352_tag <= _GEN_6496;
      end
    end else begin
      btb_352_tag <= _GEN_6496;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_352_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h160 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_352_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_352_target_address <= _GEN_11810;
      end
    end else begin
      btb_352_target_address <= _GEN_11810;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_352_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h160 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_352_bht <= 2'h1;
        end else begin
          btb_352_bht <= 2'h0;
        end
      end else begin
        btb_352_bht <= _GEN_11812;
      end
    end else begin
      btb_352_bht <= _GEN_11812;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_353_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_353_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_353_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_353_valid <= _GEN_15715;
      end
    end else begin
      btb_353_valid <= _GEN_15715;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_353_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h161 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_353_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_353_tag <= _GEN_6497;
      end
    end else begin
      btb_353_tag <= _GEN_6497;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_353_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h161 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_353_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_353_target_address <= _GEN_11813;
      end
    end else begin
      btb_353_target_address <= _GEN_11813;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_353_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h161 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_353_bht <= 2'h1;
        end else begin
          btb_353_bht <= 2'h0;
        end
      end else begin
        btb_353_bht <= _GEN_11815;
      end
    end else begin
      btb_353_bht <= _GEN_11815;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_354_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_354_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_354_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_354_valid <= _GEN_15716;
      end
    end else begin
      btb_354_valid <= _GEN_15716;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_354_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h162 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_354_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_354_tag <= _GEN_6498;
      end
    end else begin
      btb_354_tag <= _GEN_6498;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_354_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h162 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_354_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_354_target_address <= _GEN_11816;
      end
    end else begin
      btb_354_target_address <= _GEN_11816;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_354_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h162 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_354_bht <= 2'h1;
        end else begin
          btb_354_bht <= 2'h0;
        end
      end else begin
        btb_354_bht <= _GEN_11818;
      end
    end else begin
      btb_354_bht <= _GEN_11818;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_355_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_355_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_355_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_355_valid <= _GEN_15717;
      end
    end else begin
      btb_355_valid <= _GEN_15717;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_355_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h163 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_355_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_355_tag <= _GEN_6499;
      end
    end else begin
      btb_355_tag <= _GEN_6499;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_355_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h163 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_355_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_355_target_address <= _GEN_11819;
      end
    end else begin
      btb_355_target_address <= _GEN_11819;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_355_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h163 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_355_bht <= 2'h1;
        end else begin
          btb_355_bht <= 2'h0;
        end
      end else begin
        btb_355_bht <= _GEN_11821;
      end
    end else begin
      btb_355_bht <= _GEN_11821;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_356_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_356_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_356_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_356_valid <= _GEN_15718;
      end
    end else begin
      btb_356_valid <= _GEN_15718;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_356_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h164 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_356_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_356_tag <= _GEN_6500;
      end
    end else begin
      btb_356_tag <= _GEN_6500;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_356_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h164 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_356_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_356_target_address <= _GEN_11822;
      end
    end else begin
      btb_356_target_address <= _GEN_11822;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_356_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h164 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_356_bht <= 2'h1;
        end else begin
          btb_356_bht <= 2'h0;
        end
      end else begin
        btb_356_bht <= _GEN_11824;
      end
    end else begin
      btb_356_bht <= _GEN_11824;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_357_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_357_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_357_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_357_valid <= _GEN_15719;
      end
    end else begin
      btb_357_valid <= _GEN_15719;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_357_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h165 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_357_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_357_tag <= _GEN_6501;
      end
    end else begin
      btb_357_tag <= _GEN_6501;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_357_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h165 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_357_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_357_target_address <= _GEN_11825;
      end
    end else begin
      btb_357_target_address <= _GEN_11825;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_357_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h165 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_357_bht <= 2'h1;
        end else begin
          btb_357_bht <= 2'h0;
        end
      end else begin
        btb_357_bht <= _GEN_11827;
      end
    end else begin
      btb_357_bht <= _GEN_11827;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_358_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_358_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_358_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_358_valid <= _GEN_15720;
      end
    end else begin
      btb_358_valid <= _GEN_15720;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_358_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h166 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_358_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_358_tag <= _GEN_6502;
      end
    end else begin
      btb_358_tag <= _GEN_6502;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_358_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h166 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_358_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_358_target_address <= _GEN_11828;
      end
    end else begin
      btb_358_target_address <= _GEN_11828;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_358_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h166 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_358_bht <= 2'h1;
        end else begin
          btb_358_bht <= 2'h0;
        end
      end else begin
        btb_358_bht <= _GEN_11830;
      end
    end else begin
      btb_358_bht <= _GEN_11830;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_359_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_359_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_359_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_359_valid <= _GEN_15721;
      end
    end else begin
      btb_359_valid <= _GEN_15721;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_359_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h167 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_359_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_359_tag <= _GEN_6503;
      end
    end else begin
      btb_359_tag <= _GEN_6503;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_359_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h167 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_359_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_359_target_address <= _GEN_11831;
      end
    end else begin
      btb_359_target_address <= _GEN_11831;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_359_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h167 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_359_bht <= 2'h1;
        end else begin
          btb_359_bht <= 2'h0;
        end
      end else begin
        btb_359_bht <= _GEN_11833;
      end
    end else begin
      btb_359_bht <= _GEN_11833;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_360_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_360_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_360_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_360_valid <= _GEN_15722;
      end
    end else begin
      btb_360_valid <= _GEN_15722;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_360_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h168 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_360_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_360_tag <= _GEN_6504;
      end
    end else begin
      btb_360_tag <= _GEN_6504;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_360_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h168 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_360_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_360_target_address <= _GEN_11834;
      end
    end else begin
      btb_360_target_address <= _GEN_11834;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_360_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h168 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_360_bht <= 2'h1;
        end else begin
          btb_360_bht <= 2'h0;
        end
      end else begin
        btb_360_bht <= _GEN_11836;
      end
    end else begin
      btb_360_bht <= _GEN_11836;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_361_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_361_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_361_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_361_valid <= _GEN_15723;
      end
    end else begin
      btb_361_valid <= _GEN_15723;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_361_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h169 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_361_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_361_tag <= _GEN_6505;
      end
    end else begin
      btb_361_tag <= _GEN_6505;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_361_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h169 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_361_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_361_target_address <= _GEN_11837;
      end
    end else begin
      btb_361_target_address <= _GEN_11837;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_361_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h169 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_361_bht <= 2'h1;
        end else begin
          btb_361_bht <= 2'h0;
        end
      end else begin
        btb_361_bht <= _GEN_11839;
      end
    end else begin
      btb_361_bht <= _GEN_11839;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_362_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_362_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_362_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_362_valid <= _GEN_15724;
      end
    end else begin
      btb_362_valid <= _GEN_15724;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_362_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_362_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_362_tag <= _GEN_6506;
      end
    end else begin
      btb_362_tag <= _GEN_6506;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_362_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_362_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_362_target_address <= _GEN_11840;
      end
    end else begin
      btb_362_target_address <= _GEN_11840;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_362_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_362_bht <= 2'h1;
        end else begin
          btb_362_bht <= 2'h0;
        end
      end else begin
        btb_362_bht <= _GEN_11842;
      end
    end else begin
      btb_362_bht <= _GEN_11842;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_363_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_363_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_363_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_363_valid <= _GEN_15725;
      end
    end else begin
      btb_363_valid <= _GEN_15725;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_363_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_363_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_363_tag <= _GEN_6507;
      end
    end else begin
      btb_363_tag <= _GEN_6507;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_363_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_363_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_363_target_address <= _GEN_11843;
      end
    end else begin
      btb_363_target_address <= _GEN_11843;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_363_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_363_bht <= 2'h1;
        end else begin
          btb_363_bht <= 2'h0;
        end
      end else begin
        btb_363_bht <= _GEN_11845;
      end
    end else begin
      btb_363_bht <= _GEN_11845;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_364_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_364_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_364_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_364_valid <= _GEN_15726;
      end
    end else begin
      btb_364_valid <= _GEN_15726;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_364_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_364_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_364_tag <= _GEN_6508;
      end
    end else begin
      btb_364_tag <= _GEN_6508;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_364_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_364_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_364_target_address <= _GEN_11846;
      end
    end else begin
      btb_364_target_address <= _GEN_11846;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_364_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_364_bht <= 2'h1;
        end else begin
          btb_364_bht <= 2'h0;
        end
      end else begin
        btb_364_bht <= _GEN_11848;
      end
    end else begin
      btb_364_bht <= _GEN_11848;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_365_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_365_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_365_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_365_valid <= _GEN_15727;
      end
    end else begin
      btb_365_valid <= _GEN_15727;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_365_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_365_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_365_tag <= _GEN_6509;
      end
    end else begin
      btb_365_tag <= _GEN_6509;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_365_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_365_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_365_target_address <= _GEN_11849;
      end
    end else begin
      btb_365_target_address <= _GEN_11849;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_365_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_365_bht <= 2'h1;
        end else begin
          btb_365_bht <= 2'h0;
        end
      end else begin
        btb_365_bht <= _GEN_11851;
      end
    end else begin
      btb_365_bht <= _GEN_11851;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_366_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_366_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_366_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_366_valid <= _GEN_15728;
      end
    end else begin
      btb_366_valid <= _GEN_15728;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_366_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_366_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_366_tag <= _GEN_6510;
      end
    end else begin
      btb_366_tag <= _GEN_6510;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_366_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_366_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_366_target_address <= _GEN_11852;
      end
    end else begin
      btb_366_target_address <= _GEN_11852;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_366_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_366_bht <= 2'h1;
        end else begin
          btb_366_bht <= 2'h0;
        end
      end else begin
        btb_366_bht <= _GEN_11854;
      end
    end else begin
      btb_366_bht <= _GEN_11854;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_367_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_367_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_367_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_367_valid <= _GEN_15729;
      end
    end else begin
      btb_367_valid <= _GEN_15729;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_367_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_367_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_367_tag <= _GEN_6511;
      end
    end else begin
      btb_367_tag <= _GEN_6511;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_367_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_367_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_367_target_address <= _GEN_11855;
      end
    end else begin
      btb_367_target_address <= _GEN_11855;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_367_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h16f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_367_bht <= 2'h1;
        end else begin
          btb_367_bht <= 2'h0;
        end
      end else begin
        btb_367_bht <= _GEN_11857;
      end
    end else begin
      btb_367_bht <= _GEN_11857;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_368_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_368_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_368_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_368_valid <= _GEN_15730;
      end
    end else begin
      btb_368_valid <= _GEN_15730;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_368_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h170 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_368_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_368_tag <= _GEN_6512;
      end
    end else begin
      btb_368_tag <= _GEN_6512;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_368_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h170 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_368_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_368_target_address <= _GEN_11858;
      end
    end else begin
      btb_368_target_address <= _GEN_11858;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_368_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h170 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_368_bht <= 2'h1;
        end else begin
          btb_368_bht <= 2'h0;
        end
      end else begin
        btb_368_bht <= _GEN_11860;
      end
    end else begin
      btb_368_bht <= _GEN_11860;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_369_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_369_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_369_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_369_valid <= _GEN_15731;
      end
    end else begin
      btb_369_valid <= _GEN_15731;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_369_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h171 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_369_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_369_tag <= _GEN_6513;
      end
    end else begin
      btb_369_tag <= _GEN_6513;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_369_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h171 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_369_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_369_target_address <= _GEN_11861;
      end
    end else begin
      btb_369_target_address <= _GEN_11861;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_369_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h171 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_369_bht <= 2'h1;
        end else begin
          btb_369_bht <= 2'h0;
        end
      end else begin
        btb_369_bht <= _GEN_11863;
      end
    end else begin
      btb_369_bht <= _GEN_11863;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_370_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_370_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_370_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_370_valid <= _GEN_15732;
      end
    end else begin
      btb_370_valid <= _GEN_15732;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_370_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h172 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_370_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_370_tag <= _GEN_6514;
      end
    end else begin
      btb_370_tag <= _GEN_6514;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_370_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h172 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_370_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_370_target_address <= _GEN_11864;
      end
    end else begin
      btb_370_target_address <= _GEN_11864;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_370_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h172 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_370_bht <= 2'h1;
        end else begin
          btb_370_bht <= 2'h0;
        end
      end else begin
        btb_370_bht <= _GEN_11866;
      end
    end else begin
      btb_370_bht <= _GEN_11866;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_371_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_371_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_371_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_371_valid <= _GEN_15733;
      end
    end else begin
      btb_371_valid <= _GEN_15733;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_371_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h173 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_371_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_371_tag <= _GEN_6515;
      end
    end else begin
      btb_371_tag <= _GEN_6515;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_371_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h173 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_371_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_371_target_address <= _GEN_11867;
      end
    end else begin
      btb_371_target_address <= _GEN_11867;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_371_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h173 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_371_bht <= 2'h1;
        end else begin
          btb_371_bht <= 2'h0;
        end
      end else begin
        btb_371_bht <= _GEN_11869;
      end
    end else begin
      btb_371_bht <= _GEN_11869;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_372_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_372_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_372_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_372_valid <= _GEN_15734;
      end
    end else begin
      btb_372_valid <= _GEN_15734;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_372_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h174 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_372_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_372_tag <= _GEN_6516;
      end
    end else begin
      btb_372_tag <= _GEN_6516;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_372_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h174 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_372_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_372_target_address <= _GEN_11870;
      end
    end else begin
      btb_372_target_address <= _GEN_11870;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_372_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h174 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_372_bht <= 2'h1;
        end else begin
          btb_372_bht <= 2'h0;
        end
      end else begin
        btb_372_bht <= _GEN_11872;
      end
    end else begin
      btb_372_bht <= _GEN_11872;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_373_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_373_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_373_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_373_valid <= _GEN_15735;
      end
    end else begin
      btb_373_valid <= _GEN_15735;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_373_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h175 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_373_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_373_tag <= _GEN_6517;
      end
    end else begin
      btb_373_tag <= _GEN_6517;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_373_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h175 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_373_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_373_target_address <= _GEN_11873;
      end
    end else begin
      btb_373_target_address <= _GEN_11873;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_373_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h175 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_373_bht <= 2'h1;
        end else begin
          btb_373_bht <= 2'h0;
        end
      end else begin
        btb_373_bht <= _GEN_11875;
      end
    end else begin
      btb_373_bht <= _GEN_11875;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_374_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_374_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_374_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_374_valid <= _GEN_15736;
      end
    end else begin
      btb_374_valid <= _GEN_15736;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_374_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h176 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_374_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_374_tag <= _GEN_6518;
      end
    end else begin
      btb_374_tag <= _GEN_6518;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_374_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h176 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_374_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_374_target_address <= _GEN_11876;
      end
    end else begin
      btb_374_target_address <= _GEN_11876;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_374_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h176 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_374_bht <= 2'h1;
        end else begin
          btb_374_bht <= 2'h0;
        end
      end else begin
        btb_374_bht <= _GEN_11878;
      end
    end else begin
      btb_374_bht <= _GEN_11878;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_375_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_375_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_375_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_375_valid <= _GEN_15737;
      end
    end else begin
      btb_375_valid <= _GEN_15737;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_375_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h177 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_375_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_375_tag <= _GEN_6519;
      end
    end else begin
      btb_375_tag <= _GEN_6519;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_375_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h177 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_375_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_375_target_address <= _GEN_11879;
      end
    end else begin
      btb_375_target_address <= _GEN_11879;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_375_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h177 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_375_bht <= 2'h1;
        end else begin
          btb_375_bht <= 2'h0;
        end
      end else begin
        btb_375_bht <= _GEN_11881;
      end
    end else begin
      btb_375_bht <= _GEN_11881;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_376_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_376_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_376_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_376_valid <= _GEN_15738;
      end
    end else begin
      btb_376_valid <= _GEN_15738;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_376_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h178 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_376_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_376_tag <= _GEN_6520;
      end
    end else begin
      btb_376_tag <= _GEN_6520;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_376_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h178 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_376_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_376_target_address <= _GEN_11882;
      end
    end else begin
      btb_376_target_address <= _GEN_11882;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_376_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h178 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_376_bht <= 2'h1;
        end else begin
          btb_376_bht <= 2'h0;
        end
      end else begin
        btb_376_bht <= _GEN_11884;
      end
    end else begin
      btb_376_bht <= _GEN_11884;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_377_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_377_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_377_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_377_valid <= _GEN_15739;
      end
    end else begin
      btb_377_valid <= _GEN_15739;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_377_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h179 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_377_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_377_tag <= _GEN_6521;
      end
    end else begin
      btb_377_tag <= _GEN_6521;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_377_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h179 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_377_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_377_target_address <= _GEN_11885;
      end
    end else begin
      btb_377_target_address <= _GEN_11885;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_377_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h179 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_377_bht <= 2'h1;
        end else begin
          btb_377_bht <= 2'h0;
        end
      end else begin
        btb_377_bht <= _GEN_11887;
      end
    end else begin
      btb_377_bht <= _GEN_11887;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_378_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_378_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_378_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_378_valid <= _GEN_15740;
      end
    end else begin
      btb_378_valid <= _GEN_15740;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_378_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_378_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_378_tag <= _GEN_6522;
      end
    end else begin
      btb_378_tag <= _GEN_6522;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_378_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_378_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_378_target_address <= _GEN_11888;
      end
    end else begin
      btb_378_target_address <= _GEN_11888;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_378_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_378_bht <= 2'h1;
        end else begin
          btb_378_bht <= 2'h0;
        end
      end else begin
        btb_378_bht <= _GEN_11890;
      end
    end else begin
      btb_378_bht <= _GEN_11890;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_379_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_379_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_379_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_379_valid <= _GEN_15741;
      end
    end else begin
      btb_379_valid <= _GEN_15741;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_379_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_379_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_379_tag <= _GEN_6523;
      end
    end else begin
      btb_379_tag <= _GEN_6523;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_379_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_379_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_379_target_address <= _GEN_11891;
      end
    end else begin
      btb_379_target_address <= _GEN_11891;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_379_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_379_bht <= 2'h1;
        end else begin
          btb_379_bht <= 2'h0;
        end
      end else begin
        btb_379_bht <= _GEN_11893;
      end
    end else begin
      btb_379_bht <= _GEN_11893;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_380_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_380_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_380_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_380_valid <= _GEN_15742;
      end
    end else begin
      btb_380_valid <= _GEN_15742;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_380_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_380_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_380_tag <= _GEN_6524;
      end
    end else begin
      btb_380_tag <= _GEN_6524;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_380_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_380_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_380_target_address <= _GEN_11894;
      end
    end else begin
      btb_380_target_address <= _GEN_11894;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_380_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_380_bht <= 2'h1;
        end else begin
          btb_380_bht <= 2'h0;
        end
      end else begin
        btb_380_bht <= _GEN_11896;
      end
    end else begin
      btb_380_bht <= _GEN_11896;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_381_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_381_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_381_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_381_valid <= _GEN_15743;
      end
    end else begin
      btb_381_valid <= _GEN_15743;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_381_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_381_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_381_tag <= _GEN_6525;
      end
    end else begin
      btb_381_tag <= _GEN_6525;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_381_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_381_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_381_target_address <= _GEN_11897;
      end
    end else begin
      btb_381_target_address <= _GEN_11897;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_381_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_381_bht <= 2'h1;
        end else begin
          btb_381_bht <= 2'h0;
        end
      end else begin
        btb_381_bht <= _GEN_11899;
      end
    end else begin
      btb_381_bht <= _GEN_11899;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_382_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_382_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_382_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_382_valid <= _GEN_15744;
      end
    end else begin
      btb_382_valid <= _GEN_15744;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_382_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_382_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_382_tag <= _GEN_6526;
      end
    end else begin
      btb_382_tag <= _GEN_6526;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_382_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_382_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_382_target_address <= _GEN_11900;
      end
    end else begin
      btb_382_target_address <= _GEN_11900;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_382_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_382_bht <= 2'h1;
        end else begin
          btb_382_bht <= 2'h0;
        end
      end else begin
        btb_382_bht <= _GEN_11902;
      end
    end else begin
      btb_382_bht <= _GEN_11902;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_383_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_383_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_383_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_383_valid <= _GEN_15745;
      end
    end else begin
      btb_383_valid <= _GEN_15745;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_383_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_383_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_383_tag <= _GEN_6527;
      end
    end else begin
      btb_383_tag <= _GEN_6527;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_383_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_383_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_383_target_address <= _GEN_11903;
      end
    end else begin
      btb_383_target_address <= _GEN_11903;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_383_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h17f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_383_bht <= 2'h1;
        end else begin
          btb_383_bht <= 2'h0;
        end
      end else begin
        btb_383_bht <= _GEN_11905;
      end
    end else begin
      btb_383_bht <= _GEN_11905;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_384_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_384_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_384_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_384_valid <= _GEN_15746;
      end
    end else begin
      btb_384_valid <= _GEN_15746;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_384_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h180 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_384_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_384_tag <= _GEN_6528;
      end
    end else begin
      btb_384_tag <= _GEN_6528;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_384_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h180 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_384_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_384_target_address <= _GEN_11906;
      end
    end else begin
      btb_384_target_address <= _GEN_11906;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_384_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h180 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_384_bht <= 2'h1;
        end else begin
          btb_384_bht <= 2'h0;
        end
      end else begin
        btb_384_bht <= _GEN_11908;
      end
    end else begin
      btb_384_bht <= _GEN_11908;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_385_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_385_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_385_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_385_valid <= _GEN_15747;
      end
    end else begin
      btb_385_valid <= _GEN_15747;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_385_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h181 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_385_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_385_tag <= _GEN_6529;
      end
    end else begin
      btb_385_tag <= _GEN_6529;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_385_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h181 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_385_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_385_target_address <= _GEN_11909;
      end
    end else begin
      btb_385_target_address <= _GEN_11909;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_385_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h181 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_385_bht <= 2'h1;
        end else begin
          btb_385_bht <= 2'h0;
        end
      end else begin
        btb_385_bht <= _GEN_11911;
      end
    end else begin
      btb_385_bht <= _GEN_11911;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_386_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_386_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_386_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_386_valid <= _GEN_15748;
      end
    end else begin
      btb_386_valid <= _GEN_15748;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_386_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h182 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_386_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_386_tag <= _GEN_6530;
      end
    end else begin
      btb_386_tag <= _GEN_6530;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_386_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h182 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_386_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_386_target_address <= _GEN_11912;
      end
    end else begin
      btb_386_target_address <= _GEN_11912;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_386_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h182 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_386_bht <= 2'h1;
        end else begin
          btb_386_bht <= 2'h0;
        end
      end else begin
        btb_386_bht <= _GEN_11914;
      end
    end else begin
      btb_386_bht <= _GEN_11914;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_387_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_387_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_387_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_387_valid <= _GEN_15749;
      end
    end else begin
      btb_387_valid <= _GEN_15749;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_387_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h183 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_387_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_387_tag <= _GEN_6531;
      end
    end else begin
      btb_387_tag <= _GEN_6531;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_387_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h183 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_387_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_387_target_address <= _GEN_11915;
      end
    end else begin
      btb_387_target_address <= _GEN_11915;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_387_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h183 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_387_bht <= 2'h1;
        end else begin
          btb_387_bht <= 2'h0;
        end
      end else begin
        btb_387_bht <= _GEN_11917;
      end
    end else begin
      btb_387_bht <= _GEN_11917;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_388_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_388_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_388_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_388_valid <= _GEN_15750;
      end
    end else begin
      btb_388_valid <= _GEN_15750;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_388_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h184 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_388_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_388_tag <= _GEN_6532;
      end
    end else begin
      btb_388_tag <= _GEN_6532;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_388_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h184 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_388_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_388_target_address <= _GEN_11918;
      end
    end else begin
      btb_388_target_address <= _GEN_11918;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_388_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h184 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_388_bht <= 2'h1;
        end else begin
          btb_388_bht <= 2'h0;
        end
      end else begin
        btb_388_bht <= _GEN_11920;
      end
    end else begin
      btb_388_bht <= _GEN_11920;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_389_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_389_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_389_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_389_valid <= _GEN_15751;
      end
    end else begin
      btb_389_valid <= _GEN_15751;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_389_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h185 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_389_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_389_tag <= _GEN_6533;
      end
    end else begin
      btb_389_tag <= _GEN_6533;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_389_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h185 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_389_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_389_target_address <= _GEN_11921;
      end
    end else begin
      btb_389_target_address <= _GEN_11921;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_389_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h185 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_389_bht <= 2'h1;
        end else begin
          btb_389_bht <= 2'h0;
        end
      end else begin
        btb_389_bht <= _GEN_11923;
      end
    end else begin
      btb_389_bht <= _GEN_11923;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_390_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_390_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_390_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_390_valid <= _GEN_15752;
      end
    end else begin
      btb_390_valid <= _GEN_15752;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_390_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h186 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_390_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_390_tag <= _GEN_6534;
      end
    end else begin
      btb_390_tag <= _GEN_6534;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_390_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h186 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_390_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_390_target_address <= _GEN_11924;
      end
    end else begin
      btb_390_target_address <= _GEN_11924;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_390_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h186 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_390_bht <= 2'h1;
        end else begin
          btb_390_bht <= 2'h0;
        end
      end else begin
        btb_390_bht <= _GEN_11926;
      end
    end else begin
      btb_390_bht <= _GEN_11926;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_391_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_391_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_391_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_391_valid <= _GEN_15753;
      end
    end else begin
      btb_391_valid <= _GEN_15753;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_391_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h187 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_391_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_391_tag <= _GEN_6535;
      end
    end else begin
      btb_391_tag <= _GEN_6535;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_391_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h187 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_391_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_391_target_address <= _GEN_11927;
      end
    end else begin
      btb_391_target_address <= _GEN_11927;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_391_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h187 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_391_bht <= 2'h1;
        end else begin
          btb_391_bht <= 2'h0;
        end
      end else begin
        btb_391_bht <= _GEN_11929;
      end
    end else begin
      btb_391_bht <= _GEN_11929;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_392_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_392_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_392_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_392_valid <= _GEN_15754;
      end
    end else begin
      btb_392_valid <= _GEN_15754;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_392_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h188 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_392_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_392_tag <= _GEN_6536;
      end
    end else begin
      btb_392_tag <= _GEN_6536;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_392_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h188 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_392_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_392_target_address <= _GEN_11930;
      end
    end else begin
      btb_392_target_address <= _GEN_11930;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_392_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h188 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_392_bht <= 2'h1;
        end else begin
          btb_392_bht <= 2'h0;
        end
      end else begin
        btb_392_bht <= _GEN_11932;
      end
    end else begin
      btb_392_bht <= _GEN_11932;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_393_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_393_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_393_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_393_valid <= _GEN_15755;
      end
    end else begin
      btb_393_valid <= _GEN_15755;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_393_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h189 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_393_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_393_tag <= _GEN_6537;
      end
    end else begin
      btb_393_tag <= _GEN_6537;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_393_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h189 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_393_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_393_target_address <= _GEN_11933;
      end
    end else begin
      btb_393_target_address <= _GEN_11933;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_393_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h189 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_393_bht <= 2'h1;
        end else begin
          btb_393_bht <= 2'h0;
        end
      end else begin
        btb_393_bht <= _GEN_11935;
      end
    end else begin
      btb_393_bht <= _GEN_11935;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_394_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_394_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_394_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_394_valid <= _GEN_15756;
      end
    end else begin
      btb_394_valid <= _GEN_15756;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_394_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_394_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_394_tag <= _GEN_6538;
      end
    end else begin
      btb_394_tag <= _GEN_6538;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_394_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_394_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_394_target_address <= _GEN_11936;
      end
    end else begin
      btb_394_target_address <= _GEN_11936;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_394_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_394_bht <= 2'h1;
        end else begin
          btb_394_bht <= 2'h0;
        end
      end else begin
        btb_394_bht <= _GEN_11938;
      end
    end else begin
      btb_394_bht <= _GEN_11938;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_395_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_395_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_395_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_395_valid <= _GEN_15757;
      end
    end else begin
      btb_395_valid <= _GEN_15757;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_395_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_395_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_395_tag <= _GEN_6539;
      end
    end else begin
      btb_395_tag <= _GEN_6539;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_395_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_395_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_395_target_address <= _GEN_11939;
      end
    end else begin
      btb_395_target_address <= _GEN_11939;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_395_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_395_bht <= 2'h1;
        end else begin
          btb_395_bht <= 2'h0;
        end
      end else begin
        btb_395_bht <= _GEN_11941;
      end
    end else begin
      btb_395_bht <= _GEN_11941;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_396_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_396_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_396_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_396_valid <= _GEN_15758;
      end
    end else begin
      btb_396_valid <= _GEN_15758;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_396_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_396_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_396_tag <= _GEN_6540;
      end
    end else begin
      btb_396_tag <= _GEN_6540;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_396_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_396_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_396_target_address <= _GEN_11942;
      end
    end else begin
      btb_396_target_address <= _GEN_11942;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_396_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_396_bht <= 2'h1;
        end else begin
          btb_396_bht <= 2'h0;
        end
      end else begin
        btb_396_bht <= _GEN_11944;
      end
    end else begin
      btb_396_bht <= _GEN_11944;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_397_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_397_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_397_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_397_valid <= _GEN_15759;
      end
    end else begin
      btb_397_valid <= _GEN_15759;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_397_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_397_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_397_tag <= _GEN_6541;
      end
    end else begin
      btb_397_tag <= _GEN_6541;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_397_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_397_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_397_target_address <= _GEN_11945;
      end
    end else begin
      btb_397_target_address <= _GEN_11945;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_397_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_397_bht <= 2'h1;
        end else begin
          btb_397_bht <= 2'h0;
        end
      end else begin
        btb_397_bht <= _GEN_11947;
      end
    end else begin
      btb_397_bht <= _GEN_11947;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_398_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_398_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_398_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_398_valid <= _GEN_15760;
      end
    end else begin
      btb_398_valid <= _GEN_15760;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_398_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_398_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_398_tag <= _GEN_6542;
      end
    end else begin
      btb_398_tag <= _GEN_6542;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_398_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_398_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_398_target_address <= _GEN_11948;
      end
    end else begin
      btb_398_target_address <= _GEN_11948;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_398_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_398_bht <= 2'h1;
        end else begin
          btb_398_bht <= 2'h0;
        end
      end else begin
        btb_398_bht <= _GEN_11950;
      end
    end else begin
      btb_398_bht <= _GEN_11950;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_399_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_399_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_399_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_399_valid <= _GEN_15761;
      end
    end else begin
      btb_399_valid <= _GEN_15761;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_399_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_399_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_399_tag <= _GEN_6543;
      end
    end else begin
      btb_399_tag <= _GEN_6543;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_399_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_399_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_399_target_address <= _GEN_11951;
      end
    end else begin
      btb_399_target_address <= _GEN_11951;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_399_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h18f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_399_bht <= 2'h1;
        end else begin
          btb_399_bht <= 2'h0;
        end
      end else begin
        btb_399_bht <= _GEN_11953;
      end
    end else begin
      btb_399_bht <= _GEN_11953;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_400_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_400_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_400_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_400_valid <= _GEN_15762;
      end
    end else begin
      btb_400_valid <= _GEN_15762;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_400_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h190 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_400_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_400_tag <= _GEN_6544;
      end
    end else begin
      btb_400_tag <= _GEN_6544;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_400_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h190 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_400_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_400_target_address <= _GEN_11954;
      end
    end else begin
      btb_400_target_address <= _GEN_11954;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_400_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h190 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_400_bht <= 2'h1;
        end else begin
          btb_400_bht <= 2'h0;
        end
      end else begin
        btb_400_bht <= _GEN_11956;
      end
    end else begin
      btb_400_bht <= _GEN_11956;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_401_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_401_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_401_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_401_valid <= _GEN_15763;
      end
    end else begin
      btb_401_valid <= _GEN_15763;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_401_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h191 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_401_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_401_tag <= _GEN_6545;
      end
    end else begin
      btb_401_tag <= _GEN_6545;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_401_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h191 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_401_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_401_target_address <= _GEN_11957;
      end
    end else begin
      btb_401_target_address <= _GEN_11957;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_401_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h191 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_401_bht <= 2'h1;
        end else begin
          btb_401_bht <= 2'h0;
        end
      end else begin
        btb_401_bht <= _GEN_11959;
      end
    end else begin
      btb_401_bht <= _GEN_11959;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_402_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_402_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_402_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_402_valid <= _GEN_15764;
      end
    end else begin
      btb_402_valid <= _GEN_15764;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_402_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h192 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_402_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_402_tag <= _GEN_6546;
      end
    end else begin
      btb_402_tag <= _GEN_6546;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_402_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h192 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_402_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_402_target_address <= _GEN_11960;
      end
    end else begin
      btb_402_target_address <= _GEN_11960;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_402_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h192 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_402_bht <= 2'h1;
        end else begin
          btb_402_bht <= 2'h0;
        end
      end else begin
        btb_402_bht <= _GEN_11962;
      end
    end else begin
      btb_402_bht <= _GEN_11962;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_403_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_403_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_403_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_403_valid <= _GEN_15765;
      end
    end else begin
      btb_403_valid <= _GEN_15765;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_403_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h193 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_403_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_403_tag <= _GEN_6547;
      end
    end else begin
      btb_403_tag <= _GEN_6547;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_403_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h193 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_403_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_403_target_address <= _GEN_11963;
      end
    end else begin
      btb_403_target_address <= _GEN_11963;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_403_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h193 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_403_bht <= 2'h1;
        end else begin
          btb_403_bht <= 2'h0;
        end
      end else begin
        btb_403_bht <= _GEN_11965;
      end
    end else begin
      btb_403_bht <= _GEN_11965;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_404_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_404_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_404_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_404_valid <= _GEN_15766;
      end
    end else begin
      btb_404_valid <= _GEN_15766;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_404_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h194 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_404_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_404_tag <= _GEN_6548;
      end
    end else begin
      btb_404_tag <= _GEN_6548;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_404_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h194 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_404_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_404_target_address <= _GEN_11966;
      end
    end else begin
      btb_404_target_address <= _GEN_11966;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_404_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h194 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_404_bht <= 2'h1;
        end else begin
          btb_404_bht <= 2'h0;
        end
      end else begin
        btb_404_bht <= _GEN_11968;
      end
    end else begin
      btb_404_bht <= _GEN_11968;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_405_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_405_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_405_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_405_valid <= _GEN_15767;
      end
    end else begin
      btb_405_valid <= _GEN_15767;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_405_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h195 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_405_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_405_tag <= _GEN_6549;
      end
    end else begin
      btb_405_tag <= _GEN_6549;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_405_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h195 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_405_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_405_target_address <= _GEN_11969;
      end
    end else begin
      btb_405_target_address <= _GEN_11969;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_405_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h195 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_405_bht <= 2'h1;
        end else begin
          btb_405_bht <= 2'h0;
        end
      end else begin
        btb_405_bht <= _GEN_11971;
      end
    end else begin
      btb_405_bht <= _GEN_11971;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_406_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_406_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_406_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_406_valid <= _GEN_15768;
      end
    end else begin
      btb_406_valid <= _GEN_15768;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_406_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h196 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_406_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_406_tag <= _GEN_6550;
      end
    end else begin
      btb_406_tag <= _GEN_6550;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_406_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h196 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_406_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_406_target_address <= _GEN_11972;
      end
    end else begin
      btb_406_target_address <= _GEN_11972;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_406_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h196 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_406_bht <= 2'h1;
        end else begin
          btb_406_bht <= 2'h0;
        end
      end else begin
        btb_406_bht <= _GEN_11974;
      end
    end else begin
      btb_406_bht <= _GEN_11974;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_407_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_407_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_407_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_407_valid <= _GEN_15769;
      end
    end else begin
      btb_407_valid <= _GEN_15769;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_407_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h197 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_407_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_407_tag <= _GEN_6551;
      end
    end else begin
      btb_407_tag <= _GEN_6551;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_407_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h197 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_407_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_407_target_address <= _GEN_11975;
      end
    end else begin
      btb_407_target_address <= _GEN_11975;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_407_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h197 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_407_bht <= 2'h1;
        end else begin
          btb_407_bht <= 2'h0;
        end
      end else begin
        btb_407_bht <= _GEN_11977;
      end
    end else begin
      btb_407_bht <= _GEN_11977;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_408_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_408_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_408_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_408_valid <= _GEN_15770;
      end
    end else begin
      btb_408_valid <= _GEN_15770;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_408_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h198 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_408_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_408_tag <= _GEN_6552;
      end
    end else begin
      btb_408_tag <= _GEN_6552;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_408_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h198 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_408_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_408_target_address <= _GEN_11978;
      end
    end else begin
      btb_408_target_address <= _GEN_11978;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_408_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h198 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_408_bht <= 2'h1;
        end else begin
          btb_408_bht <= 2'h0;
        end
      end else begin
        btb_408_bht <= _GEN_11980;
      end
    end else begin
      btb_408_bht <= _GEN_11980;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_409_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_409_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_409_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_409_valid <= _GEN_15771;
      end
    end else begin
      btb_409_valid <= _GEN_15771;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_409_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h199 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_409_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_409_tag <= _GEN_6553;
      end
    end else begin
      btb_409_tag <= _GEN_6553;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_409_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h199 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_409_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_409_target_address <= _GEN_11981;
      end
    end else begin
      btb_409_target_address <= _GEN_11981;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_409_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h199 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_409_bht <= 2'h1;
        end else begin
          btb_409_bht <= 2'h0;
        end
      end else begin
        btb_409_bht <= _GEN_11983;
      end
    end else begin
      btb_409_bht <= _GEN_11983;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_410_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_410_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_410_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_410_valid <= _GEN_15772;
      end
    end else begin
      btb_410_valid <= _GEN_15772;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_410_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19a == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_410_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_410_tag <= _GEN_6554;
      end
    end else begin
      btb_410_tag <= _GEN_6554;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_410_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19a == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_410_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_410_target_address <= _GEN_11984;
      end
    end else begin
      btb_410_target_address <= _GEN_11984;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_410_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19a == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_410_bht <= 2'h1;
        end else begin
          btb_410_bht <= 2'h0;
        end
      end else begin
        btb_410_bht <= _GEN_11986;
      end
    end else begin
      btb_410_bht <= _GEN_11986;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_411_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_411_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_411_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_411_valid <= _GEN_15773;
      end
    end else begin
      btb_411_valid <= _GEN_15773;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_411_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19b == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_411_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_411_tag <= _GEN_6555;
      end
    end else begin
      btb_411_tag <= _GEN_6555;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_411_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19b == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_411_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_411_target_address <= _GEN_11987;
      end
    end else begin
      btb_411_target_address <= _GEN_11987;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_411_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19b == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_411_bht <= 2'h1;
        end else begin
          btb_411_bht <= 2'h0;
        end
      end else begin
        btb_411_bht <= _GEN_11989;
      end
    end else begin
      btb_411_bht <= _GEN_11989;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_412_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_412_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_412_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_412_valid <= _GEN_15774;
      end
    end else begin
      btb_412_valid <= _GEN_15774;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_412_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19c == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_412_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_412_tag <= _GEN_6556;
      end
    end else begin
      btb_412_tag <= _GEN_6556;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_412_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19c == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_412_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_412_target_address <= _GEN_11990;
      end
    end else begin
      btb_412_target_address <= _GEN_11990;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_412_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19c == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_412_bht <= 2'h1;
        end else begin
          btb_412_bht <= 2'h0;
        end
      end else begin
        btb_412_bht <= _GEN_11992;
      end
    end else begin
      btb_412_bht <= _GEN_11992;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_413_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_413_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_413_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_413_valid <= _GEN_15775;
      end
    end else begin
      btb_413_valid <= _GEN_15775;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_413_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19d == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_413_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_413_tag <= _GEN_6557;
      end
    end else begin
      btb_413_tag <= _GEN_6557;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_413_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19d == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_413_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_413_target_address <= _GEN_11993;
      end
    end else begin
      btb_413_target_address <= _GEN_11993;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_413_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19d == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_413_bht <= 2'h1;
        end else begin
          btb_413_bht <= 2'h0;
        end
      end else begin
        btb_413_bht <= _GEN_11995;
      end
    end else begin
      btb_413_bht <= _GEN_11995;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_414_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_414_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_414_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_414_valid <= _GEN_15776;
      end
    end else begin
      btb_414_valid <= _GEN_15776;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_414_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19e == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_414_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_414_tag <= _GEN_6558;
      end
    end else begin
      btb_414_tag <= _GEN_6558;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_414_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19e == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_414_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_414_target_address <= _GEN_11996;
      end
    end else begin
      btb_414_target_address <= _GEN_11996;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_414_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19e == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_414_bht <= 2'h1;
        end else begin
          btb_414_bht <= 2'h0;
        end
      end else begin
        btb_414_bht <= _GEN_11998;
      end
    end else begin
      btb_414_bht <= _GEN_11998;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_415_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_415_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_415_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_415_valid <= _GEN_15777;
      end
    end else begin
      btb_415_valid <= _GEN_15777;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_415_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19f == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_415_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_415_tag <= _GEN_6559;
      end
    end else begin
      btb_415_tag <= _GEN_6559;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_415_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19f == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_415_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_415_target_address <= _GEN_11999;
      end
    end else begin
      btb_415_target_address <= _GEN_11999;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_415_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h19f == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_415_bht <= 2'h1;
        end else begin
          btb_415_bht <= 2'h0;
        end
      end else begin
        btb_415_bht <= _GEN_12001;
      end
    end else begin
      btb_415_bht <= _GEN_12001;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_416_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_416_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_416_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_416_valid <= _GEN_15778;
      end
    end else begin
      btb_416_valid <= _GEN_15778;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_416_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_416_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_416_tag <= _GEN_6560;
      end
    end else begin
      btb_416_tag <= _GEN_6560;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_416_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_416_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_416_target_address <= _GEN_12002;
      end
    end else begin
      btb_416_target_address <= _GEN_12002;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_416_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_416_bht <= 2'h1;
        end else begin
          btb_416_bht <= 2'h0;
        end
      end else begin
        btb_416_bht <= _GEN_12004;
      end
    end else begin
      btb_416_bht <= _GEN_12004;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_417_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_417_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_417_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_417_valid <= _GEN_15779;
      end
    end else begin
      btb_417_valid <= _GEN_15779;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_417_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_417_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_417_tag <= _GEN_6561;
      end
    end else begin
      btb_417_tag <= _GEN_6561;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_417_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_417_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_417_target_address <= _GEN_12005;
      end
    end else begin
      btb_417_target_address <= _GEN_12005;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_417_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_417_bht <= 2'h1;
        end else begin
          btb_417_bht <= 2'h0;
        end
      end else begin
        btb_417_bht <= _GEN_12007;
      end
    end else begin
      btb_417_bht <= _GEN_12007;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_418_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_418_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_418_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_418_valid <= _GEN_15780;
      end
    end else begin
      btb_418_valid <= _GEN_15780;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_418_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_418_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_418_tag <= _GEN_6562;
      end
    end else begin
      btb_418_tag <= _GEN_6562;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_418_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_418_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_418_target_address <= _GEN_12008;
      end
    end else begin
      btb_418_target_address <= _GEN_12008;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_418_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_418_bht <= 2'h1;
        end else begin
          btb_418_bht <= 2'h0;
        end
      end else begin
        btb_418_bht <= _GEN_12010;
      end
    end else begin
      btb_418_bht <= _GEN_12010;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_419_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_419_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_419_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_419_valid <= _GEN_15781;
      end
    end else begin
      btb_419_valid <= _GEN_15781;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_419_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_419_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_419_tag <= _GEN_6563;
      end
    end else begin
      btb_419_tag <= _GEN_6563;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_419_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_419_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_419_target_address <= _GEN_12011;
      end
    end else begin
      btb_419_target_address <= _GEN_12011;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_419_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_419_bht <= 2'h1;
        end else begin
          btb_419_bht <= 2'h0;
        end
      end else begin
        btb_419_bht <= _GEN_12013;
      end
    end else begin
      btb_419_bht <= _GEN_12013;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_420_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_420_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_420_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_420_valid <= _GEN_15782;
      end
    end else begin
      btb_420_valid <= _GEN_15782;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_420_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_420_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_420_tag <= _GEN_6564;
      end
    end else begin
      btb_420_tag <= _GEN_6564;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_420_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_420_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_420_target_address <= _GEN_12014;
      end
    end else begin
      btb_420_target_address <= _GEN_12014;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_420_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_420_bht <= 2'h1;
        end else begin
          btb_420_bht <= 2'h0;
        end
      end else begin
        btb_420_bht <= _GEN_12016;
      end
    end else begin
      btb_420_bht <= _GEN_12016;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_421_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_421_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_421_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_421_valid <= _GEN_15783;
      end
    end else begin
      btb_421_valid <= _GEN_15783;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_421_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_421_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_421_tag <= _GEN_6565;
      end
    end else begin
      btb_421_tag <= _GEN_6565;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_421_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_421_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_421_target_address <= _GEN_12017;
      end
    end else begin
      btb_421_target_address <= _GEN_12017;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_421_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_421_bht <= 2'h1;
        end else begin
          btb_421_bht <= 2'h0;
        end
      end else begin
        btb_421_bht <= _GEN_12019;
      end
    end else begin
      btb_421_bht <= _GEN_12019;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_422_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_422_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_422_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_422_valid <= _GEN_15784;
      end
    end else begin
      btb_422_valid <= _GEN_15784;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_422_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_422_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_422_tag <= _GEN_6566;
      end
    end else begin
      btb_422_tag <= _GEN_6566;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_422_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_422_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_422_target_address <= _GEN_12020;
      end
    end else begin
      btb_422_target_address <= _GEN_12020;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_422_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_422_bht <= 2'h1;
        end else begin
          btb_422_bht <= 2'h0;
        end
      end else begin
        btb_422_bht <= _GEN_12022;
      end
    end else begin
      btb_422_bht <= _GEN_12022;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_423_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_423_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_423_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_423_valid <= _GEN_15785;
      end
    end else begin
      btb_423_valid <= _GEN_15785;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_423_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_423_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_423_tag <= _GEN_6567;
      end
    end else begin
      btb_423_tag <= _GEN_6567;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_423_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_423_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_423_target_address <= _GEN_12023;
      end
    end else begin
      btb_423_target_address <= _GEN_12023;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_423_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_423_bht <= 2'h1;
        end else begin
          btb_423_bht <= 2'h0;
        end
      end else begin
        btb_423_bht <= _GEN_12025;
      end
    end else begin
      btb_423_bht <= _GEN_12025;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_424_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_424_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_424_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_424_valid <= _GEN_15786;
      end
    end else begin
      btb_424_valid <= _GEN_15786;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_424_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_424_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_424_tag <= _GEN_6568;
      end
    end else begin
      btb_424_tag <= _GEN_6568;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_424_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_424_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_424_target_address <= _GEN_12026;
      end
    end else begin
      btb_424_target_address <= _GEN_12026;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_424_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_424_bht <= 2'h1;
        end else begin
          btb_424_bht <= 2'h0;
        end
      end else begin
        btb_424_bht <= _GEN_12028;
      end
    end else begin
      btb_424_bht <= _GEN_12028;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_425_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_425_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_425_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_425_valid <= _GEN_15787;
      end
    end else begin
      btb_425_valid <= _GEN_15787;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_425_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_425_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_425_tag <= _GEN_6569;
      end
    end else begin
      btb_425_tag <= _GEN_6569;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_425_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_425_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_425_target_address <= _GEN_12029;
      end
    end else begin
      btb_425_target_address <= _GEN_12029;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_425_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1a9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_425_bht <= 2'h1;
        end else begin
          btb_425_bht <= 2'h0;
        end
      end else begin
        btb_425_bht <= _GEN_12031;
      end
    end else begin
      btb_425_bht <= _GEN_12031;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_426_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_426_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_426_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_426_valid <= _GEN_15788;
      end
    end else begin
      btb_426_valid <= _GEN_15788;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_426_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1aa == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_426_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_426_tag <= _GEN_6570;
      end
    end else begin
      btb_426_tag <= _GEN_6570;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_426_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1aa == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_426_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_426_target_address <= _GEN_12032;
      end
    end else begin
      btb_426_target_address <= _GEN_12032;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_426_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1aa == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_426_bht <= 2'h1;
        end else begin
          btb_426_bht <= 2'h0;
        end
      end else begin
        btb_426_bht <= _GEN_12034;
      end
    end else begin
      btb_426_bht <= _GEN_12034;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_427_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_427_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_427_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_427_valid <= _GEN_15789;
      end
    end else begin
      btb_427_valid <= _GEN_15789;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_427_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ab == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_427_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_427_tag <= _GEN_6571;
      end
    end else begin
      btb_427_tag <= _GEN_6571;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_427_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ab == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_427_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_427_target_address <= _GEN_12035;
      end
    end else begin
      btb_427_target_address <= _GEN_12035;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_427_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ab == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_427_bht <= 2'h1;
        end else begin
          btb_427_bht <= 2'h0;
        end
      end else begin
        btb_427_bht <= _GEN_12037;
      end
    end else begin
      btb_427_bht <= _GEN_12037;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_428_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_428_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_428_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_428_valid <= _GEN_15790;
      end
    end else begin
      btb_428_valid <= _GEN_15790;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_428_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ac == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_428_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_428_tag <= _GEN_6572;
      end
    end else begin
      btb_428_tag <= _GEN_6572;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_428_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ac == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_428_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_428_target_address <= _GEN_12038;
      end
    end else begin
      btb_428_target_address <= _GEN_12038;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_428_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ac == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_428_bht <= 2'h1;
        end else begin
          btb_428_bht <= 2'h0;
        end
      end else begin
        btb_428_bht <= _GEN_12040;
      end
    end else begin
      btb_428_bht <= _GEN_12040;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_429_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_429_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_429_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_429_valid <= _GEN_15791;
      end
    end else begin
      btb_429_valid <= _GEN_15791;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_429_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ad == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_429_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_429_tag <= _GEN_6573;
      end
    end else begin
      btb_429_tag <= _GEN_6573;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_429_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ad == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_429_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_429_target_address <= _GEN_12041;
      end
    end else begin
      btb_429_target_address <= _GEN_12041;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_429_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ad == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_429_bht <= 2'h1;
        end else begin
          btb_429_bht <= 2'h0;
        end
      end else begin
        btb_429_bht <= _GEN_12043;
      end
    end else begin
      btb_429_bht <= _GEN_12043;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_430_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_430_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_430_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_430_valid <= _GEN_15792;
      end
    end else begin
      btb_430_valid <= _GEN_15792;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_430_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ae == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_430_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_430_tag <= _GEN_6574;
      end
    end else begin
      btb_430_tag <= _GEN_6574;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_430_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ae == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_430_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_430_target_address <= _GEN_12044;
      end
    end else begin
      btb_430_target_address <= _GEN_12044;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_430_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ae == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_430_bht <= 2'h1;
        end else begin
          btb_430_bht <= 2'h0;
        end
      end else begin
        btb_430_bht <= _GEN_12046;
      end
    end else begin
      btb_430_bht <= _GEN_12046;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_431_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_431_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_431_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_431_valid <= _GEN_15793;
      end
    end else begin
      btb_431_valid <= _GEN_15793;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_431_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1af == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_431_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_431_tag <= _GEN_6575;
      end
    end else begin
      btb_431_tag <= _GEN_6575;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_431_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1af == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_431_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_431_target_address <= _GEN_12047;
      end
    end else begin
      btb_431_target_address <= _GEN_12047;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_431_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1af == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_431_bht <= 2'h1;
        end else begin
          btb_431_bht <= 2'h0;
        end
      end else begin
        btb_431_bht <= _GEN_12049;
      end
    end else begin
      btb_431_bht <= _GEN_12049;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_432_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_432_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_432_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_432_valid <= _GEN_15794;
      end
    end else begin
      btb_432_valid <= _GEN_15794;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_432_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_432_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_432_tag <= _GEN_6576;
      end
    end else begin
      btb_432_tag <= _GEN_6576;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_432_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_432_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_432_target_address <= _GEN_12050;
      end
    end else begin
      btb_432_target_address <= _GEN_12050;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_432_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_432_bht <= 2'h1;
        end else begin
          btb_432_bht <= 2'h0;
        end
      end else begin
        btb_432_bht <= _GEN_12052;
      end
    end else begin
      btb_432_bht <= _GEN_12052;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_433_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_433_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_433_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_433_valid <= _GEN_15795;
      end
    end else begin
      btb_433_valid <= _GEN_15795;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_433_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_433_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_433_tag <= _GEN_6577;
      end
    end else begin
      btb_433_tag <= _GEN_6577;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_433_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_433_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_433_target_address <= _GEN_12053;
      end
    end else begin
      btb_433_target_address <= _GEN_12053;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_433_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_433_bht <= 2'h1;
        end else begin
          btb_433_bht <= 2'h0;
        end
      end else begin
        btb_433_bht <= _GEN_12055;
      end
    end else begin
      btb_433_bht <= _GEN_12055;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_434_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_434_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_434_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_434_valid <= _GEN_15796;
      end
    end else begin
      btb_434_valid <= _GEN_15796;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_434_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_434_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_434_tag <= _GEN_6578;
      end
    end else begin
      btb_434_tag <= _GEN_6578;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_434_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_434_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_434_target_address <= _GEN_12056;
      end
    end else begin
      btb_434_target_address <= _GEN_12056;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_434_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_434_bht <= 2'h1;
        end else begin
          btb_434_bht <= 2'h0;
        end
      end else begin
        btb_434_bht <= _GEN_12058;
      end
    end else begin
      btb_434_bht <= _GEN_12058;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_435_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_435_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_435_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_435_valid <= _GEN_15797;
      end
    end else begin
      btb_435_valid <= _GEN_15797;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_435_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_435_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_435_tag <= _GEN_6579;
      end
    end else begin
      btb_435_tag <= _GEN_6579;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_435_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_435_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_435_target_address <= _GEN_12059;
      end
    end else begin
      btb_435_target_address <= _GEN_12059;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_435_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_435_bht <= 2'h1;
        end else begin
          btb_435_bht <= 2'h0;
        end
      end else begin
        btb_435_bht <= _GEN_12061;
      end
    end else begin
      btb_435_bht <= _GEN_12061;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_436_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_436_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_436_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_436_valid <= _GEN_15798;
      end
    end else begin
      btb_436_valid <= _GEN_15798;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_436_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_436_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_436_tag <= _GEN_6580;
      end
    end else begin
      btb_436_tag <= _GEN_6580;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_436_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_436_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_436_target_address <= _GEN_12062;
      end
    end else begin
      btb_436_target_address <= _GEN_12062;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_436_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_436_bht <= 2'h1;
        end else begin
          btb_436_bht <= 2'h0;
        end
      end else begin
        btb_436_bht <= _GEN_12064;
      end
    end else begin
      btb_436_bht <= _GEN_12064;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_437_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_437_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_437_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_437_valid <= _GEN_15799;
      end
    end else begin
      btb_437_valid <= _GEN_15799;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_437_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_437_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_437_tag <= _GEN_6581;
      end
    end else begin
      btb_437_tag <= _GEN_6581;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_437_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_437_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_437_target_address <= _GEN_12065;
      end
    end else begin
      btb_437_target_address <= _GEN_12065;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_437_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_437_bht <= 2'h1;
        end else begin
          btb_437_bht <= 2'h0;
        end
      end else begin
        btb_437_bht <= _GEN_12067;
      end
    end else begin
      btb_437_bht <= _GEN_12067;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_438_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_438_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_438_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_438_valid <= _GEN_15800;
      end
    end else begin
      btb_438_valid <= _GEN_15800;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_438_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_438_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_438_tag <= _GEN_6582;
      end
    end else begin
      btb_438_tag <= _GEN_6582;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_438_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_438_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_438_target_address <= _GEN_12068;
      end
    end else begin
      btb_438_target_address <= _GEN_12068;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_438_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_438_bht <= 2'h1;
        end else begin
          btb_438_bht <= 2'h0;
        end
      end else begin
        btb_438_bht <= _GEN_12070;
      end
    end else begin
      btb_438_bht <= _GEN_12070;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_439_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_439_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_439_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_439_valid <= _GEN_15801;
      end
    end else begin
      btb_439_valid <= _GEN_15801;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_439_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_439_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_439_tag <= _GEN_6583;
      end
    end else begin
      btb_439_tag <= _GEN_6583;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_439_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_439_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_439_target_address <= _GEN_12071;
      end
    end else begin
      btb_439_target_address <= _GEN_12071;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_439_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_439_bht <= 2'h1;
        end else begin
          btb_439_bht <= 2'h0;
        end
      end else begin
        btb_439_bht <= _GEN_12073;
      end
    end else begin
      btb_439_bht <= _GEN_12073;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_440_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_440_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_440_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_440_valid <= _GEN_15802;
      end
    end else begin
      btb_440_valid <= _GEN_15802;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_440_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_440_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_440_tag <= _GEN_6584;
      end
    end else begin
      btb_440_tag <= _GEN_6584;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_440_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_440_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_440_target_address <= _GEN_12074;
      end
    end else begin
      btb_440_target_address <= _GEN_12074;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_440_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_440_bht <= 2'h1;
        end else begin
          btb_440_bht <= 2'h0;
        end
      end else begin
        btb_440_bht <= _GEN_12076;
      end
    end else begin
      btb_440_bht <= _GEN_12076;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_441_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_441_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_441_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_441_valid <= _GEN_15803;
      end
    end else begin
      btb_441_valid <= _GEN_15803;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_441_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_441_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_441_tag <= _GEN_6585;
      end
    end else begin
      btb_441_tag <= _GEN_6585;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_441_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_441_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_441_target_address <= _GEN_12077;
      end
    end else begin
      btb_441_target_address <= _GEN_12077;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_441_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1b9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_441_bht <= 2'h1;
        end else begin
          btb_441_bht <= 2'h0;
        end
      end else begin
        btb_441_bht <= _GEN_12079;
      end
    end else begin
      btb_441_bht <= _GEN_12079;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_442_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_442_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_442_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_442_valid <= _GEN_15804;
      end
    end else begin
      btb_442_valid <= _GEN_15804;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_442_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ba == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_442_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_442_tag <= _GEN_6586;
      end
    end else begin
      btb_442_tag <= _GEN_6586;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_442_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ba == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_442_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_442_target_address <= _GEN_12080;
      end
    end else begin
      btb_442_target_address <= _GEN_12080;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_442_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ba == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_442_bht <= 2'h1;
        end else begin
          btb_442_bht <= 2'h0;
        end
      end else begin
        btb_442_bht <= _GEN_12082;
      end
    end else begin
      btb_442_bht <= _GEN_12082;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_443_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_443_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_443_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_443_valid <= _GEN_15805;
      end
    end else begin
      btb_443_valid <= _GEN_15805;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_443_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_443_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_443_tag <= _GEN_6587;
      end
    end else begin
      btb_443_tag <= _GEN_6587;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_443_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_443_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_443_target_address <= _GEN_12083;
      end
    end else begin
      btb_443_target_address <= _GEN_12083;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_443_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_443_bht <= 2'h1;
        end else begin
          btb_443_bht <= 2'h0;
        end
      end else begin
        btb_443_bht <= _GEN_12085;
      end
    end else begin
      btb_443_bht <= _GEN_12085;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_444_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_444_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_444_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_444_valid <= _GEN_15806;
      end
    end else begin
      btb_444_valid <= _GEN_15806;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_444_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_444_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_444_tag <= _GEN_6588;
      end
    end else begin
      btb_444_tag <= _GEN_6588;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_444_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_444_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_444_target_address <= _GEN_12086;
      end
    end else begin
      btb_444_target_address <= _GEN_12086;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_444_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_444_bht <= 2'h1;
        end else begin
          btb_444_bht <= 2'h0;
        end
      end else begin
        btb_444_bht <= _GEN_12088;
      end
    end else begin
      btb_444_bht <= _GEN_12088;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_445_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_445_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_445_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_445_valid <= _GEN_15807;
      end
    end else begin
      btb_445_valid <= _GEN_15807;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_445_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_445_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_445_tag <= _GEN_6589;
      end
    end else begin
      btb_445_tag <= _GEN_6589;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_445_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_445_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_445_target_address <= _GEN_12089;
      end
    end else begin
      btb_445_target_address <= _GEN_12089;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_445_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_445_bht <= 2'h1;
        end else begin
          btb_445_bht <= 2'h0;
        end
      end else begin
        btb_445_bht <= _GEN_12091;
      end
    end else begin
      btb_445_bht <= _GEN_12091;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_446_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_446_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_446_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_446_valid <= _GEN_15808;
      end
    end else begin
      btb_446_valid <= _GEN_15808;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_446_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1be == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_446_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_446_tag <= _GEN_6590;
      end
    end else begin
      btb_446_tag <= _GEN_6590;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_446_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1be == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_446_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_446_target_address <= _GEN_12092;
      end
    end else begin
      btb_446_target_address <= _GEN_12092;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_446_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1be == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_446_bht <= 2'h1;
        end else begin
          btb_446_bht <= 2'h0;
        end
      end else begin
        btb_446_bht <= _GEN_12094;
      end
    end else begin
      btb_446_bht <= _GEN_12094;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_447_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_447_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_447_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_447_valid <= _GEN_15809;
      end
    end else begin
      btb_447_valid <= _GEN_15809;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_447_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_447_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_447_tag <= _GEN_6591;
      end
    end else begin
      btb_447_tag <= _GEN_6591;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_447_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_447_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_447_target_address <= _GEN_12095;
      end
    end else begin
      btb_447_target_address <= _GEN_12095;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_447_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1bf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_447_bht <= 2'h1;
        end else begin
          btb_447_bht <= 2'h0;
        end
      end else begin
        btb_447_bht <= _GEN_12097;
      end
    end else begin
      btb_447_bht <= _GEN_12097;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_448_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_448_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_448_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_448_valid <= _GEN_15810;
      end
    end else begin
      btb_448_valid <= _GEN_15810;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_448_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_448_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_448_tag <= _GEN_6592;
      end
    end else begin
      btb_448_tag <= _GEN_6592;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_448_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_448_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_448_target_address <= _GEN_12098;
      end
    end else begin
      btb_448_target_address <= _GEN_12098;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_448_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_448_bht <= 2'h1;
        end else begin
          btb_448_bht <= 2'h0;
        end
      end else begin
        btb_448_bht <= _GEN_12100;
      end
    end else begin
      btb_448_bht <= _GEN_12100;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_449_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_449_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_449_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_449_valid <= _GEN_15811;
      end
    end else begin
      btb_449_valid <= _GEN_15811;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_449_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_449_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_449_tag <= _GEN_6593;
      end
    end else begin
      btb_449_tag <= _GEN_6593;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_449_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_449_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_449_target_address <= _GEN_12101;
      end
    end else begin
      btb_449_target_address <= _GEN_12101;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_449_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_449_bht <= 2'h1;
        end else begin
          btb_449_bht <= 2'h0;
        end
      end else begin
        btb_449_bht <= _GEN_12103;
      end
    end else begin
      btb_449_bht <= _GEN_12103;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_450_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_450_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_450_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_450_valid <= _GEN_15812;
      end
    end else begin
      btb_450_valid <= _GEN_15812;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_450_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_450_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_450_tag <= _GEN_6594;
      end
    end else begin
      btb_450_tag <= _GEN_6594;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_450_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_450_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_450_target_address <= _GEN_12104;
      end
    end else begin
      btb_450_target_address <= _GEN_12104;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_450_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_450_bht <= 2'h1;
        end else begin
          btb_450_bht <= 2'h0;
        end
      end else begin
        btb_450_bht <= _GEN_12106;
      end
    end else begin
      btb_450_bht <= _GEN_12106;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_451_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_451_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_451_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_451_valid <= _GEN_15813;
      end
    end else begin
      btb_451_valid <= _GEN_15813;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_451_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_451_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_451_tag <= _GEN_6595;
      end
    end else begin
      btb_451_tag <= _GEN_6595;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_451_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_451_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_451_target_address <= _GEN_12107;
      end
    end else begin
      btb_451_target_address <= _GEN_12107;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_451_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_451_bht <= 2'h1;
        end else begin
          btb_451_bht <= 2'h0;
        end
      end else begin
        btb_451_bht <= _GEN_12109;
      end
    end else begin
      btb_451_bht <= _GEN_12109;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_452_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_452_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_452_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_452_valid <= _GEN_15814;
      end
    end else begin
      btb_452_valid <= _GEN_15814;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_452_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_452_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_452_tag <= _GEN_6596;
      end
    end else begin
      btb_452_tag <= _GEN_6596;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_452_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_452_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_452_target_address <= _GEN_12110;
      end
    end else begin
      btb_452_target_address <= _GEN_12110;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_452_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_452_bht <= 2'h1;
        end else begin
          btb_452_bht <= 2'h0;
        end
      end else begin
        btb_452_bht <= _GEN_12112;
      end
    end else begin
      btb_452_bht <= _GEN_12112;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_453_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_453_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_453_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_453_valid <= _GEN_15815;
      end
    end else begin
      btb_453_valid <= _GEN_15815;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_453_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_453_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_453_tag <= _GEN_6597;
      end
    end else begin
      btb_453_tag <= _GEN_6597;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_453_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_453_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_453_target_address <= _GEN_12113;
      end
    end else begin
      btb_453_target_address <= _GEN_12113;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_453_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_453_bht <= 2'h1;
        end else begin
          btb_453_bht <= 2'h0;
        end
      end else begin
        btb_453_bht <= _GEN_12115;
      end
    end else begin
      btb_453_bht <= _GEN_12115;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_454_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_454_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_454_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_454_valid <= _GEN_15816;
      end
    end else begin
      btb_454_valid <= _GEN_15816;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_454_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_454_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_454_tag <= _GEN_6598;
      end
    end else begin
      btb_454_tag <= _GEN_6598;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_454_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_454_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_454_target_address <= _GEN_12116;
      end
    end else begin
      btb_454_target_address <= _GEN_12116;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_454_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_454_bht <= 2'h1;
        end else begin
          btb_454_bht <= 2'h0;
        end
      end else begin
        btb_454_bht <= _GEN_12118;
      end
    end else begin
      btb_454_bht <= _GEN_12118;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_455_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_455_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_455_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_455_valid <= _GEN_15817;
      end
    end else begin
      btb_455_valid <= _GEN_15817;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_455_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_455_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_455_tag <= _GEN_6599;
      end
    end else begin
      btb_455_tag <= _GEN_6599;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_455_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_455_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_455_target_address <= _GEN_12119;
      end
    end else begin
      btb_455_target_address <= _GEN_12119;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_455_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_455_bht <= 2'h1;
        end else begin
          btb_455_bht <= 2'h0;
        end
      end else begin
        btb_455_bht <= _GEN_12121;
      end
    end else begin
      btb_455_bht <= _GEN_12121;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_456_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_456_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_456_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_456_valid <= _GEN_15818;
      end
    end else begin
      btb_456_valid <= _GEN_15818;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_456_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_456_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_456_tag <= _GEN_6600;
      end
    end else begin
      btb_456_tag <= _GEN_6600;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_456_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_456_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_456_target_address <= _GEN_12122;
      end
    end else begin
      btb_456_target_address <= _GEN_12122;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_456_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_456_bht <= 2'h1;
        end else begin
          btb_456_bht <= 2'h0;
        end
      end else begin
        btb_456_bht <= _GEN_12124;
      end
    end else begin
      btb_456_bht <= _GEN_12124;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_457_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_457_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_457_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_457_valid <= _GEN_15819;
      end
    end else begin
      btb_457_valid <= _GEN_15819;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_457_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_457_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_457_tag <= _GEN_6601;
      end
    end else begin
      btb_457_tag <= _GEN_6601;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_457_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_457_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_457_target_address <= _GEN_12125;
      end
    end else begin
      btb_457_target_address <= _GEN_12125;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_457_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1c9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_457_bht <= 2'h1;
        end else begin
          btb_457_bht <= 2'h0;
        end
      end else begin
        btb_457_bht <= _GEN_12127;
      end
    end else begin
      btb_457_bht <= _GEN_12127;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_458_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_458_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_458_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_458_valid <= _GEN_15820;
      end
    end else begin
      btb_458_valid <= _GEN_15820;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_458_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ca == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_458_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_458_tag <= _GEN_6602;
      end
    end else begin
      btb_458_tag <= _GEN_6602;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_458_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ca == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_458_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_458_target_address <= _GEN_12128;
      end
    end else begin
      btb_458_target_address <= _GEN_12128;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_458_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ca == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_458_bht <= 2'h1;
        end else begin
          btb_458_bht <= 2'h0;
        end
      end else begin
        btb_458_bht <= _GEN_12130;
      end
    end else begin
      btb_458_bht <= _GEN_12130;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_459_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_459_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_459_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_459_valid <= _GEN_15821;
      end
    end else begin
      btb_459_valid <= _GEN_15821;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_459_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_459_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_459_tag <= _GEN_6603;
      end
    end else begin
      btb_459_tag <= _GEN_6603;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_459_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_459_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_459_target_address <= _GEN_12131;
      end
    end else begin
      btb_459_target_address <= _GEN_12131;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_459_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_459_bht <= 2'h1;
        end else begin
          btb_459_bht <= 2'h0;
        end
      end else begin
        btb_459_bht <= _GEN_12133;
      end
    end else begin
      btb_459_bht <= _GEN_12133;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_460_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_460_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_460_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_460_valid <= _GEN_15822;
      end
    end else begin
      btb_460_valid <= _GEN_15822;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_460_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_460_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_460_tag <= _GEN_6604;
      end
    end else begin
      btb_460_tag <= _GEN_6604;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_460_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_460_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_460_target_address <= _GEN_12134;
      end
    end else begin
      btb_460_target_address <= _GEN_12134;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_460_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_460_bht <= 2'h1;
        end else begin
          btb_460_bht <= 2'h0;
        end
      end else begin
        btb_460_bht <= _GEN_12136;
      end
    end else begin
      btb_460_bht <= _GEN_12136;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_461_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_461_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_461_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_461_valid <= _GEN_15823;
      end
    end else begin
      btb_461_valid <= _GEN_15823;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_461_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_461_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_461_tag <= _GEN_6605;
      end
    end else begin
      btb_461_tag <= _GEN_6605;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_461_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_461_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_461_target_address <= _GEN_12137;
      end
    end else begin
      btb_461_target_address <= _GEN_12137;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_461_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_461_bht <= 2'h1;
        end else begin
          btb_461_bht <= 2'h0;
        end
      end else begin
        btb_461_bht <= _GEN_12139;
      end
    end else begin
      btb_461_bht <= _GEN_12139;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_462_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_462_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_462_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_462_valid <= _GEN_15824;
      end
    end else begin
      btb_462_valid <= _GEN_15824;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_462_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ce == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_462_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_462_tag <= _GEN_6606;
      end
    end else begin
      btb_462_tag <= _GEN_6606;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_462_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ce == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_462_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_462_target_address <= _GEN_12140;
      end
    end else begin
      btb_462_target_address <= _GEN_12140;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_462_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ce == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_462_bht <= 2'h1;
        end else begin
          btb_462_bht <= 2'h0;
        end
      end else begin
        btb_462_bht <= _GEN_12142;
      end
    end else begin
      btb_462_bht <= _GEN_12142;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_463_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_463_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_463_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_463_valid <= _GEN_15825;
      end
    end else begin
      btb_463_valid <= _GEN_15825;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_463_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cf == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_463_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_463_tag <= _GEN_6607;
      end
    end else begin
      btb_463_tag <= _GEN_6607;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_463_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cf == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_463_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_463_target_address <= _GEN_12143;
      end
    end else begin
      btb_463_target_address <= _GEN_12143;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_463_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1cf == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_463_bht <= 2'h1;
        end else begin
          btb_463_bht <= 2'h0;
        end
      end else begin
        btb_463_bht <= _GEN_12145;
      end
    end else begin
      btb_463_bht <= _GEN_12145;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_464_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_464_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_464_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_464_valid <= _GEN_15826;
      end
    end else begin
      btb_464_valid <= _GEN_15826;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_464_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_464_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_464_tag <= _GEN_6608;
      end
    end else begin
      btb_464_tag <= _GEN_6608;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_464_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_464_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_464_target_address <= _GEN_12146;
      end
    end else begin
      btb_464_target_address <= _GEN_12146;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_464_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_464_bht <= 2'h1;
        end else begin
          btb_464_bht <= 2'h0;
        end
      end else begin
        btb_464_bht <= _GEN_12148;
      end
    end else begin
      btb_464_bht <= _GEN_12148;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_465_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_465_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_465_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_465_valid <= _GEN_15827;
      end
    end else begin
      btb_465_valid <= _GEN_15827;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_465_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_465_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_465_tag <= _GEN_6609;
      end
    end else begin
      btb_465_tag <= _GEN_6609;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_465_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_465_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_465_target_address <= _GEN_12149;
      end
    end else begin
      btb_465_target_address <= _GEN_12149;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_465_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_465_bht <= 2'h1;
        end else begin
          btb_465_bht <= 2'h0;
        end
      end else begin
        btb_465_bht <= _GEN_12151;
      end
    end else begin
      btb_465_bht <= _GEN_12151;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_466_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_466_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_466_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_466_valid <= _GEN_15828;
      end
    end else begin
      btb_466_valid <= _GEN_15828;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_466_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_466_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_466_tag <= _GEN_6610;
      end
    end else begin
      btb_466_tag <= _GEN_6610;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_466_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_466_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_466_target_address <= _GEN_12152;
      end
    end else begin
      btb_466_target_address <= _GEN_12152;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_466_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_466_bht <= 2'h1;
        end else begin
          btb_466_bht <= 2'h0;
        end
      end else begin
        btb_466_bht <= _GEN_12154;
      end
    end else begin
      btb_466_bht <= _GEN_12154;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_467_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_467_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_467_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_467_valid <= _GEN_15829;
      end
    end else begin
      btb_467_valid <= _GEN_15829;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_467_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_467_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_467_tag <= _GEN_6611;
      end
    end else begin
      btb_467_tag <= _GEN_6611;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_467_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_467_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_467_target_address <= _GEN_12155;
      end
    end else begin
      btb_467_target_address <= _GEN_12155;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_467_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_467_bht <= 2'h1;
        end else begin
          btb_467_bht <= 2'h0;
        end
      end else begin
        btb_467_bht <= _GEN_12157;
      end
    end else begin
      btb_467_bht <= _GEN_12157;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_468_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_468_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_468_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_468_valid <= _GEN_15830;
      end
    end else begin
      btb_468_valid <= _GEN_15830;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_468_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_468_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_468_tag <= _GEN_6612;
      end
    end else begin
      btb_468_tag <= _GEN_6612;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_468_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_468_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_468_target_address <= _GEN_12158;
      end
    end else begin
      btb_468_target_address <= _GEN_12158;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_468_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_468_bht <= 2'h1;
        end else begin
          btb_468_bht <= 2'h0;
        end
      end else begin
        btb_468_bht <= _GEN_12160;
      end
    end else begin
      btb_468_bht <= _GEN_12160;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_469_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_469_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_469_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_469_valid <= _GEN_15831;
      end
    end else begin
      btb_469_valid <= _GEN_15831;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_469_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_469_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_469_tag <= _GEN_6613;
      end
    end else begin
      btb_469_tag <= _GEN_6613;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_469_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_469_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_469_target_address <= _GEN_12161;
      end
    end else begin
      btb_469_target_address <= _GEN_12161;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_469_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_469_bht <= 2'h1;
        end else begin
          btb_469_bht <= 2'h0;
        end
      end else begin
        btb_469_bht <= _GEN_12163;
      end
    end else begin
      btb_469_bht <= _GEN_12163;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_470_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_470_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_470_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_470_valid <= _GEN_15832;
      end
    end else begin
      btb_470_valid <= _GEN_15832;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_470_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_470_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_470_tag <= _GEN_6614;
      end
    end else begin
      btb_470_tag <= _GEN_6614;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_470_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_470_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_470_target_address <= _GEN_12164;
      end
    end else begin
      btb_470_target_address <= _GEN_12164;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_470_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_470_bht <= 2'h1;
        end else begin
          btb_470_bht <= 2'h0;
        end
      end else begin
        btb_470_bht <= _GEN_12166;
      end
    end else begin
      btb_470_bht <= _GEN_12166;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_471_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_471_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_471_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_471_valid <= _GEN_15833;
      end
    end else begin
      btb_471_valid <= _GEN_15833;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_471_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_471_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_471_tag <= _GEN_6615;
      end
    end else begin
      btb_471_tag <= _GEN_6615;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_471_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_471_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_471_target_address <= _GEN_12167;
      end
    end else begin
      btb_471_target_address <= _GEN_12167;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_471_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_471_bht <= 2'h1;
        end else begin
          btb_471_bht <= 2'h0;
        end
      end else begin
        btb_471_bht <= _GEN_12169;
      end
    end else begin
      btb_471_bht <= _GEN_12169;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_472_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_472_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_472_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_472_valid <= _GEN_15834;
      end
    end else begin
      btb_472_valid <= _GEN_15834;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_472_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_472_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_472_tag <= _GEN_6616;
      end
    end else begin
      btb_472_tag <= _GEN_6616;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_472_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_472_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_472_target_address <= _GEN_12170;
      end
    end else begin
      btb_472_target_address <= _GEN_12170;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_472_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_472_bht <= 2'h1;
        end else begin
          btb_472_bht <= 2'h0;
        end
      end else begin
        btb_472_bht <= _GEN_12172;
      end
    end else begin
      btb_472_bht <= _GEN_12172;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_473_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_473_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_473_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_473_valid <= _GEN_15835;
      end
    end else begin
      btb_473_valid <= _GEN_15835;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_473_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_473_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_473_tag <= _GEN_6617;
      end
    end else begin
      btb_473_tag <= _GEN_6617;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_473_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_473_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_473_target_address <= _GEN_12173;
      end
    end else begin
      btb_473_target_address <= _GEN_12173;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_473_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1d9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_473_bht <= 2'h1;
        end else begin
          btb_473_bht <= 2'h0;
        end
      end else begin
        btb_473_bht <= _GEN_12175;
      end
    end else begin
      btb_473_bht <= _GEN_12175;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_474_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_474_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_474_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_474_valid <= _GEN_15836;
      end
    end else begin
      btb_474_valid <= _GEN_15836;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_474_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1da == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_474_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_474_tag <= _GEN_6618;
      end
    end else begin
      btb_474_tag <= _GEN_6618;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_474_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1da == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_474_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_474_target_address <= _GEN_12176;
      end
    end else begin
      btb_474_target_address <= _GEN_12176;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_474_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1da == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_474_bht <= 2'h1;
        end else begin
          btb_474_bht <= 2'h0;
        end
      end else begin
        btb_474_bht <= _GEN_12178;
      end
    end else begin
      btb_474_bht <= _GEN_12178;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_475_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_475_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_475_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_475_valid <= _GEN_15837;
      end
    end else begin
      btb_475_valid <= _GEN_15837;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_475_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1db == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_475_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_475_tag <= _GEN_6619;
      end
    end else begin
      btb_475_tag <= _GEN_6619;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_475_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1db == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_475_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_475_target_address <= _GEN_12179;
      end
    end else begin
      btb_475_target_address <= _GEN_12179;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_475_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1db == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_475_bht <= 2'h1;
        end else begin
          btb_475_bht <= 2'h0;
        end
      end else begin
        btb_475_bht <= _GEN_12181;
      end
    end else begin
      btb_475_bht <= _GEN_12181;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_476_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_476_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_476_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_476_valid <= _GEN_15838;
      end
    end else begin
      btb_476_valid <= _GEN_15838;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_476_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1dc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_476_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_476_tag <= _GEN_6620;
      end
    end else begin
      btb_476_tag <= _GEN_6620;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_476_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1dc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_476_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_476_target_address <= _GEN_12182;
      end
    end else begin
      btb_476_target_address <= _GEN_12182;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_476_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1dc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_476_bht <= 2'h1;
        end else begin
          btb_476_bht <= 2'h0;
        end
      end else begin
        btb_476_bht <= _GEN_12184;
      end
    end else begin
      btb_476_bht <= _GEN_12184;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_477_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_477_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_477_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_477_valid <= _GEN_15839;
      end
    end else begin
      btb_477_valid <= _GEN_15839;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_477_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1dd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_477_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_477_tag <= _GEN_6621;
      end
    end else begin
      btb_477_tag <= _GEN_6621;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_477_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1dd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_477_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_477_target_address <= _GEN_12185;
      end
    end else begin
      btb_477_target_address <= _GEN_12185;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_477_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1dd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_477_bht <= 2'h1;
        end else begin
          btb_477_bht <= 2'h0;
        end
      end else begin
        btb_477_bht <= _GEN_12187;
      end
    end else begin
      btb_477_bht <= _GEN_12187;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_478_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_478_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_478_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_478_valid <= _GEN_15840;
      end
    end else begin
      btb_478_valid <= _GEN_15840;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_478_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1de == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_478_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_478_tag <= _GEN_6622;
      end
    end else begin
      btb_478_tag <= _GEN_6622;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_478_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1de == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_478_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_478_target_address <= _GEN_12188;
      end
    end else begin
      btb_478_target_address <= _GEN_12188;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_478_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1de == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_478_bht <= 2'h1;
        end else begin
          btb_478_bht <= 2'h0;
        end
      end else begin
        btb_478_bht <= _GEN_12190;
      end
    end else begin
      btb_478_bht <= _GEN_12190;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_479_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_479_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_479_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_479_valid <= _GEN_15841;
      end
    end else begin
      btb_479_valid <= _GEN_15841;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_479_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1df == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_479_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_479_tag <= _GEN_6623;
      end
    end else begin
      btb_479_tag <= _GEN_6623;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_479_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1df == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_479_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_479_target_address <= _GEN_12191;
      end
    end else begin
      btb_479_target_address <= _GEN_12191;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_479_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1df == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_479_bht <= 2'h1;
        end else begin
          btb_479_bht <= 2'h0;
        end
      end else begin
        btb_479_bht <= _GEN_12193;
      end
    end else begin
      btb_479_bht <= _GEN_12193;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_480_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_480_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_480_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_480_valid <= _GEN_15842;
      end
    end else begin
      btb_480_valid <= _GEN_15842;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_480_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_480_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_480_tag <= _GEN_6624;
      end
    end else begin
      btb_480_tag <= _GEN_6624;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_480_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_480_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_480_target_address <= _GEN_12194;
      end
    end else begin
      btb_480_target_address <= _GEN_12194;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_480_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_480_bht <= 2'h1;
        end else begin
          btb_480_bht <= 2'h0;
        end
      end else begin
        btb_480_bht <= _GEN_12196;
      end
    end else begin
      btb_480_bht <= _GEN_12196;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_481_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_481_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_481_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_481_valid <= _GEN_15843;
      end
    end else begin
      btb_481_valid <= _GEN_15843;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_481_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_481_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_481_tag <= _GEN_6625;
      end
    end else begin
      btb_481_tag <= _GEN_6625;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_481_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_481_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_481_target_address <= _GEN_12197;
      end
    end else begin
      btb_481_target_address <= _GEN_12197;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_481_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_481_bht <= 2'h1;
        end else begin
          btb_481_bht <= 2'h0;
        end
      end else begin
        btb_481_bht <= _GEN_12199;
      end
    end else begin
      btb_481_bht <= _GEN_12199;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_482_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_482_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_482_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_482_valid <= _GEN_15844;
      end
    end else begin
      btb_482_valid <= _GEN_15844;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_482_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_482_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_482_tag <= _GEN_6626;
      end
    end else begin
      btb_482_tag <= _GEN_6626;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_482_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_482_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_482_target_address <= _GEN_12200;
      end
    end else begin
      btb_482_target_address <= _GEN_12200;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_482_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_482_bht <= 2'h1;
        end else begin
          btb_482_bht <= 2'h0;
        end
      end else begin
        btb_482_bht <= _GEN_12202;
      end
    end else begin
      btb_482_bht <= _GEN_12202;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_483_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_483_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_483_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_483_valid <= _GEN_15845;
      end
    end else begin
      btb_483_valid <= _GEN_15845;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_483_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_483_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_483_tag <= _GEN_6627;
      end
    end else begin
      btb_483_tag <= _GEN_6627;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_483_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_483_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_483_target_address <= _GEN_12203;
      end
    end else begin
      btb_483_target_address <= _GEN_12203;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_483_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_483_bht <= 2'h1;
        end else begin
          btb_483_bht <= 2'h0;
        end
      end else begin
        btb_483_bht <= _GEN_12205;
      end
    end else begin
      btb_483_bht <= _GEN_12205;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_484_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_484_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_484_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_484_valid <= _GEN_15846;
      end
    end else begin
      btb_484_valid <= _GEN_15846;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_484_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_484_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_484_tag <= _GEN_6628;
      end
    end else begin
      btb_484_tag <= _GEN_6628;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_484_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_484_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_484_target_address <= _GEN_12206;
      end
    end else begin
      btb_484_target_address <= _GEN_12206;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_484_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_484_bht <= 2'h1;
        end else begin
          btb_484_bht <= 2'h0;
        end
      end else begin
        btb_484_bht <= _GEN_12208;
      end
    end else begin
      btb_484_bht <= _GEN_12208;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_485_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_485_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_485_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_485_valid <= _GEN_15847;
      end
    end else begin
      btb_485_valid <= _GEN_15847;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_485_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_485_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_485_tag <= _GEN_6629;
      end
    end else begin
      btb_485_tag <= _GEN_6629;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_485_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_485_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_485_target_address <= _GEN_12209;
      end
    end else begin
      btb_485_target_address <= _GEN_12209;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_485_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_485_bht <= 2'h1;
        end else begin
          btb_485_bht <= 2'h0;
        end
      end else begin
        btb_485_bht <= _GEN_12211;
      end
    end else begin
      btb_485_bht <= _GEN_12211;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_486_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_486_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_486_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_486_valid <= _GEN_15848;
      end
    end else begin
      btb_486_valid <= _GEN_15848;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_486_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_486_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_486_tag <= _GEN_6630;
      end
    end else begin
      btb_486_tag <= _GEN_6630;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_486_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_486_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_486_target_address <= _GEN_12212;
      end
    end else begin
      btb_486_target_address <= _GEN_12212;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_486_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_486_bht <= 2'h1;
        end else begin
          btb_486_bht <= 2'h0;
        end
      end else begin
        btb_486_bht <= _GEN_12214;
      end
    end else begin
      btb_486_bht <= _GEN_12214;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_487_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_487_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_487_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_487_valid <= _GEN_15849;
      end
    end else begin
      btb_487_valid <= _GEN_15849;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_487_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_487_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_487_tag <= _GEN_6631;
      end
    end else begin
      btb_487_tag <= _GEN_6631;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_487_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_487_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_487_target_address <= _GEN_12215;
      end
    end else begin
      btb_487_target_address <= _GEN_12215;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_487_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_487_bht <= 2'h1;
        end else begin
          btb_487_bht <= 2'h0;
        end
      end else begin
        btb_487_bht <= _GEN_12217;
      end
    end else begin
      btb_487_bht <= _GEN_12217;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_488_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_488_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_488_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_488_valid <= _GEN_15850;
      end
    end else begin
      btb_488_valid <= _GEN_15850;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_488_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_488_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_488_tag <= _GEN_6632;
      end
    end else begin
      btb_488_tag <= _GEN_6632;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_488_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_488_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_488_target_address <= _GEN_12218;
      end
    end else begin
      btb_488_target_address <= _GEN_12218;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_488_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_488_bht <= 2'h1;
        end else begin
          btb_488_bht <= 2'h0;
        end
      end else begin
        btb_488_bht <= _GEN_12220;
      end
    end else begin
      btb_488_bht <= _GEN_12220;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_489_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_489_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_489_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_489_valid <= _GEN_15851;
      end
    end else begin
      btb_489_valid <= _GEN_15851;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_489_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_489_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_489_tag <= _GEN_6633;
      end
    end else begin
      btb_489_tag <= _GEN_6633;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_489_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_489_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_489_target_address <= _GEN_12221;
      end
    end else begin
      btb_489_target_address <= _GEN_12221;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_489_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1e9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_489_bht <= 2'h1;
        end else begin
          btb_489_bht <= 2'h0;
        end
      end else begin
        btb_489_bht <= _GEN_12223;
      end
    end else begin
      btb_489_bht <= _GEN_12223;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_490_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_490_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_490_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_490_valid <= _GEN_15852;
      end
    end else begin
      btb_490_valid <= _GEN_15852;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_490_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ea == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_490_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_490_tag <= _GEN_6634;
      end
    end else begin
      btb_490_tag <= _GEN_6634;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_490_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ea == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_490_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_490_target_address <= _GEN_12224;
      end
    end else begin
      btb_490_target_address <= _GEN_12224;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_490_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ea == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_490_bht <= 2'h1;
        end else begin
          btb_490_bht <= 2'h0;
        end
      end else begin
        btb_490_bht <= _GEN_12226;
      end
    end else begin
      btb_490_bht <= _GEN_12226;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_491_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_491_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_491_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_491_valid <= _GEN_15853;
      end
    end else begin
      btb_491_valid <= _GEN_15853;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_491_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1eb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_491_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_491_tag <= _GEN_6635;
      end
    end else begin
      btb_491_tag <= _GEN_6635;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_491_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1eb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_491_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_491_target_address <= _GEN_12227;
      end
    end else begin
      btb_491_target_address <= _GEN_12227;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_491_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1eb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_491_bht <= 2'h1;
        end else begin
          btb_491_bht <= 2'h0;
        end
      end else begin
        btb_491_bht <= _GEN_12229;
      end
    end else begin
      btb_491_bht <= _GEN_12229;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_492_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_492_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_492_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_492_valid <= _GEN_15854;
      end
    end else begin
      btb_492_valid <= _GEN_15854;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_492_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ec == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_492_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_492_tag <= _GEN_6636;
      end
    end else begin
      btb_492_tag <= _GEN_6636;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_492_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ec == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_492_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_492_target_address <= _GEN_12230;
      end
    end else begin
      btb_492_target_address <= _GEN_12230;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_492_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ec == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_492_bht <= 2'h1;
        end else begin
          btb_492_bht <= 2'h0;
        end
      end else begin
        btb_492_bht <= _GEN_12232;
      end
    end else begin
      btb_492_bht <= _GEN_12232;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_493_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_493_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_493_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_493_valid <= _GEN_15855;
      end
    end else begin
      btb_493_valid <= _GEN_15855;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_493_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ed == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_493_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_493_tag <= _GEN_6637;
      end
    end else begin
      btb_493_tag <= _GEN_6637;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_493_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ed == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_493_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_493_target_address <= _GEN_12233;
      end
    end else begin
      btb_493_target_address <= _GEN_12233;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_493_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ed == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_493_bht <= 2'h1;
        end else begin
          btb_493_bht <= 2'h0;
        end
      end else begin
        btb_493_bht <= _GEN_12235;
      end
    end else begin
      btb_493_bht <= _GEN_12235;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_494_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_494_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_494_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_494_valid <= _GEN_15856;
      end
    end else begin
      btb_494_valid <= _GEN_15856;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_494_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ee == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_494_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_494_tag <= _GEN_6638;
      end
    end else begin
      btb_494_tag <= _GEN_6638;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_494_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ee == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_494_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_494_target_address <= _GEN_12236;
      end
    end else begin
      btb_494_target_address <= _GEN_12236;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_494_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ee == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_494_bht <= 2'h1;
        end else begin
          btb_494_bht <= 2'h0;
        end
      end else begin
        btb_494_bht <= _GEN_12238;
      end
    end else begin
      btb_494_bht <= _GEN_12238;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_495_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_495_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_495_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_495_valid <= _GEN_15857;
      end
    end else begin
      btb_495_valid <= _GEN_15857;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_495_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ef == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_495_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_495_tag <= _GEN_6639;
      end
    end else begin
      btb_495_tag <= _GEN_6639;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_495_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ef == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_495_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_495_target_address <= _GEN_12239;
      end
    end else begin
      btb_495_target_address <= _GEN_12239;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_495_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ef == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_495_bht <= 2'h1;
        end else begin
          btb_495_bht <= 2'h0;
        end
      end else begin
        btb_495_bht <= _GEN_12241;
      end
    end else begin
      btb_495_bht <= _GEN_12241;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_496_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_496_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_496_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_496_valid <= _GEN_15858;
      end
    end else begin
      btb_496_valid <= _GEN_15858;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_496_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f0 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_496_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_496_tag <= _GEN_6640;
      end
    end else begin
      btb_496_tag <= _GEN_6640;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_496_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f0 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_496_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_496_target_address <= _GEN_12242;
      end
    end else begin
      btb_496_target_address <= _GEN_12242;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_496_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f0 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_496_bht <= 2'h1;
        end else begin
          btb_496_bht <= 2'h0;
        end
      end else begin
        btb_496_bht <= _GEN_12244;
      end
    end else begin
      btb_496_bht <= _GEN_12244;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_497_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_497_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_497_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_497_valid <= _GEN_15859;
      end
    end else begin
      btb_497_valid <= _GEN_15859;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_497_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f1 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_497_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_497_tag <= _GEN_6641;
      end
    end else begin
      btb_497_tag <= _GEN_6641;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_497_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f1 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_497_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_497_target_address <= _GEN_12245;
      end
    end else begin
      btb_497_target_address <= _GEN_12245;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_497_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f1 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_497_bht <= 2'h1;
        end else begin
          btb_497_bht <= 2'h0;
        end
      end else begin
        btb_497_bht <= _GEN_12247;
      end
    end else begin
      btb_497_bht <= _GEN_12247;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_498_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_498_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_498_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_498_valid <= _GEN_15860;
      end
    end else begin
      btb_498_valid <= _GEN_15860;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_498_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f2 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_498_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_498_tag <= _GEN_6642;
      end
    end else begin
      btb_498_tag <= _GEN_6642;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_498_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f2 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_498_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_498_target_address <= _GEN_12248;
      end
    end else begin
      btb_498_target_address <= _GEN_12248;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_498_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f2 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_498_bht <= 2'h1;
        end else begin
          btb_498_bht <= 2'h0;
        end
      end else begin
        btb_498_bht <= _GEN_12250;
      end
    end else begin
      btb_498_bht <= _GEN_12250;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_499_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_499_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_499_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_499_valid <= _GEN_15861;
      end
    end else begin
      btb_499_valid <= _GEN_15861;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_499_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f3 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_499_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_499_tag <= _GEN_6643;
      end
    end else begin
      btb_499_tag <= _GEN_6643;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_499_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f3 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_499_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_499_target_address <= _GEN_12251;
      end
    end else begin
      btb_499_target_address <= _GEN_12251;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_499_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f3 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_499_bht <= 2'h1;
        end else begin
          btb_499_bht <= 2'h0;
        end
      end else begin
        btb_499_bht <= _GEN_12253;
      end
    end else begin
      btb_499_bht <= _GEN_12253;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_500_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_500_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_500_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_500_valid <= _GEN_15862;
      end
    end else begin
      btb_500_valid <= _GEN_15862;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_500_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f4 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_500_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_500_tag <= _GEN_6644;
      end
    end else begin
      btb_500_tag <= _GEN_6644;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_500_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f4 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_500_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_500_target_address <= _GEN_12254;
      end
    end else begin
      btb_500_target_address <= _GEN_12254;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_500_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f4 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_500_bht <= 2'h1;
        end else begin
          btb_500_bht <= 2'h0;
        end
      end else begin
        btb_500_bht <= _GEN_12256;
      end
    end else begin
      btb_500_bht <= _GEN_12256;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_501_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_501_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_501_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_501_valid <= _GEN_15863;
      end
    end else begin
      btb_501_valid <= _GEN_15863;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_501_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f5 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_501_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_501_tag <= _GEN_6645;
      end
    end else begin
      btb_501_tag <= _GEN_6645;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_501_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f5 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_501_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_501_target_address <= _GEN_12257;
      end
    end else begin
      btb_501_target_address <= _GEN_12257;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_501_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f5 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_501_bht <= 2'h1;
        end else begin
          btb_501_bht <= 2'h0;
        end
      end else begin
        btb_501_bht <= _GEN_12259;
      end
    end else begin
      btb_501_bht <= _GEN_12259;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_502_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_502_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_502_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_502_valid <= _GEN_15864;
      end
    end else begin
      btb_502_valid <= _GEN_15864;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_502_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f6 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_502_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_502_tag <= _GEN_6646;
      end
    end else begin
      btb_502_tag <= _GEN_6646;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_502_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f6 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_502_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_502_target_address <= _GEN_12260;
      end
    end else begin
      btb_502_target_address <= _GEN_12260;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_502_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f6 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_502_bht <= 2'h1;
        end else begin
          btb_502_bht <= 2'h0;
        end
      end else begin
        btb_502_bht <= _GEN_12262;
      end
    end else begin
      btb_502_bht <= _GEN_12262;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_503_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_503_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_503_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_503_valid <= _GEN_15865;
      end
    end else begin
      btb_503_valid <= _GEN_15865;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_503_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f7 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_503_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_503_tag <= _GEN_6647;
      end
    end else begin
      btb_503_tag <= _GEN_6647;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_503_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f7 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_503_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_503_target_address <= _GEN_12263;
      end
    end else begin
      btb_503_target_address <= _GEN_12263;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_503_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f7 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_503_bht <= 2'h1;
        end else begin
          btb_503_bht <= 2'h0;
        end
      end else begin
        btb_503_bht <= _GEN_12265;
      end
    end else begin
      btb_503_bht <= _GEN_12265;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_504_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_504_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_504_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_504_valid <= _GEN_15866;
      end
    end else begin
      btb_504_valid <= _GEN_15866;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_504_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f8 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_504_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_504_tag <= _GEN_6648;
      end
    end else begin
      btb_504_tag <= _GEN_6648;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_504_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f8 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_504_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_504_target_address <= _GEN_12266;
      end
    end else begin
      btb_504_target_address <= _GEN_12266;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_504_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f8 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_504_bht <= 2'h1;
        end else begin
          btb_504_bht <= 2'h0;
        end
      end else begin
        btb_504_bht <= _GEN_12268;
      end
    end else begin
      btb_504_bht <= _GEN_12268;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_505_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_505_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_505_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_505_valid <= _GEN_15867;
      end
    end else begin
      btb_505_valid <= _GEN_15867;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_505_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f9 == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_505_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_505_tag <= _GEN_6649;
      end
    end else begin
      btb_505_tag <= _GEN_6649;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_505_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f9 == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_505_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_505_target_address <= _GEN_12269;
      end
    end else begin
      btb_505_target_address <= _GEN_12269;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_505_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1f9 == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_505_bht <= 2'h1;
        end else begin
          btb_505_bht <= 2'h0;
        end
      end else begin
        btb_505_bht <= _GEN_12271;
      end
    end else begin
      btb_505_bht <= _GEN_12271;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_506_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_506_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_506_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_506_valid <= _GEN_15868;
      end
    end else begin
      btb_506_valid <= _GEN_15868;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_506_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fa == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_506_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_506_tag <= _GEN_6650;
      end
    end else begin
      btb_506_tag <= _GEN_6650;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_506_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fa == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_506_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_506_target_address <= _GEN_12272;
      end
    end else begin
      btb_506_target_address <= _GEN_12272;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_506_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fa == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_506_bht <= 2'h1;
        end else begin
          btb_506_bht <= 2'h0;
        end
      end else begin
        btb_506_bht <= _GEN_12274;
      end
    end else begin
      btb_506_bht <= _GEN_12274;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_507_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_507_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_507_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_507_valid <= _GEN_15869;
      end
    end else begin
      btb_507_valid <= _GEN_15869;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_507_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fb == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_507_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_507_tag <= _GEN_6651;
      end
    end else begin
      btb_507_tag <= _GEN_6651;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_507_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fb == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_507_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_507_target_address <= _GEN_12275;
      end
    end else begin
      btb_507_target_address <= _GEN_12275;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_507_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fb == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_507_bht <= 2'h1;
        end else begin
          btb_507_bht <= 2'h0;
        end
      end else begin
        btb_507_bht <= _GEN_12277;
      end
    end else begin
      btb_507_bht <= _GEN_12277;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_508_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_508_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_508_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_508_valid <= _GEN_15870;
      end
    end else begin
      btb_508_valid <= _GEN_15870;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_508_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fc == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_508_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_508_tag <= _GEN_6652;
      end
    end else begin
      btb_508_tag <= _GEN_6652;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_508_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fc == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_508_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_508_target_address <= _GEN_12278;
      end
    end else begin
      btb_508_target_address <= _GEN_12278;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_508_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fc == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_508_bht <= 2'h1;
        end else begin
          btb_508_bht <= 2'h0;
        end
      end else begin
        btb_508_bht <= _GEN_12280;
      end
    end else begin
      btb_508_bht <= _GEN_12280;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_509_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_509_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_509_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_509_valid <= _GEN_15871;
      end
    end else begin
      btb_509_valid <= _GEN_15871;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_509_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fd == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_509_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_509_tag <= _GEN_6653;
      end
    end else begin
      btb_509_tag <= _GEN_6653;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_509_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fd == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_509_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_509_target_address <= _GEN_12281;
      end
    end else begin
      btb_509_target_address <= _GEN_12281;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_509_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fd == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_509_bht <= 2'h1;
        end else begin
          btb_509_bht <= 2'h0;
        end
      end else begin
        btb_509_bht <= _GEN_12283;
      end
    end else begin
      btb_509_bht <= _GEN_12283;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_510_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_510_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_510_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_510_valid <= _GEN_15872;
      end
    end else begin
      btb_510_valid <= _GEN_15872;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_510_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fe == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_510_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_510_tag <= _GEN_6654;
      end
    end else begin
      btb_510_tag <= _GEN_6654;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_510_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fe == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_510_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_510_target_address <= _GEN_12284;
      end
    end else begin
      btb_510_target_address <= _GEN_12284;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_510_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1fe == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_510_bht <= 2'h1;
        end else begin
          btb_510_bht <= 2'h0;
        end
      end else begin
        btb_510_bht <= _GEN_12286;
      end
    end else begin
      btb_510_bht <= _GEN_12286;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_511_valid <= 1'h0; // @[branch_predictor.scala 30:22]
    end else if (io_i_branch_presolve_pack_valid) begin // @[branch_predictor.scala 109:42]
      if (btb_511_tag == io_i_branch_presolve_pack_pc[12:3]) begin // @[branch_predictor.scala 111:68]
        btb_511_valid <= 1'h0; // @[branch_predictor.scala 112:30]
      end else begin
        btb_511_valid <= _GEN_15873;
      end
    end else begin
      btb_511_valid <= _GEN_15873;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_511_tag <= 10'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ff == btb_victim_ptr) begin // @[branch_predictor.scala 100:33]
        btb_511_tag <= io_i_branch_resolve_pack_pc[12:3]; // @[branch_predictor.scala 100:33]
      end else begin
        btb_511_tag <= _GEN_6655;
      end
    end else begin
      btb_511_tag <= _GEN_6655;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_511_target_address <= 64'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ff == btb_victim_ptr) begin // @[branch_predictor.scala 101:44]
        btb_511_target_address <= io_i_branch_resolve_pack_target; // @[branch_predictor.scala 101:44]
      end else begin
        btb_511_target_address <= _GEN_12287;
      end
    end else begin
      btb_511_target_address <= _GEN_12287;
    end
    if (reset) begin // @[branch_predictor.scala 30:22]
      btb_511_bht <= 2'h0; // @[branch_predictor.scala 30:22]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      if (9'h1ff == btb_victim_ptr) begin // @[branch_predictor.scala 104:33]
        if (io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 68:39]
          btb_511_bht <= 2'h1;
        end else begin
          btb_511_bht <= 2'h0;
        end
      end else begin
        btb_511_bht <= _GEN_12289;
      end
    end else begin
      btb_511_bht <= _GEN_12289;
    end
    if (reset) begin // @[branch_predictor.scala 32:33]
      btb_victim_ptr <= 9'h0; // @[branch_predictor.scala 32:33]
    end else if (_T_1027 & ~entry_found) begin // @[branch_predictor.scala 98:103]
      btb_victim_ptr <= _btb_victim_ptr_T_1; // @[branch_predictor.scala 107:24]
    end else if (io_i_branch_resolve_pack_valid & ~io_i_branch_resolve_pack_prediction_valid &
      io_i_branch_resolve_pack_taken) begin // @[branch_predictor.scala 62:121]
      btb_victim_ptr <= _btb_victim_ptr_T_1; // @[branch_predictor.scala 71:24]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_0_tag = _RAND_1[9:0];
  _RAND_2 = {2{`RANDOM}};
  btb_0_target_address = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  btb_0_bht = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  btb_1_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  btb_1_tag = _RAND_5[9:0];
  _RAND_6 = {2{`RANDOM}};
  btb_1_target_address = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  btb_1_bht = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  btb_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  btb_2_tag = _RAND_9[9:0];
  _RAND_10 = {2{`RANDOM}};
  btb_2_target_address = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  btb_2_bht = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  btb_3_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btb_3_tag = _RAND_13[9:0];
  _RAND_14 = {2{`RANDOM}};
  btb_3_target_address = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  btb_3_bht = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  btb_4_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  btb_4_tag = _RAND_17[9:0];
  _RAND_18 = {2{`RANDOM}};
  btb_4_target_address = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  btb_4_bht = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  btb_5_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  btb_5_tag = _RAND_21[9:0];
  _RAND_22 = {2{`RANDOM}};
  btb_5_target_address = _RAND_22[63:0];
  _RAND_23 = {1{`RANDOM}};
  btb_5_bht = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  btb_6_valid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  btb_6_tag = _RAND_25[9:0];
  _RAND_26 = {2{`RANDOM}};
  btb_6_target_address = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  btb_6_bht = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  btb_7_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  btb_7_tag = _RAND_29[9:0];
  _RAND_30 = {2{`RANDOM}};
  btb_7_target_address = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  btb_7_bht = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  btb_8_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  btb_8_tag = _RAND_33[9:0];
  _RAND_34 = {2{`RANDOM}};
  btb_8_target_address = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  btb_8_bht = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  btb_9_valid = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  btb_9_tag = _RAND_37[9:0];
  _RAND_38 = {2{`RANDOM}};
  btb_9_target_address = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  btb_9_bht = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  btb_10_valid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  btb_10_tag = _RAND_41[9:0];
  _RAND_42 = {2{`RANDOM}};
  btb_10_target_address = _RAND_42[63:0];
  _RAND_43 = {1{`RANDOM}};
  btb_10_bht = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  btb_11_valid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  btb_11_tag = _RAND_45[9:0];
  _RAND_46 = {2{`RANDOM}};
  btb_11_target_address = _RAND_46[63:0];
  _RAND_47 = {1{`RANDOM}};
  btb_11_bht = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  btb_12_valid = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  btb_12_tag = _RAND_49[9:0];
  _RAND_50 = {2{`RANDOM}};
  btb_12_target_address = _RAND_50[63:0];
  _RAND_51 = {1{`RANDOM}};
  btb_12_bht = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  btb_13_valid = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  btb_13_tag = _RAND_53[9:0];
  _RAND_54 = {2{`RANDOM}};
  btb_13_target_address = _RAND_54[63:0];
  _RAND_55 = {1{`RANDOM}};
  btb_13_bht = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  btb_14_valid = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  btb_14_tag = _RAND_57[9:0];
  _RAND_58 = {2{`RANDOM}};
  btb_14_target_address = _RAND_58[63:0];
  _RAND_59 = {1{`RANDOM}};
  btb_14_bht = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  btb_15_valid = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  btb_15_tag = _RAND_61[9:0];
  _RAND_62 = {2{`RANDOM}};
  btb_15_target_address = _RAND_62[63:0];
  _RAND_63 = {1{`RANDOM}};
  btb_15_bht = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  btb_16_valid = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  btb_16_tag = _RAND_65[9:0];
  _RAND_66 = {2{`RANDOM}};
  btb_16_target_address = _RAND_66[63:0];
  _RAND_67 = {1{`RANDOM}};
  btb_16_bht = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  btb_17_valid = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  btb_17_tag = _RAND_69[9:0];
  _RAND_70 = {2{`RANDOM}};
  btb_17_target_address = _RAND_70[63:0];
  _RAND_71 = {1{`RANDOM}};
  btb_17_bht = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  btb_18_valid = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  btb_18_tag = _RAND_73[9:0];
  _RAND_74 = {2{`RANDOM}};
  btb_18_target_address = _RAND_74[63:0];
  _RAND_75 = {1{`RANDOM}};
  btb_18_bht = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  btb_19_valid = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  btb_19_tag = _RAND_77[9:0];
  _RAND_78 = {2{`RANDOM}};
  btb_19_target_address = _RAND_78[63:0];
  _RAND_79 = {1{`RANDOM}};
  btb_19_bht = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  btb_20_valid = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  btb_20_tag = _RAND_81[9:0];
  _RAND_82 = {2{`RANDOM}};
  btb_20_target_address = _RAND_82[63:0];
  _RAND_83 = {1{`RANDOM}};
  btb_20_bht = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  btb_21_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  btb_21_tag = _RAND_85[9:0];
  _RAND_86 = {2{`RANDOM}};
  btb_21_target_address = _RAND_86[63:0];
  _RAND_87 = {1{`RANDOM}};
  btb_21_bht = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  btb_22_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  btb_22_tag = _RAND_89[9:0];
  _RAND_90 = {2{`RANDOM}};
  btb_22_target_address = _RAND_90[63:0];
  _RAND_91 = {1{`RANDOM}};
  btb_22_bht = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  btb_23_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  btb_23_tag = _RAND_93[9:0];
  _RAND_94 = {2{`RANDOM}};
  btb_23_target_address = _RAND_94[63:0];
  _RAND_95 = {1{`RANDOM}};
  btb_23_bht = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  btb_24_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  btb_24_tag = _RAND_97[9:0];
  _RAND_98 = {2{`RANDOM}};
  btb_24_target_address = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  btb_24_bht = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  btb_25_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  btb_25_tag = _RAND_101[9:0];
  _RAND_102 = {2{`RANDOM}};
  btb_25_target_address = _RAND_102[63:0];
  _RAND_103 = {1{`RANDOM}};
  btb_25_bht = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  btb_26_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  btb_26_tag = _RAND_105[9:0];
  _RAND_106 = {2{`RANDOM}};
  btb_26_target_address = _RAND_106[63:0];
  _RAND_107 = {1{`RANDOM}};
  btb_26_bht = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  btb_27_valid = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  btb_27_tag = _RAND_109[9:0];
  _RAND_110 = {2{`RANDOM}};
  btb_27_target_address = _RAND_110[63:0];
  _RAND_111 = {1{`RANDOM}};
  btb_27_bht = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  btb_28_valid = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  btb_28_tag = _RAND_113[9:0];
  _RAND_114 = {2{`RANDOM}};
  btb_28_target_address = _RAND_114[63:0];
  _RAND_115 = {1{`RANDOM}};
  btb_28_bht = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  btb_29_valid = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  btb_29_tag = _RAND_117[9:0];
  _RAND_118 = {2{`RANDOM}};
  btb_29_target_address = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  btb_29_bht = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  btb_30_valid = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  btb_30_tag = _RAND_121[9:0];
  _RAND_122 = {2{`RANDOM}};
  btb_30_target_address = _RAND_122[63:0];
  _RAND_123 = {1{`RANDOM}};
  btb_30_bht = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  btb_31_valid = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  btb_31_tag = _RAND_125[9:0];
  _RAND_126 = {2{`RANDOM}};
  btb_31_target_address = _RAND_126[63:0];
  _RAND_127 = {1{`RANDOM}};
  btb_31_bht = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  btb_32_valid = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  btb_32_tag = _RAND_129[9:0];
  _RAND_130 = {2{`RANDOM}};
  btb_32_target_address = _RAND_130[63:0];
  _RAND_131 = {1{`RANDOM}};
  btb_32_bht = _RAND_131[1:0];
  _RAND_132 = {1{`RANDOM}};
  btb_33_valid = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  btb_33_tag = _RAND_133[9:0];
  _RAND_134 = {2{`RANDOM}};
  btb_33_target_address = _RAND_134[63:0];
  _RAND_135 = {1{`RANDOM}};
  btb_33_bht = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  btb_34_valid = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  btb_34_tag = _RAND_137[9:0];
  _RAND_138 = {2{`RANDOM}};
  btb_34_target_address = _RAND_138[63:0];
  _RAND_139 = {1{`RANDOM}};
  btb_34_bht = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  btb_35_valid = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  btb_35_tag = _RAND_141[9:0];
  _RAND_142 = {2{`RANDOM}};
  btb_35_target_address = _RAND_142[63:0];
  _RAND_143 = {1{`RANDOM}};
  btb_35_bht = _RAND_143[1:0];
  _RAND_144 = {1{`RANDOM}};
  btb_36_valid = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  btb_36_tag = _RAND_145[9:0];
  _RAND_146 = {2{`RANDOM}};
  btb_36_target_address = _RAND_146[63:0];
  _RAND_147 = {1{`RANDOM}};
  btb_36_bht = _RAND_147[1:0];
  _RAND_148 = {1{`RANDOM}};
  btb_37_valid = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  btb_37_tag = _RAND_149[9:0];
  _RAND_150 = {2{`RANDOM}};
  btb_37_target_address = _RAND_150[63:0];
  _RAND_151 = {1{`RANDOM}};
  btb_37_bht = _RAND_151[1:0];
  _RAND_152 = {1{`RANDOM}};
  btb_38_valid = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  btb_38_tag = _RAND_153[9:0];
  _RAND_154 = {2{`RANDOM}};
  btb_38_target_address = _RAND_154[63:0];
  _RAND_155 = {1{`RANDOM}};
  btb_38_bht = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  btb_39_valid = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  btb_39_tag = _RAND_157[9:0];
  _RAND_158 = {2{`RANDOM}};
  btb_39_target_address = _RAND_158[63:0];
  _RAND_159 = {1{`RANDOM}};
  btb_39_bht = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  btb_40_valid = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  btb_40_tag = _RAND_161[9:0];
  _RAND_162 = {2{`RANDOM}};
  btb_40_target_address = _RAND_162[63:0];
  _RAND_163 = {1{`RANDOM}};
  btb_40_bht = _RAND_163[1:0];
  _RAND_164 = {1{`RANDOM}};
  btb_41_valid = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  btb_41_tag = _RAND_165[9:0];
  _RAND_166 = {2{`RANDOM}};
  btb_41_target_address = _RAND_166[63:0];
  _RAND_167 = {1{`RANDOM}};
  btb_41_bht = _RAND_167[1:0];
  _RAND_168 = {1{`RANDOM}};
  btb_42_valid = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  btb_42_tag = _RAND_169[9:0];
  _RAND_170 = {2{`RANDOM}};
  btb_42_target_address = _RAND_170[63:0];
  _RAND_171 = {1{`RANDOM}};
  btb_42_bht = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  btb_43_valid = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  btb_43_tag = _RAND_173[9:0];
  _RAND_174 = {2{`RANDOM}};
  btb_43_target_address = _RAND_174[63:0];
  _RAND_175 = {1{`RANDOM}};
  btb_43_bht = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  btb_44_valid = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  btb_44_tag = _RAND_177[9:0];
  _RAND_178 = {2{`RANDOM}};
  btb_44_target_address = _RAND_178[63:0];
  _RAND_179 = {1{`RANDOM}};
  btb_44_bht = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  btb_45_valid = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  btb_45_tag = _RAND_181[9:0];
  _RAND_182 = {2{`RANDOM}};
  btb_45_target_address = _RAND_182[63:0];
  _RAND_183 = {1{`RANDOM}};
  btb_45_bht = _RAND_183[1:0];
  _RAND_184 = {1{`RANDOM}};
  btb_46_valid = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  btb_46_tag = _RAND_185[9:0];
  _RAND_186 = {2{`RANDOM}};
  btb_46_target_address = _RAND_186[63:0];
  _RAND_187 = {1{`RANDOM}};
  btb_46_bht = _RAND_187[1:0];
  _RAND_188 = {1{`RANDOM}};
  btb_47_valid = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  btb_47_tag = _RAND_189[9:0];
  _RAND_190 = {2{`RANDOM}};
  btb_47_target_address = _RAND_190[63:0];
  _RAND_191 = {1{`RANDOM}};
  btb_47_bht = _RAND_191[1:0];
  _RAND_192 = {1{`RANDOM}};
  btb_48_valid = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  btb_48_tag = _RAND_193[9:0];
  _RAND_194 = {2{`RANDOM}};
  btb_48_target_address = _RAND_194[63:0];
  _RAND_195 = {1{`RANDOM}};
  btb_48_bht = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  btb_49_valid = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  btb_49_tag = _RAND_197[9:0];
  _RAND_198 = {2{`RANDOM}};
  btb_49_target_address = _RAND_198[63:0];
  _RAND_199 = {1{`RANDOM}};
  btb_49_bht = _RAND_199[1:0];
  _RAND_200 = {1{`RANDOM}};
  btb_50_valid = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  btb_50_tag = _RAND_201[9:0];
  _RAND_202 = {2{`RANDOM}};
  btb_50_target_address = _RAND_202[63:0];
  _RAND_203 = {1{`RANDOM}};
  btb_50_bht = _RAND_203[1:0];
  _RAND_204 = {1{`RANDOM}};
  btb_51_valid = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  btb_51_tag = _RAND_205[9:0];
  _RAND_206 = {2{`RANDOM}};
  btb_51_target_address = _RAND_206[63:0];
  _RAND_207 = {1{`RANDOM}};
  btb_51_bht = _RAND_207[1:0];
  _RAND_208 = {1{`RANDOM}};
  btb_52_valid = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  btb_52_tag = _RAND_209[9:0];
  _RAND_210 = {2{`RANDOM}};
  btb_52_target_address = _RAND_210[63:0];
  _RAND_211 = {1{`RANDOM}};
  btb_52_bht = _RAND_211[1:0];
  _RAND_212 = {1{`RANDOM}};
  btb_53_valid = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  btb_53_tag = _RAND_213[9:0];
  _RAND_214 = {2{`RANDOM}};
  btb_53_target_address = _RAND_214[63:0];
  _RAND_215 = {1{`RANDOM}};
  btb_53_bht = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  btb_54_valid = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  btb_54_tag = _RAND_217[9:0];
  _RAND_218 = {2{`RANDOM}};
  btb_54_target_address = _RAND_218[63:0];
  _RAND_219 = {1{`RANDOM}};
  btb_54_bht = _RAND_219[1:0];
  _RAND_220 = {1{`RANDOM}};
  btb_55_valid = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  btb_55_tag = _RAND_221[9:0];
  _RAND_222 = {2{`RANDOM}};
  btb_55_target_address = _RAND_222[63:0];
  _RAND_223 = {1{`RANDOM}};
  btb_55_bht = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  btb_56_valid = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  btb_56_tag = _RAND_225[9:0];
  _RAND_226 = {2{`RANDOM}};
  btb_56_target_address = _RAND_226[63:0];
  _RAND_227 = {1{`RANDOM}};
  btb_56_bht = _RAND_227[1:0];
  _RAND_228 = {1{`RANDOM}};
  btb_57_valid = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  btb_57_tag = _RAND_229[9:0];
  _RAND_230 = {2{`RANDOM}};
  btb_57_target_address = _RAND_230[63:0];
  _RAND_231 = {1{`RANDOM}};
  btb_57_bht = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  btb_58_valid = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  btb_58_tag = _RAND_233[9:0];
  _RAND_234 = {2{`RANDOM}};
  btb_58_target_address = _RAND_234[63:0];
  _RAND_235 = {1{`RANDOM}};
  btb_58_bht = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  btb_59_valid = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  btb_59_tag = _RAND_237[9:0];
  _RAND_238 = {2{`RANDOM}};
  btb_59_target_address = _RAND_238[63:0];
  _RAND_239 = {1{`RANDOM}};
  btb_59_bht = _RAND_239[1:0];
  _RAND_240 = {1{`RANDOM}};
  btb_60_valid = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  btb_60_tag = _RAND_241[9:0];
  _RAND_242 = {2{`RANDOM}};
  btb_60_target_address = _RAND_242[63:0];
  _RAND_243 = {1{`RANDOM}};
  btb_60_bht = _RAND_243[1:0];
  _RAND_244 = {1{`RANDOM}};
  btb_61_valid = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  btb_61_tag = _RAND_245[9:0];
  _RAND_246 = {2{`RANDOM}};
  btb_61_target_address = _RAND_246[63:0];
  _RAND_247 = {1{`RANDOM}};
  btb_61_bht = _RAND_247[1:0];
  _RAND_248 = {1{`RANDOM}};
  btb_62_valid = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  btb_62_tag = _RAND_249[9:0];
  _RAND_250 = {2{`RANDOM}};
  btb_62_target_address = _RAND_250[63:0];
  _RAND_251 = {1{`RANDOM}};
  btb_62_bht = _RAND_251[1:0];
  _RAND_252 = {1{`RANDOM}};
  btb_63_valid = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  btb_63_tag = _RAND_253[9:0];
  _RAND_254 = {2{`RANDOM}};
  btb_63_target_address = _RAND_254[63:0];
  _RAND_255 = {1{`RANDOM}};
  btb_63_bht = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  btb_64_valid = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  btb_64_tag = _RAND_257[9:0];
  _RAND_258 = {2{`RANDOM}};
  btb_64_target_address = _RAND_258[63:0];
  _RAND_259 = {1{`RANDOM}};
  btb_64_bht = _RAND_259[1:0];
  _RAND_260 = {1{`RANDOM}};
  btb_65_valid = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  btb_65_tag = _RAND_261[9:0];
  _RAND_262 = {2{`RANDOM}};
  btb_65_target_address = _RAND_262[63:0];
  _RAND_263 = {1{`RANDOM}};
  btb_65_bht = _RAND_263[1:0];
  _RAND_264 = {1{`RANDOM}};
  btb_66_valid = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  btb_66_tag = _RAND_265[9:0];
  _RAND_266 = {2{`RANDOM}};
  btb_66_target_address = _RAND_266[63:0];
  _RAND_267 = {1{`RANDOM}};
  btb_66_bht = _RAND_267[1:0];
  _RAND_268 = {1{`RANDOM}};
  btb_67_valid = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  btb_67_tag = _RAND_269[9:0];
  _RAND_270 = {2{`RANDOM}};
  btb_67_target_address = _RAND_270[63:0];
  _RAND_271 = {1{`RANDOM}};
  btb_67_bht = _RAND_271[1:0];
  _RAND_272 = {1{`RANDOM}};
  btb_68_valid = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  btb_68_tag = _RAND_273[9:0];
  _RAND_274 = {2{`RANDOM}};
  btb_68_target_address = _RAND_274[63:0];
  _RAND_275 = {1{`RANDOM}};
  btb_68_bht = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  btb_69_valid = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  btb_69_tag = _RAND_277[9:0];
  _RAND_278 = {2{`RANDOM}};
  btb_69_target_address = _RAND_278[63:0];
  _RAND_279 = {1{`RANDOM}};
  btb_69_bht = _RAND_279[1:0];
  _RAND_280 = {1{`RANDOM}};
  btb_70_valid = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  btb_70_tag = _RAND_281[9:0];
  _RAND_282 = {2{`RANDOM}};
  btb_70_target_address = _RAND_282[63:0];
  _RAND_283 = {1{`RANDOM}};
  btb_70_bht = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  btb_71_valid = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  btb_71_tag = _RAND_285[9:0];
  _RAND_286 = {2{`RANDOM}};
  btb_71_target_address = _RAND_286[63:0];
  _RAND_287 = {1{`RANDOM}};
  btb_71_bht = _RAND_287[1:0];
  _RAND_288 = {1{`RANDOM}};
  btb_72_valid = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  btb_72_tag = _RAND_289[9:0];
  _RAND_290 = {2{`RANDOM}};
  btb_72_target_address = _RAND_290[63:0];
  _RAND_291 = {1{`RANDOM}};
  btb_72_bht = _RAND_291[1:0];
  _RAND_292 = {1{`RANDOM}};
  btb_73_valid = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  btb_73_tag = _RAND_293[9:0];
  _RAND_294 = {2{`RANDOM}};
  btb_73_target_address = _RAND_294[63:0];
  _RAND_295 = {1{`RANDOM}};
  btb_73_bht = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  btb_74_valid = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  btb_74_tag = _RAND_297[9:0];
  _RAND_298 = {2{`RANDOM}};
  btb_74_target_address = _RAND_298[63:0];
  _RAND_299 = {1{`RANDOM}};
  btb_74_bht = _RAND_299[1:0];
  _RAND_300 = {1{`RANDOM}};
  btb_75_valid = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  btb_75_tag = _RAND_301[9:0];
  _RAND_302 = {2{`RANDOM}};
  btb_75_target_address = _RAND_302[63:0];
  _RAND_303 = {1{`RANDOM}};
  btb_75_bht = _RAND_303[1:0];
  _RAND_304 = {1{`RANDOM}};
  btb_76_valid = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  btb_76_tag = _RAND_305[9:0];
  _RAND_306 = {2{`RANDOM}};
  btb_76_target_address = _RAND_306[63:0];
  _RAND_307 = {1{`RANDOM}};
  btb_76_bht = _RAND_307[1:0];
  _RAND_308 = {1{`RANDOM}};
  btb_77_valid = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  btb_77_tag = _RAND_309[9:0];
  _RAND_310 = {2{`RANDOM}};
  btb_77_target_address = _RAND_310[63:0];
  _RAND_311 = {1{`RANDOM}};
  btb_77_bht = _RAND_311[1:0];
  _RAND_312 = {1{`RANDOM}};
  btb_78_valid = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  btb_78_tag = _RAND_313[9:0];
  _RAND_314 = {2{`RANDOM}};
  btb_78_target_address = _RAND_314[63:0];
  _RAND_315 = {1{`RANDOM}};
  btb_78_bht = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  btb_79_valid = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  btb_79_tag = _RAND_317[9:0];
  _RAND_318 = {2{`RANDOM}};
  btb_79_target_address = _RAND_318[63:0];
  _RAND_319 = {1{`RANDOM}};
  btb_79_bht = _RAND_319[1:0];
  _RAND_320 = {1{`RANDOM}};
  btb_80_valid = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  btb_80_tag = _RAND_321[9:0];
  _RAND_322 = {2{`RANDOM}};
  btb_80_target_address = _RAND_322[63:0];
  _RAND_323 = {1{`RANDOM}};
  btb_80_bht = _RAND_323[1:0];
  _RAND_324 = {1{`RANDOM}};
  btb_81_valid = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  btb_81_tag = _RAND_325[9:0];
  _RAND_326 = {2{`RANDOM}};
  btb_81_target_address = _RAND_326[63:0];
  _RAND_327 = {1{`RANDOM}};
  btb_81_bht = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  btb_82_valid = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  btb_82_tag = _RAND_329[9:0];
  _RAND_330 = {2{`RANDOM}};
  btb_82_target_address = _RAND_330[63:0];
  _RAND_331 = {1{`RANDOM}};
  btb_82_bht = _RAND_331[1:0];
  _RAND_332 = {1{`RANDOM}};
  btb_83_valid = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  btb_83_tag = _RAND_333[9:0];
  _RAND_334 = {2{`RANDOM}};
  btb_83_target_address = _RAND_334[63:0];
  _RAND_335 = {1{`RANDOM}};
  btb_83_bht = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  btb_84_valid = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  btb_84_tag = _RAND_337[9:0];
  _RAND_338 = {2{`RANDOM}};
  btb_84_target_address = _RAND_338[63:0];
  _RAND_339 = {1{`RANDOM}};
  btb_84_bht = _RAND_339[1:0];
  _RAND_340 = {1{`RANDOM}};
  btb_85_valid = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  btb_85_tag = _RAND_341[9:0];
  _RAND_342 = {2{`RANDOM}};
  btb_85_target_address = _RAND_342[63:0];
  _RAND_343 = {1{`RANDOM}};
  btb_85_bht = _RAND_343[1:0];
  _RAND_344 = {1{`RANDOM}};
  btb_86_valid = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  btb_86_tag = _RAND_345[9:0];
  _RAND_346 = {2{`RANDOM}};
  btb_86_target_address = _RAND_346[63:0];
  _RAND_347 = {1{`RANDOM}};
  btb_86_bht = _RAND_347[1:0];
  _RAND_348 = {1{`RANDOM}};
  btb_87_valid = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  btb_87_tag = _RAND_349[9:0];
  _RAND_350 = {2{`RANDOM}};
  btb_87_target_address = _RAND_350[63:0];
  _RAND_351 = {1{`RANDOM}};
  btb_87_bht = _RAND_351[1:0];
  _RAND_352 = {1{`RANDOM}};
  btb_88_valid = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  btb_88_tag = _RAND_353[9:0];
  _RAND_354 = {2{`RANDOM}};
  btb_88_target_address = _RAND_354[63:0];
  _RAND_355 = {1{`RANDOM}};
  btb_88_bht = _RAND_355[1:0];
  _RAND_356 = {1{`RANDOM}};
  btb_89_valid = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  btb_89_tag = _RAND_357[9:0];
  _RAND_358 = {2{`RANDOM}};
  btb_89_target_address = _RAND_358[63:0];
  _RAND_359 = {1{`RANDOM}};
  btb_89_bht = _RAND_359[1:0];
  _RAND_360 = {1{`RANDOM}};
  btb_90_valid = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  btb_90_tag = _RAND_361[9:0];
  _RAND_362 = {2{`RANDOM}};
  btb_90_target_address = _RAND_362[63:0];
  _RAND_363 = {1{`RANDOM}};
  btb_90_bht = _RAND_363[1:0];
  _RAND_364 = {1{`RANDOM}};
  btb_91_valid = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  btb_91_tag = _RAND_365[9:0];
  _RAND_366 = {2{`RANDOM}};
  btb_91_target_address = _RAND_366[63:0];
  _RAND_367 = {1{`RANDOM}};
  btb_91_bht = _RAND_367[1:0];
  _RAND_368 = {1{`RANDOM}};
  btb_92_valid = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  btb_92_tag = _RAND_369[9:0];
  _RAND_370 = {2{`RANDOM}};
  btb_92_target_address = _RAND_370[63:0];
  _RAND_371 = {1{`RANDOM}};
  btb_92_bht = _RAND_371[1:0];
  _RAND_372 = {1{`RANDOM}};
  btb_93_valid = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  btb_93_tag = _RAND_373[9:0];
  _RAND_374 = {2{`RANDOM}};
  btb_93_target_address = _RAND_374[63:0];
  _RAND_375 = {1{`RANDOM}};
  btb_93_bht = _RAND_375[1:0];
  _RAND_376 = {1{`RANDOM}};
  btb_94_valid = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  btb_94_tag = _RAND_377[9:0];
  _RAND_378 = {2{`RANDOM}};
  btb_94_target_address = _RAND_378[63:0];
  _RAND_379 = {1{`RANDOM}};
  btb_94_bht = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  btb_95_valid = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  btb_95_tag = _RAND_381[9:0];
  _RAND_382 = {2{`RANDOM}};
  btb_95_target_address = _RAND_382[63:0];
  _RAND_383 = {1{`RANDOM}};
  btb_95_bht = _RAND_383[1:0];
  _RAND_384 = {1{`RANDOM}};
  btb_96_valid = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  btb_96_tag = _RAND_385[9:0];
  _RAND_386 = {2{`RANDOM}};
  btb_96_target_address = _RAND_386[63:0];
  _RAND_387 = {1{`RANDOM}};
  btb_96_bht = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  btb_97_valid = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  btb_97_tag = _RAND_389[9:0];
  _RAND_390 = {2{`RANDOM}};
  btb_97_target_address = _RAND_390[63:0];
  _RAND_391 = {1{`RANDOM}};
  btb_97_bht = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  btb_98_valid = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  btb_98_tag = _RAND_393[9:0];
  _RAND_394 = {2{`RANDOM}};
  btb_98_target_address = _RAND_394[63:0];
  _RAND_395 = {1{`RANDOM}};
  btb_98_bht = _RAND_395[1:0];
  _RAND_396 = {1{`RANDOM}};
  btb_99_valid = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  btb_99_tag = _RAND_397[9:0];
  _RAND_398 = {2{`RANDOM}};
  btb_99_target_address = _RAND_398[63:0];
  _RAND_399 = {1{`RANDOM}};
  btb_99_bht = _RAND_399[1:0];
  _RAND_400 = {1{`RANDOM}};
  btb_100_valid = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  btb_100_tag = _RAND_401[9:0];
  _RAND_402 = {2{`RANDOM}};
  btb_100_target_address = _RAND_402[63:0];
  _RAND_403 = {1{`RANDOM}};
  btb_100_bht = _RAND_403[1:0];
  _RAND_404 = {1{`RANDOM}};
  btb_101_valid = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  btb_101_tag = _RAND_405[9:0];
  _RAND_406 = {2{`RANDOM}};
  btb_101_target_address = _RAND_406[63:0];
  _RAND_407 = {1{`RANDOM}};
  btb_101_bht = _RAND_407[1:0];
  _RAND_408 = {1{`RANDOM}};
  btb_102_valid = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  btb_102_tag = _RAND_409[9:0];
  _RAND_410 = {2{`RANDOM}};
  btb_102_target_address = _RAND_410[63:0];
  _RAND_411 = {1{`RANDOM}};
  btb_102_bht = _RAND_411[1:0];
  _RAND_412 = {1{`RANDOM}};
  btb_103_valid = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  btb_103_tag = _RAND_413[9:0];
  _RAND_414 = {2{`RANDOM}};
  btb_103_target_address = _RAND_414[63:0];
  _RAND_415 = {1{`RANDOM}};
  btb_103_bht = _RAND_415[1:0];
  _RAND_416 = {1{`RANDOM}};
  btb_104_valid = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  btb_104_tag = _RAND_417[9:0];
  _RAND_418 = {2{`RANDOM}};
  btb_104_target_address = _RAND_418[63:0];
  _RAND_419 = {1{`RANDOM}};
  btb_104_bht = _RAND_419[1:0];
  _RAND_420 = {1{`RANDOM}};
  btb_105_valid = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  btb_105_tag = _RAND_421[9:0];
  _RAND_422 = {2{`RANDOM}};
  btb_105_target_address = _RAND_422[63:0];
  _RAND_423 = {1{`RANDOM}};
  btb_105_bht = _RAND_423[1:0];
  _RAND_424 = {1{`RANDOM}};
  btb_106_valid = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  btb_106_tag = _RAND_425[9:0];
  _RAND_426 = {2{`RANDOM}};
  btb_106_target_address = _RAND_426[63:0];
  _RAND_427 = {1{`RANDOM}};
  btb_106_bht = _RAND_427[1:0];
  _RAND_428 = {1{`RANDOM}};
  btb_107_valid = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  btb_107_tag = _RAND_429[9:0];
  _RAND_430 = {2{`RANDOM}};
  btb_107_target_address = _RAND_430[63:0];
  _RAND_431 = {1{`RANDOM}};
  btb_107_bht = _RAND_431[1:0];
  _RAND_432 = {1{`RANDOM}};
  btb_108_valid = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  btb_108_tag = _RAND_433[9:0];
  _RAND_434 = {2{`RANDOM}};
  btb_108_target_address = _RAND_434[63:0];
  _RAND_435 = {1{`RANDOM}};
  btb_108_bht = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  btb_109_valid = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  btb_109_tag = _RAND_437[9:0];
  _RAND_438 = {2{`RANDOM}};
  btb_109_target_address = _RAND_438[63:0];
  _RAND_439 = {1{`RANDOM}};
  btb_109_bht = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  btb_110_valid = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  btb_110_tag = _RAND_441[9:0];
  _RAND_442 = {2{`RANDOM}};
  btb_110_target_address = _RAND_442[63:0];
  _RAND_443 = {1{`RANDOM}};
  btb_110_bht = _RAND_443[1:0];
  _RAND_444 = {1{`RANDOM}};
  btb_111_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  btb_111_tag = _RAND_445[9:0];
  _RAND_446 = {2{`RANDOM}};
  btb_111_target_address = _RAND_446[63:0];
  _RAND_447 = {1{`RANDOM}};
  btb_111_bht = _RAND_447[1:0];
  _RAND_448 = {1{`RANDOM}};
  btb_112_valid = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  btb_112_tag = _RAND_449[9:0];
  _RAND_450 = {2{`RANDOM}};
  btb_112_target_address = _RAND_450[63:0];
  _RAND_451 = {1{`RANDOM}};
  btb_112_bht = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  btb_113_valid = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  btb_113_tag = _RAND_453[9:0];
  _RAND_454 = {2{`RANDOM}};
  btb_113_target_address = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  btb_113_bht = _RAND_455[1:0];
  _RAND_456 = {1{`RANDOM}};
  btb_114_valid = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  btb_114_tag = _RAND_457[9:0];
  _RAND_458 = {2{`RANDOM}};
  btb_114_target_address = _RAND_458[63:0];
  _RAND_459 = {1{`RANDOM}};
  btb_114_bht = _RAND_459[1:0];
  _RAND_460 = {1{`RANDOM}};
  btb_115_valid = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  btb_115_tag = _RAND_461[9:0];
  _RAND_462 = {2{`RANDOM}};
  btb_115_target_address = _RAND_462[63:0];
  _RAND_463 = {1{`RANDOM}};
  btb_115_bht = _RAND_463[1:0];
  _RAND_464 = {1{`RANDOM}};
  btb_116_valid = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  btb_116_tag = _RAND_465[9:0];
  _RAND_466 = {2{`RANDOM}};
  btb_116_target_address = _RAND_466[63:0];
  _RAND_467 = {1{`RANDOM}};
  btb_116_bht = _RAND_467[1:0];
  _RAND_468 = {1{`RANDOM}};
  btb_117_valid = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  btb_117_tag = _RAND_469[9:0];
  _RAND_470 = {2{`RANDOM}};
  btb_117_target_address = _RAND_470[63:0];
  _RAND_471 = {1{`RANDOM}};
  btb_117_bht = _RAND_471[1:0];
  _RAND_472 = {1{`RANDOM}};
  btb_118_valid = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  btb_118_tag = _RAND_473[9:0];
  _RAND_474 = {2{`RANDOM}};
  btb_118_target_address = _RAND_474[63:0];
  _RAND_475 = {1{`RANDOM}};
  btb_118_bht = _RAND_475[1:0];
  _RAND_476 = {1{`RANDOM}};
  btb_119_valid = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  btb_119_tag = _RAND_477[9:0];
  _RAND_478 = {2{`RANDOM}};
  btb_119_target_address = _RAND_478[63:0];
  _RAND_479 = {1{`RANDOM}};
  btb_119_bht = _RAND_479[1:0];
  _RAND_480 = {1{`RANDOM}};
  btb_120_valid = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  btb_120_tag = _RAND_481[9:0];
  _RAND_482 = {2{`RANDOM}};
  btb_120_target_address = _RAND_482[63:0];
  _RAND_483 = {1{`RANDOM}};
  btb_120_bht = _RAND_483[1:0];
  _RAND_484 = {1{`RANDOM}};
  btb_121_valid = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  btb_121_tag = _RAND_485[9:0];
  _RAND_486 = {2{`RANDOM}};
  btb_121_target_address = _RAND_486[63:0];
  _RAND_487 = {1{`RANDOM}};
  btb_121_bht = _RAND_487[1:0];
  _RAND_488 = {1{`RANDOM}};
  btb_122_valid = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  btb_122_tag = _RAND_489[9:0];
  _RAND_490 = {2{`RANDOM}};
  btb_122_target_address = _RAND_490[63:0];
  _RAND_491 = {1{`RANDOM}};
  btb_122_bht = _RAND_491[1:0];
  _RAND_492 = {1{`RANDOM}};
  btb_123_valid = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  btb_123_tag = _RAND_493[9:0];
  _RAND_494 = {2{`RANDOM}};
  btb_123_target_address = _RAND_494[63:0];
  _RAND_495 = {1{`RANDOM}};
  btb_123_bht = _RAND_495[1:0];
  _RAND_496 = {1{`RANDOM}};
  btb_124_valid = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  btb_124_tag = _RAND_497[9:0];
  _RAND_498 = {2{`RANDOM}};
  btb_124_target_address = _RAND_498[63:0];
  _RAND_499 = {1{`RANDOM}};
  btb_124_bht = _RAND_499[1:0];
  _RAND_500 = {1{`RANDOM}};
  btb_125_valid = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  btb_125_tag = _RAND_501[9:0];
  _RAND_502 = {2{`RANDOM}};
  btb_125_target_address = _RAND_502[63:0];
  _RAND_503 = {1{`RANDOM}};
  btb_125_bht = _RAND_503[1:0];
  _RAND_504 = {1{`RANDOM}};
  btb_126_valid = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  btb_126_tag = _RAND_505[9:0];
  _RAND_506 = {2{`RANDOM}};
  btb_126_target_address = _RAND_506[63:0];
  _RAND_507 = {1{`RANDOM}};
  btb_126_bht = _RAND_507[1:0];
  _RAND_508 = {1{`RANDOM}};
  btb_127_valid = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  btb_127_tag = _RAND_509[9:0];
  _RAND_510 = {2{`RANDOM}};
  btb_127_target_address = _RAND_510[63:0];
  _RAND_511 = {1{`RANDOM}};
  btb_127_bht = _RAND_511[1:0];
  _RAND_512 = {1{`RANDOM}};
  btb_128_valid = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  btb_128_tag = _RAND_513[9:0];
  _RAND_514 = {2{`RANDOM}};
  btb_128_target_address = _RAND_514[63:0];
  _RAND_515 = {1{`RANDOM}};
  btb_128_bht = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  btb_129_valid = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  btb_129_tag = _RAND_517[9:0];
  _RAND_518 = {2{`RANDOM}};
  btb_129_target_address = _RAND_518[63:0];
  _RAND_519 = {1{`RANDOM}};
  btb_129_bht = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  btb_130_valid = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  btb_130_tag = _RAND_521[9:0];
  _RAND_522 = {2{`RANDOM}};
  btb_130_target_address = _RAND_522[63:0];
  _RAND_523 = {1{`RANDOM}};
  btb_130_bht = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  btb_131_valid = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  btb_131_tag = _RAND_525[9:0];
  _RAND_526 = {2{`RANDOM}};
  btb_131_target_address = _RAND_526[63:0];
  _RAND_527 = {1{`RANDOM}};
  btb_131_bht = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  btb_132_valid = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  btb_132_tag = _RAND_529[9:0];
  _RAND_530 = {2{`RANDOM}};
  btb_132_target_address = _RAND_530[63:0];
  _RAND_531 = {1{`RANDOM}};
  btb_132_bht = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  btb_133_valid = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  btb_133_tag = _RAND_533[9:0];
  _RAND_534 = {2{`RANDOM}};
  btb_133_target_address = _RAND_534[63:0];
  _RAND_535 = {1{`RANDOM}};
  btb_133_bht = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  btb_134_valid = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  btb_134_tag = _RAND_537[9:0];
  _RAND_538 = {2{`RANDOM}};
  btb_134_target_address = _RAND_538[63:0];
  _RAND_539 = {1{`RANDOM}};
  btb_134_bht = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  btb_135_valid = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  btb_135_tag = _RAND_541[9:0];
  _RAND_542 = {2{`RANDOM}};
  btb_135_target_address = _RAND_542[63:0];
  _RAND_543 = {1{`RANDOM}};
  btb_135_bht = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  btb_136_valid = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  btb_136_tag = _RAND_545[9:0];
  _RAND_546 = {2{`RANDOM}};
  btb_136_target_address = _RAND_546[63:0];
  _RAND_547 = {1{`RANDOM}};
  btb_136_bht = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  btb_137_valid = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  btb_137_tag = _RAND_549[9:0];
  _RAND_550 = {2{`RANDOM}};
  btb_137_target_address = _RAND_550[63:0];
  _RAND_551 = {1{`RANDOM}};
  btb_137_bht = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  btb_138_valid = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  btb_138_tag = _RAND_553[9:0];
  _RAND_554 = {2{`RANDOM}};
  btb_138_target_address = _RAND_554[63:0];
  _RAND_555 = {1{`RANDOM}};
  btb_138_bht = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  btb_139_valid = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  btb_139_tag = _RAND_557[9:0];
  _RAND_558 = {2{`RANDOM}};
  btb_139_target_address = _RAND_558[63:0];
  _RAND_559 = {1{`RANDOM}};
  btb_139_bht = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  btb_140_valid = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  btb_140_tag = _RAND_561[9:0];
  _RAND_562 = {2{`RANDOM}};
  btb_140_target_address = _RAND_562[63:0];
  _RAND_563 = {1{`RANDOM}};
  btb_140_bht = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  btb_141_valid = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  btb_141_tag = _RAND_565[9:0];
  _RAND_566 = {2{`RANDOM}};
  btb_141_target_address = _RAND_566[63:0];
  _RAND_567 = {1{`RANDOM}};
  btb_141_bht = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  btb_142_valid = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  btb_142_tag = _RAND_569[9:0];
  _RAND_570 = {2{`RANDOM}};
  btb_142_target_address = _RAND_570[63:0];
  _RAND_571 = {1{`RANDOM}};
  btb_142_bht = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  btb_143_valid = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  btb_143_tag = _RAND_573[9:0];
  _RAND_574 = {2{`RANDOM}};
  btb_143_target_address = _RAND_574[63:0];
  _RAND_575 = {1{`RANDOM}};
  btb_143_bht = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  btb_144_valid = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  btb_144_tag = _RAND_577[9:0];
  _RAND_578 = {2{`RANDOM}};
  btb_144_target_address = _RAND_578[63:0];
  _RAND_579 = {1{`RANDOM}};
  btb_144_bht = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  btb_145_valid = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  btb_145_tag = _RAND_581[9:0];
  _RAND_582 = {2{`RANDOM}};
  btb_145_target_address = _RAND_582[63:0];
  _RAND_583 = {1{`RANDOM}};
  btb_145_bht = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  btb_146_valid = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  btb_146_tag = _RAND_585[9:0];
  _RAND_586 = {2{`RANDOM}};
  btb_146_target_address = _RAND_586[63:0];
  _RAND_587 = {1{`RANDOM}};
  btb_146_bht = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  btb_147_valid = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  btb_147_tag = _RAND_589[9:0];
  _RAND_590 = {2{`RANDOM}};
  btb_147_target_address = _RAND_590[63:0];
  _RAND_591 = {1{`RANDOM}};
  btb_147_bht = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  btb_148_valid = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  btb_148_tag = _RAND_593[9:0];
  _RAND_594 = {2{`RANDOM}};
  btb_148_target_address = _RAND_594[63:0];
  _RAND_595 = {1{`RANDOM}};
  btb_148_bht = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  btb_149_valid = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  btb_149_tag = _RAND_597[9:0];
  _RAND_598 = {2{`RANDOM}};
  btb_149_target_address = _RAND_598[63:0];
  _RAND_599 = {1{`RANDOM}};
  btb_149_bht = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  btb_150_valid = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  btb_150_tag = _RAND_601[9:0];
  _RAND_602 = {2{`RANDOM}};
  btb_150_target_address = _RAND_602[63:0];
  _RAND_603 = {1{`RANDOM}};
  btb_150_bht = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  btb_151_valid = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  btb_151_tag = _RAND_605[9:0];
  _RAND_606 = {2{`RANDOM}};
  btb_151_target_address = _RAND_606[63:0];
  _RAND_607 = {1{`RANDOM}};
  btb_151_bht = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  btb_152_valid = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  btb_152_tag = _RAND_609[9:0];
  _RAND_610 = {2{`RANDOM}};
  btb_152_target_address = _RAND_610[63:0];
  _RAND_611 = {1{`RANDOM}};
  btb_152_bht = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  btb_153_valid = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  btb_153_tag = _RAND_613[9:0];
  _RAND_614 = {2{`RANDOM}};
  btb_153_target_address = _RAND_614[63:0];
  _RAND_615 = {1{`RANDOM}};
  btb_153_bht = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  btb_154_valid = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  btb_154_tag = _RAND_617[9:0];
  _RAND_618 = {2{`RANDOM}};
  btb_154_target_address = _RAND_618[63:0];
  _RAND_619 = {1{`RANDOM}};
  btb_154_bht = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  btb_155_valid = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  btb_155_tag = _RAND_621[9:0];
  _RAND_622 = {2{`RANDOM}};
  btb_155_target_address = _RAND_622[63:0];
  _RAND_623 = {1{`RANDOM}};
  btb_155_bht = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  btb_156_valid = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  btb_156_tag = _RAND_625[9:0];
  _RAND_626 = {2{`RANDOM}};
  btb_156_target_address = _RAND_626[63:0];
  _RAND_627 = {1{`RANDOM}};
  btb_156_bht = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  btb_157_valid = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  btb_157_tag = _RAND_629[9:0];
  _RAND_630 = {2{`RANDOM}};
  btb_157_target_address = _RAND_630[63:0];
  _RAND_631 = {1{`RANDOM}};
  btb_157_bht = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  btb_158_valid = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  btb_158_tag = _RAND_633[9:0];
  _RAND_634 = {2{`RANDOM}};
  btb_158_target_address = _RAND_634[63:0];
  _RAND_635 = {1{`RANDOM}};
  btb_158_bht = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  btb_159_valid = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  btb_159_tag = _RAND_637[9:0];
  _RAND_638 = {2{`RANDOM}};
  btb_159_target_address = _RAND_638[63:0];
  _RAND_639 = {1{`RANDOM}};
  btb_159_bht = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  btb_160_valid = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  btb_160_tag = _RAND_641[9:0];
  _RAND_642 = {2{`RANDOM}};
  btb_160_target_address = _RAND_642[63:0];
  _RAND_643 = {1{`RANDOM}};
  btb_160_bht = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  btb_161_valid = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  btb_161_tag = _RAND_645[9:0];
  _RAND_646 = {2{`RANDOM}};
  btb_161_target_address = _RAND_646[63:0];
  _RAND_647 = {1{`RANDOM}};
  btb_161_bht = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  btb_162_valid = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  btb_162_tag = _RAND_649[9:0];
  _RAND_650 = {2{`RANDOM}};
  btb_162_target_address = _RAND_650[63:0];
  _RAND_651 = {1{`RANDOM}};
  btb_162_bht = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  btb_163_valid = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  btb_163_tag = _RAND_653[9:0];
  _RAND_654 = {2{`RANDOM}};
  btb_163_target_address = _RAND_654[63:0];
  _RAND_655 = {1{`RANDOM}};
  btb_163_bht = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  btb_164_valid = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  btb_164_tag = _RAND_657[9:0];
  _RAND_658 = {2{`RANDOM}};
  btb_164_target_address = _RAND_658[63:0];
  _RAND_659 = {1{`RANDOM}};
  btb_164_bht = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  btb_165_valid = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  btb_165_tag = _RAND_661[9:0];
  _RAND_662 = {2{`RANDOM}};
  btb_165_target_address = _RAND_662[63:0];
  _RAND_663 = {1{`RANDOM}};
  btb_165_bht = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  btb_166_valid = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  btb_166_tag = _RAND_665[9:0];
  _RAND_666 = {2{`RANDOM}};
  btb_166_target_address = _RAND_666[63:0];
  _RAND_667 = {1{`RANDOM}};
  btb_166_bht = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  btb_167_valid = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  btb_167_tag = _RAND_669[9:0];
  _RAND_670 = {2{`RANDOM}};
  btb_167_target_address = _RAND_670[63:0];
  _RAND_671 = {1{`RANDOM}};
  btb_167_bht = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  btb_168_valid = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  btb_168_tag = _RAND_673[9:0];
  _RAND_674 = {2{`RANDOM}};
  btb_168_target_address = _RAND_674[63:0];
  _RAND_675 = {1{`RANDOM}};
  btb_168_bht = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  btb_169_valid = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  btb_169_tag = _RAND_677[9:0];
  _RAND_678 = {2{`RANDOM}};
  btb_169_target_address = _RAND_678[63:0];
  _RAND_679 = {1{`RANDOM}};
  btb_169_bht = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  btb_170_valid = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  btb_170_tag = _RAND_681[9:0];
  _RAND_682 = {2{`RANDOM}};
  btb_170_target_address = _RAND_682[63:0];
  _RAND_683 = {1{`RANDOM}};
  btb_170_bht = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  btb_171_valid = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  btb_171_tag = _RAND_685[9:0];
  _RAND_686 = {2{`RANDOM}};
  btb_171_target_address = _RAND_686[63:0];
  _RAND_687 = {1{`RANDOM}};
  btb_171_bht = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  btb_172_valid = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  btb_172_tag = _RAND_689[9:0];
  _RAND_690 = {2{`RANDOM}};
  btb_172_target_address = _RAND_690[63:0];
  _RAND_691 = {1{`RANDOM}};
  btb_172_bht = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  btb_173_valid = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  btb_173_tag = _RAND_693[9:0];
  _RAND_694 = {2{`RANDOM}};
  btb_173_target_address = _RAND_694[63:0];
  _RAND_695 = {1{`RANDOM}};
  btb_173_bht = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  btb_174_valid = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  btb_174_tag = _RAND_697[9:0];
  _RAND_698 = {2{`RANDOM}};
  btb_174_target_address = _RAND_698[63:0];
  _RAND_699 = {1{`RANDOM}};
  btb_174_bht = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  btb_175_valid = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  btb_175_tag = _RAND_701[9:0];
  _RAND_702 = {2{`RANDOM}};
  btb_175_target_address = _RAND_702[63:0];
  _RAND_703 = {1{`RANDOM}};
  btb_175_bht = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  btb_176_valid = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  btb_176_tag = _RAND_705[9:0];
  _RAND_706 = {2{`RANDOM}};
  btb_176_target_address = _RAND_706[63:0];
  _RAND_707 = {1{`RANDOM}};
  btb_176_bht = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  btb_177_valid = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  btb_177_tag = _RAND_709[9:0];
  _RAND_710 = {2{`RANDOM}};
  btb_177_target_address = _RAND_710[63:0];
  _RAND_711 = {1{`RANDOM}};
  btb_177_bht = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  btb_178_valid = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  btb_178_tag = _RAND_713[9:0];
  _RAND_714 = {2{`RANDOM}};
  btb_178_target_address = _RAND_714[63:0];
  _RAND_715 = {1{`RANDOM}};
  btb_178_bht = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  btb_179_valid = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  btb_179_tag = _RAND_717[9:0];
  _RAND_718 = {2{`RANDOM}};
  btb_179_target_address = _RAND_718[63:0];
  _RAND_719 = {1{`RANDOM}};
  btb_179_bht = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  btb_180_valid = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  btb_180_tag = _RAND_721[9:0];
  _RAND_722 = {2{`RANDOM}};
  btb_180_target_address = _RAND_722[63:0];
  _RAND_723 = {1{`RANDOM}};
  btb_180_bht = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  btb_181_valid = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  btb_181_tag = _RAND_725[9:0];
  _RAND_726 = {2{`RANDOM}};
  btb_181_target_address = _RAND_726[63:0];
  _RAND_727 = {1{`RANDOM}};
  btb_181_bht = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  btb_182_valid = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  btb_182_tag = _RAND_729[9:0];
  _RAND_730 = {2{`RANDOM}};
  btb_182_target_address = _RAND_730[63:0];
  _RAND_731 = {1{`RANDOM}};
  btb_182_bht = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  btb_183_valid = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  btb_183_tag = _RAND_733[9:0];
  _RAND_734 = {2{`RANDOM}};
  btb_183_target_address = _RAND_734[63:0];
  _RAND_735 = {1{`RANDOM}};
  btb_183_bht = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  btb_184_valid = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  btb_184_tag = _RAND_737[9:0];
  _RAND_738 = {2{`RANDOM}};
  btb_184_target_address = _RAND_738[63:0];
  _RAND_739 = {1{`RANDOM}};
  btb_184_bht = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  btb_185_valid = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  btb_185_tag = _RAND_741[9:0];
  _RAND_742 = {2{`RANDOM}};
  btb_185_target_address = _RAND_742[63:0];
  _RAND_743 = {1{`RANDOM}};
  btb_185_bht = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  btb_186_valid = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  btb_186_tag = _RAND_745[9:0];
  _RAND_746 = {2{`RANDOM}};
  btb_186_target_address = _RAND_746[63:0];
  _RAND_747 = {1{`RANDOM}};
  btb_186_bht = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  btb_187_valid = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  btb_187_tag = _RAND_749[9:0];
  _RAND_750 = {2{`RANDOM}};
  btb_187_target_address = _RAND_750[63:0];
  _RAND_751 = {1{`RANDOM}};
  btb_187_bht = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  btb_188_valid = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  btb_188_tag = _RAND_753[9:0];
  _RAND_754 = {2{`RANDOM}};
  btb_188_target_address = _RAND_754[63:0];
  _RAND_755 = {1{`RANDOM}};
  btb_188_bht = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  btb_189_valid = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  btb_189_tag = _RAND_757[9:0];
  _RAND_758 = {2{`RANDOM}};
  btb_189_target_address = _RAND_758[63:0];
  _RAND_759 = {1{`RANDOM}};
  btb_189_bht = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  btb_190_valid = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  btb_190_tag = _RAND_761[9:0];
  _RAND_762 = {2{`RANDOM}};
  btb_190_target_address = _RAND_762[63:0];
  _RAND_763 = {1{`RANDOM}};
  btb_190_bht = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  btb_191_valid = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  btb_191_tag = _RAND_765[9:0];
  _RAND_766 = {2{`RANDOM}};
  btb_191_target_address = _RAND_766[63:0];
  _RAND_767 = {1{`RANDOM}};
  btb_191_bht = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  btb_192_valid = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  btb_192_tag = _RAND_769[9:0];
  _RAND_770 = {2{`RANDOM}};
  btb_192_target_address = _RAND_770[63:0];
  _RAND_771 = {1{`RANDOM}};
  btb_192_bht = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  btb_193_valid = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  btb_193_tag = _RAND_773[9:0];
  _RAND_774 = {2{`RANDOM}};
  btb_193_target_address = _RAND_774[63:0];
  _RAND_775 = {1{`RANDOM}};
  btb_193_bht = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  btb_194_valid = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  btb_194_tag = _RAND_777[9:0];
  _RAND_778 = {2{`RANDOM}};
  btb_194_target_address = _RAND_778[63:0];
  _RAND_779 = {1{`RANDOM}};
  btb_194_bht = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  btb_195_valid = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  btb_195_tag = _RAND_781[9:0];
  _RAND_782 = {2{`RANDOM}};
  btb_195_target_address = _RAND_782[63:0];
  _RAND_783 = {1{`RANDOM}};
  btb_195_bht = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  btb_196_valid = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  btb_196_tag = _RAND_785[9:0];
  _RAND_786 = {2{`RANDOM}};
  btb_196_target_address = _RAND_786[63:0];
  _RAND_787 = {1{`RANDOM}};
  btb_196_bht = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  btb_197_valid = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  btb_197_tag = _RAND_789[9:0];
  _RAND_790 = {2{`RANDOM}};
  btb_197_target_address = _RAND_790[63:0];
  _RAND_791 = {1{`RANDOM}};
  btb_197_bht = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  btb_198_valid = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  btb_198_tag = _RAND_793[9:0];
  _RAND_794 = {2{`RANDOM}};
  btb_198_target_address = _RAND_794[63:0];
  _RAND_795 = {1{`RANDOM}};
  btb_198_bht = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  btb_199_valid = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  btb_199_tag = _RAND_797[9:0];
  _RAND_798 = {2{`RANDOM}};
  btb_199_target_address = _RAND_798[63:0];
  _RAND_799 = {1{`RANDOM}};
  btb_199_bht = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  btb_200_valid = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  btb_200_tag = _RAND_801[9:0];
  _RAND_802 = {2{`RANDOM}};
  btb_200_target_address = _RAND_802[63:0];
  _RAND_803 = {1{`RANDOM}};
  btb_200_bht = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  btb_201_valid = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  btb_201_tag = _RAND_805[9:0];
  _RAND_806 = {2{`RANDOM}};
  btb_201_target_address = _RAND_806[63:0];
  _RAND_807 = {1{`RANDOM}};
  btb_201_bht = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  btb_202_valid = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  btb_202_tag = _RAND_809[9:0];
  _RAND_810 = {2{`RANDOM}};
  btb_202_target_address = _RAND_810[63:0];
  _RAND_811 = {1{`RANDOM}};
  btb_202_bht = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  btb_203_valid = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  btb_203_tag = _RAND_813[9:0];
  _RAND_814 = {2{`RANDOM}};
  btb_203_target_address = _RAND_814[63:0];
  _RAND_815 = {1{`RANDOM}};
  btb_203_bht = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  btb_204_valid = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  btb_204_tag = _RAND_817[9:0];
  _RAND_818 = {2{`RANDOM}};
  btb_204_target_address = _RAND_818[63:0];
  _RAND_819 = {1{`RANDOM}};
  btb_204_bht = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  btb_205_valid = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  btb_205_tag = _RAND_821[9:0];
  _RAND_822 = {2{`RANDOM}};
  btb_205_target_address = _RAND_822[63:0];
  _RAND_823 = {1{`RANDOM}};
  btb_205_bht = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  btb_206_valid = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  btb_206_tag = _RAND_825[9:0];
  _RAND_826 = {2{`RANDOM}};
  btb_206_target_address = _RAND_826[63:0];
  _RAND_827 = {1{`RANDOM}};
  btb_206_bht = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  btb_207_valid = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  btb_207_tag = _RAND_829[9:0];
  _RAND_830 = {2{`RANDOM}};
  btb_207_target_address = _RAND_830[63:0];
  _RAND_831 = {1{`RANDOM}};
  btb_207_bht = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  btb_208_valid = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  btb_208_tag = _RAND_833[9:0];
  _RAND_834 = {2{`RANDOM}};
  btb_208_target_address = _RAND_834[63:0];
  _RAND_835 = {1{`RANDOM}};
  btb_208_bht = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  btb_209_valid = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  btb_209_tag = _RAND_837[9:0];
  _RAND_838 = {2{`RANDOM}};
  btb_209_target_address = _RAND_838[63:0];
  _RAND_839 = {1{`RANDOM}};
  btb_209_bht = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  btb_210_valid = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  btb_210_tag = _RAND_841[9:0];
  _RAND_842 = {2{`RANDOM}};
  btb_210_target_address = _RAND_842[63:0];
  _RAND_843 = {1{`RANDOM}};
  btb_210_bht = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  btb_211_valid = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  btb_211_tag = _RAND_845[9:0];
  _RAND_846 = {2{`RANDOM}};
  btb_211_target_address = _RAND_846[63:0];
  _RAND_847 = {1{`RANDOM}};
  btb_211_bht = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  btb_212_valid = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  btb_212_tag = _RAND_849[9:0];
  _RAND_850 = {2{`RANDOM}};
  btb_212_target_address = _RAND_850[63:0];
  _RAND_851 = {1{`RANDOM}};
  btb_212_bht = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  btb_213_valid = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  btb_213_tag = _RAND_853[9:0];
  _RAND_854 = {2{`RANDOM}};
  btb_213_target_address = _RAND_854[63:0];
  _RAND_855 = {1{`RANDOM}};
  btb_213_bht = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  btb_214_valid = _RAND_856[0:0];
  _RAND_857 = {1{`RANDOM}};
  btb_214_tag = _RAND_857[9:0];
  _RAND_858 = {2{`RANDOM}};
  btb_214_target_address = _RAND_858[63:0];
  _RAND_859 = {1{`RANDOM}};
  btb_214_bht = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  btb_215_valid = _RAND_860[0:0];
  _RAND_861 = {1{`RANDOM}};
  btb_215_tag = _RAND_861[9:0];
  _RAND_862 = {2{`RANDOM}};
  btb_215_target_address = _RAND_862[63:0];
  _RAND_863 = {1{`RANDOM}};
  btb_215_bht = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  btb_216_valid = _RAND_864[0:0];
  _RAND_865 = {1{`RANDOM}};
  btb_216_tag = _RAND_865[9:0];
  _RAND_866 = {2{`RANDOM}};
  btb_216_target_address = _RAND_866[63:0];
  _RAND_867 = {1{`RANDOM}};
  btb_216_bht = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  btb_217_valid = _RAND_868[0:0];
  _RAND_869 = {1{`RANDOM}};
  btb_217_tag = _RAND_869[9:0];
  _RAND_870 = {2{`RANDOM}};
  btb_217_target_address = _RAND_870[63:0];
  _RAND_871 = {1{`RANDOM}};
  btb_217_bht = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  btb_218_valid = _RAND_872[0:0];
  _RAND_873 = {1{`RANDOM}};
  btb_218_tag = _RAND_873[9:0];
  _RAND_874 = {2{`RANDOM}};
  btb_218_target_address = _RAND_874[63:0];
  _RAND_875 = {1{`RANDOM}};
  btb_218_bht = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  btb_219_valid = _RAND_876[0:0];
  _RAND_877 = {1{`RANDOM}};
  btb_219_tag = _RAND_877[9:0];
  _RAND_878 = {2{`RANDOM}};
  btb_219_target_address = _RAND_878[63:0];
  _RAND_879 = {1{`RANDOM}};
  btb_219_bht = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  btb_220_valid = _RAND_880[0:0];
  _RAND_881 = {1{`RANDOM}};
  btb_220_tag = _RAND_881[9:0];
  _RAND_882 = {2{`RANDOM}};
  btb_220_target_address = _RAND_882[63:0];
  _RAND_883 = {1{`RANDOM}};
  btb_220_bht = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  btb_221_valid = _RAND_884[0:0];
  _RAND_885 = {1{`RANDOM}};
  btb_221_tag = _RAND_885[9:0];
  _RAND_886 = {2{`RANDOM}};
  btb_221_target_address = _RAND_886[63:0];
  _RAND_887 = {1{`RANDOM}};
  btb_221_bht = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  btb_222_valid = _RAND_888[0:0];
  _RAND_889 = {1{`RANDOM}};
  btb_222_tag = _RAND_889[9:0];
  _RAND_890 = {2{`RANDOM}};
  btb_222_target_address = _RAND_890[63:0];
  _RAND_891 = {1{`RANDOM}};
  btb_222_bht = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  btb_223_valid = _RAND_892[0:0];
  _RAND_893 = {1{`RANDOM}};
  btb_223_tag = _RAND_893[9:0];
  _RAND_894 = {2{`RANDOM}};
  btb_223_target_address = _RAND_894[63:0];
  _RAND_895 = {1{`RANDOM}};
  btb_223_bht = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  btb_224_valid = _RAND_896[0:0];
  _RAND_897 = {1{`RANDOM}};
  btb_224_tag = _RAND_897[9:0];
  _RAND_898 = {2{`RANDOM}};
  btb_224_target_address = _RAND_898[63:0];
  _RAND_899 = {1{`RANDOM}};
  btb_224_bht = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  btb_225_valid = _RAND_900[0:0];
  _RAND_901 = {1{`RANDOM}};
  btb_225_tag = _RAND_901[9:0];
  _RAND_902 = {2{`RANDOM}};
  btb_225_target_address = _RAND_902[63:0];
  _RAND_903 = {1{`RANDOM}};
  btb_225_bht = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  btb_226_valid = _RAND_904[0:0];
  _RAND_905 = {1{`RANDOM}};
  btb_226_tag = _RAND_905[9:0];
  _RAND_906 = {2{`RANDOM}};
  btb_226_target_address = _RAND_906[63:0];
  _RAND_907 = {1{`RANDOM}};
  btb_226_bht = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  btb_227_valid = _RAND_908[0:0];
  _RAND_909 = {1{`RANDOM}};
  btb_227_tag = _RAND_909[9:0];
  _RAND_910 = {2{`RANDOM}};
  btb_227_target_address = _RAND_910[63:0];
  _RAND_911 = {1{`RANDOM}};
  btb_227_bht = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  btb_228_valid = _RAND_912[0:0];
  _RAND_913 = {1{`RANDOM}};
  btb_228_tag = _RAND_913[9:0];
  _RAND_914 = {2{`RANDOM}};
  btb_228_target_address = _RAND_914[63:0];
  _RAND_915 = {1{`RANDOM}};
  btb_228_bht = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  btb_229_valid = _RAND_916[0:0];
  _RAND_917 = {1{`RANDOM}};
  btb_229_tag = _RAND_917[9:0];
  _RAND_918 = {2{`RANDOM}};
  btb_229_target_address = _RAND_918[63:0];
  _RAND_919 = {1{`RANDOM}};
  btb_229_bht = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  btb_230_valid = _RAND_920[0:0];
  _RAND_921 = {1{`RANDOM}};
  btb_230_tag = _RAND_921[9:0];
  _RAND_922 = {2{`RANDOM}};
  btb_230_target_address = _RAND_922[63:0];
  _RAND_923 = {1{`RANDOM}};
  btb_230_bht = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  btb_231_valid = _RAND_924[0:0];
  _RAND_925 = {1{`RANDOM}};
  btb_231_tag = _RAND_925[9:0];
  _RAND_926 = {2{`RANDOM}};
  btb_231_target_address = _RAND_926[63:0];
  _RAND_927 = {1{`RANDOM}};
  btb_231_bht = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  btb_232_valid = _RAND_928[0:0];
  _RAND_929 = {1{`RANDOM}};
  btb_232_tag = _RAND_929[9:0];
  _RAND_930 = {2{`RANDOM}};
  btb_232_target_address = _RAND_930[63:0];
  _RAND_931 = {1{`RANDOM}};
  btb_232_bht = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  btb_233_valid = _RAND_932[0:0];
  _RAND_933 = {1{`RANDOM}};
  btb_233_tag = _RAND_933[9:0];
  _RAND_934 = {2{`RANDOM}};
  btb_233_target_address = _RAND_934[63:0];
  _RAND_935 = {1{`RANDOM}};
  btb_233_bht = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  btb_234_valid = _RAND_936[0:0];
  _RAND_937 = {1{`RANDOM}};
  btb_234_tag = _RAND_937[9:0];
  _RAND_938 = {2{`RANDOM}};
  btb_234_target_address = _RAND_938[63:0];
  _RAND_939 = {1{`RANDOM}};
  btb_234_bht = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  btb_235_valid = _RAND_940[0:0];
  _RAND_941 = {1{`RANDOM}};
  btb_235_tag = _RAND_941[9:0];
  _RAND_942 = {2{`RANDOM}};
  btb_235_target_address = _RAND_942[63:0];
  _RAND_943 = {1{`RANDOM}};
  btb_235_bht = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  btb_236_valid = _RAND_944[0:0];
  _RAND_945 = {1{`RANDOM}};
  btb_236_tag = _RAND_945[9:0];
  _RAND_946 = {2{`RANDOM}};
  btb_236_target_address = _RAND_946[63:0];
  _RAND_947 = {1{`RANDOM}};
  btb_236_bht = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  btb_237_valid = _RAND_948[0:0];
  _RAND_949 = {1{`RANDOM}};
  btb_237_tag = _RAND_949[9:0];
  _RAND_950 = {2{`RANDOM}};
  btb_237_target_address = _RAND_950[63:0];
  _RAND_951 = {1{`RANDOM}};
  btb_237_bht = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  btb_238_valid = _RAND_952[0:0];
  _RAND_953 = {1{`RANDOM}};
  btb_238_tag = _RAND_953[9:0];
  _RAND_954 = {2{`RANDOM}};
  btb_238_target_address = _RAND_954[63:0];
  _RAND_955 = {1{`RANDOM}};
  btb_238_bht = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  btb_239_valid = _RAND_956[0:0];
  _RAND_957 = {1{`RANDOM}};
  btb_239_tag = _RAND_957[9:0];
  _RAND_958 = {2{`RANDOM}};
  btb_239_target_address = _RAND_958[63:0];
  _RAND_959 = {1{`RANDOM}};
  btb_239_bht = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  btb_240_valid = _RAND_960[0:0];
  _RAND_961 = {1{`RANDOM}};
  btb_240_tag = _RAND_961[9:0];
  _RAND_962 = {2{`RANDOM}};
  btb_240_target_address = _RAND_962[63:0];
  _RAND_963 = {1{`RANDOM}};
  btb_240_bht = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  btb_241_valid = _RAND_964[0:0];
  _RAND_965 = {1{`RANDOM}};
  btb_241_tag = _RAND_965[9:0];
  _RAND_966 = {2{`RANDOM}};
  btb_241_target_address = _RAND_966[63:0];
  _RAND_967 = {1{`RANDOM}};
  btb_241_bht = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  btb_242_valid = _RAND_968[0:0];
  _RAND_969 = {1{`RANDOM}};
  btb_242_tag = _RAND_969[9:0];
  _RAND_970 = {2{`RANDOM}};
  btb_242_target_address = _RAND_970[63:0];
  _RAND_971 = {1{`RANDOM}};
  btb_242_bht = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  btb_243_valid = _RAND_972[0:0];
  _RAND_973 = {1{`RANDOM}};
  btb_243_tag = _RAND_973[9:0];
  _RAND_974 = {2{`RANDOM}};
  btb_243_target_address = _RAND_974[63:0];
  _RAND_975 = {1{`RANDOM}};
  btb_243_bht = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  btb_244_valid = _RAND_976[0:0];
  _RAND_977 = {1{`RANDOM}};
  btb_244_tag = _RAND_977[9:0];
  _RAND_978 = {2{`RANDOM}};
  btb_244_target_address = _RAND_978[63:0];
  _RAND_979 = {1{`RANDOM}};
  btb_244_bht = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  btb_245_valid = _RAND_980[0:0];
  _RAND_981 = {1{`RANDOM}};
  btb_245_tag = _RAND_981[9:0];
  _RAND_982 = {2{`RANDOM}};
  btb_245_target_address = _RAND_982[63:0];
  _RAND_983 = {1{`RANDOM}};
  btb_245_bht = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  btb_246_valid = _RAND_984[0:0];
  _RAND_985 = {1{`RANDOM}};
  btb_246_tag = _RAND_985[9:0];
  _RAND_986 = {2{`RANDOM}};
  btb_246_target_address = _RAND_986[63:0];
  _RAND_987 = {1{`RANDOM}};
  btb_246_bht = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  btb_247_valid = _RAND_988[0:0];
  _RAND_989 = {1{`RANDOM}};
  btb_247_tag = _RAND_989[9:0];
  _RAND_990 = {2{`RANDOM}};
  btb_247_target_address = _RAND_990[63:0];
  _RAND_991 = {1{`RANDOM}};
  btb_247_bht = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  btb_248_valid = _RAND_992[0:0];
  _RAND_993 = {1{`RANDOM}};
  btb_248_tag = _RAND_993[9:0];
  _RAND_994 = {2{`RANDOM}};
  btb_248_target_address = _RAND_994[63:0];
  _RAND_995 = {1{`RANDOM}};
  btb_248_bht = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  btb_249_valid = _RAND_996[0:0];
  _RAND_997 = {1{`RANDOM}};
  btb_249_tag = _RAND_997[9:0];
  _RAND_998 = {2{`RANDOM}};
  btb_249_target_address = _RAND_998[63:0];
  _RAND_999 = {1{`RANDOM}};
  btb_249_bht = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  btb_250_valid = _RAND_1000[0:0];
  _RAND_1001 = {1{`RANDOM}};
  btb_250_tag = _RAND_1001[9:0];
  _RAND_1002 = {2{`RANDOM}};
  btb_250_target_address = _RAND_1002[63:0];
  _RAND_1003 = {1{`RANDOM}};
  btb_250_bht = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  btb_251_valid = _RAND_1004[0:0];
  _RAND_1005 = {1{`RANDOM}};
  btb_251_tag = _RAND_1005[9:0];
  _RAND_1006 = {2{`RANDOM}};
  btb_251_target_address = _RAND_1006[63:0];
  _RAND_1007 = {1{`RANDOM}};
  btb_251_bht = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  btb_252_valid = _RAND_1008[0:0];
  _RAND_1009 = {1{`RANDOM}};
  btb_252_tag = _RAND_1009[9:0];
  _RAND_1010 = {2{`RANDOM}};
  btb_252_target_address = _RAND_1010[63:0];
  _RAND_1011 = {1{`RANDOM}};
  btb_252_bht = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  btb_253_valid = _RAND_1012[0:0];
  _RAND_1013 = {1{`RANDOM}};
  btb_253_tag = _RAND_1013[9:0];
  _RAND_1014 = {2{`RANDOM}};
  btb_253_target_address = _RAND_1014[63:0];
  _RAND_1015 = {1{`RANDOM}};
  btb_253_bht = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  btb_254_valid = _RAND_1016[0:0];
  _RAND_1017 = {1{`RANDOM}};
  btb_254_tag = _RAND_1017[9:0];
  _RAND_1018 = {2{`RANDOM}};
  btb_254_target_address = _RAND_1018[63:0];
  _RAND_1019 = {1{`RANDOM}};
  btb_254_bht = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  btb_255_valid = _RAND_1020[0:0];
  _RAND_1021 = {1{`RANDOM}};
  btb_255_tag = _RAND_1021[9:0];
  _RAND_1022 = {2{`RANDOM}};
  btb_255_target_address = _RAND_1022[63:0];
  _RAND_1023 = {1{`RANDOM}};
  btb_255_bht = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  btb_256_valid = _RAND_1024[0:0];
  _RAND_1025 = {1{`RANDOM}};
  btb_256_tag = _RAND_1025[9:0];
  _RAND_1026 = {2{`RANDOM}};
  btb_256_target_address = _RAND_1026[63:0];
  _RAND_1027 = {1{`RANDOM}};
  btb_256_bht = _RAND_1027[1:0];
  _RAND_1028 = {1{`RANDOM}};
  btb_257_valid = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  btb_257_tag = _RAND_1029[9:0];
  _RAND_1030 = {2{`RANDOM}};
  btb_257_target_address = _RAND_1030[63:0];
  _RAND_1031 = {1{`RANDOM}};
  btb_257_bht = _RAND_1031[1:0];
  _RAND_1032 = {1{`RANDOM}};
  btb_258_valid = _RAND_1032[0:0];
  _RAND_1033 = {1{`RANDOM}};
  btb_258_tag = _RAND_1033[9:0];
  _RAND_1034 = {2{`RANDOM}};
  btb_258_target_address = _RAND_1034[63:0];
  _RAND_1035 = {1{`RANDOM}};
  btb_258_bht = _RAND_1035[1:0];
  _RAND_1036 = {1{`RANDOM}};
  btb_259_valid = _RAND_1036[0:0];
  _RAND_1037 = {1{`RANDOM}};
  btb_259_tag = _RAND_1037[9:0];
  _RAND_1038 = {2{`RANDOM}};
  btb_259_target_address = _RAND_1038[63:0];
  _RAND_1039 = {1{`RANDOM}};
  btb_259_bht = _RAND_1039[1:0];
  _RAND_1040 = {1{`RANDOM}};
  btb_260_valid = _RAND_1040[0:0];
  _RAND_1041 = {1{`RANDOM}};
  btb_260_tag = _RAND_1041[9:0];
  _RAND_1042 = {2{`RANDOM}};
  btb_260_target_address = _RAND_1042[63:0];
  _RAND_1043 = {1{`RANDOM}};
  btb_260_bht = _RAND_1043[1:0];
  _RAND_1044 = {1{`RANDOM}};
  btb_261_valid = _RAND_1044[0:0];
  _RAND_1045 = {1{`RANDOM}};
  btb_261_tag = _RAND_1045[9:0];
  _RAND_1046 = {2{`RANDOM}};
  btb_261_target_address = _RAND_1046[63:0];
  _RAND_1047 = {1{`RANDOM}};
  btb_261_bht = _RAND_1047[1:0];
  _RAND_1048 = {1{`RANDOM}};
  btb_262_valid = _RAND_1048[0:0];
  _RAND_1049 = {1{`RANDOM}};
  btb_262_tag = _RAND_1049[9:0];
  _RAND_1050 = {2{`RANDOM}};
  btb_262_target_address = _RAND_1050[63:0];
  _RAND_1051 = {1{`RANDOM}};
  btb_262_bht = _RAND_1051[1:0];
  _RAND_1052 = {1{`RANDOM}};
  btb_263_valid = _RAND_1052[0:0];
  _RAND_1053 = {1{`RANDOM}};
  btb_263_tag = _RAND_1053[9:0];
  _RAND_1054 = {2{`RANDOM}};
  btb_263_target_address = _RAND_1054[63:0];
  _RAND_1055 = {1{`RANDOM}};
  btb_263_bht = _RAND_1055[1:0];
  _RAND_1056 = {1{`RANDOM}};
  btb_264_valid = _RAND_1056[0:0];
  _RAND_1057 = {1{`RANDOM}};
  btb_264_tag = _RAND_1057[9:0];
  _RAND_1058 = {2{`RANDOM}};
  btb_264_target_address = _RAND_1058[63:0];
  _RAND_1059 = {1{`RANDOM}};
  btb_264_bht = _RAND_1059[1:0];
  _RAND_1060 = {1{`RANDOM}};
  btb_265_valid = _RAND_1060[0:0];
  _RAND_1061 = {1{`RANDOM}};
  btb_265_tag = _RAND_1061[9:0];
  _RAND_1062 = {2{`RANDOM}};
  btb_265_target_address = _RAND_1062[63:0];
  _RAND_1063 = {1{`RANDOM}};
  btb_265_bht = _RAND_1063[1:0];
  _RAND_1064 = {1{`RANDOM}};
  btb_266_valid = _RAND_1064[0:0];
  _RAND_1065 = {1{`RANDOM}};
  btb_266_tag = _RAND_1065[9:0];
  _RAND_1066 = {2{`RANDOM}};
  btb_266_target_address = _RAND_1066[63:0];
  _RAND_1067 = {1{`RANDOM}};
  btb_266_bht = _RAND_1067[1:0];
  _RAND_1068 = {1{`RANDOM}};
  btb_267_valid = _RAND_1068[0:0];
  _RAND_1069 = {1{`RANDOM}};
  btb_267_tag = _RAND_1069[9:0];
  _RAND_1070 = {2{`RANDOM}};
  btb_267_target_address = _RAND_1070[63:0];
  _RAND_1071 = {1{`RANDOM}};
  btb_267_bht = _RAND_1071[1:0];
  _RAND_1072 = {1{`RANDOM}};
  btb_268_valid = _RAND_1072[0:0];
  _RAND_1073 = {1{`RANDOM}};
  btb_268_tag = _RAND_1073[9:0];
  _RAND_1074 = {2{`RANDOM}};
  btb_268_target_address = _RAND_1074[63:0];
  _RAND_1075 = {1{`RANDOM}};
  btb_268_bht = _RAND_1075[1:0];
  _RAND_1076 = {1{`RANDOM}};
  btb_269_valid = _RAND_1076[0:0];
  _RAND_1077 = {1{`RANDOM}};
  btb_269_tag = _RAND_1077[9:0];
  _RAND_1078 = {2{`RANDOM}};
  btb_269_target_address = _RAND_1078[63:0];
  _RAND_1079 = {1{`RANDOM}};
  btb_269_bht = _RAND_1079[1:0];
  _RAND_1080 = {1{`RANDOM}};
  btb_270_valid = _RAND_1080[0:0];
  _RAND_1081 = {1{`RANDOM}};
  btb_270_tag = _RAND_1081[9:0];
  _RAND_1082 = {2{`RANDOM}};
  btb_270_target_address = _RAND_1082[63:0];
  _RAND_1083 = {1{`RANDOM}};
  btb_270_bht = _RAND_1083[1:0];
  _RAND_1084 = {1{`RANDOM}};
  btb_271_valid = _RAND_1084[0:0];
  _RAND_1085 = {1{`RANDOM}};
  btb_271_tag = _RAND_1085[9:0];
  _RAND_1086 = {2{`RANDOM}};
  btb_271_target_address = _RAND_1086[63:0];
  _RAND_1087 = {1{`RANDOM}};
  btb_271_bht = _RAND_1087[1:0];
  _RAND_1088 = {1{`RANDOM}};
  btb_272_valid = _RAND_1088[0:0];
  _RAND_1089 = {1{`RANDOM}};
  btb_272_tag = _RAND_1089[9:0];
  _RAND_1090 = {2{`RANDOM}};
  btb_272_target_address = _RAND_1090[63:0];
  _RAND_1091 = {1{`RANDOM}};
  btb_272_bht = _RAND_1091[1:0];
  _RAND_1092 = {1{`RANDOM}};
  btb_273_valid = _RAND_1092[0:0];
  _RAND_1093 = {1{`RANDOM}};
  btb_273_tag = _RAND_1093[9:0];
  _RAND_1094 = {2{`RANDOM}};
  btb_273_target_address = _RAND_1094[63:0];
  _RAND_1095 = {1{`RANDOM}};
  btb_273_bht = _RAND_1095[1:0];
  _RAND_1096 = {1{`RANDOM}};
  btb_274_valid = _RAND_1096[0:0];
  _RAND_1097 = {1{`RANDOM}};
  btb_274_tag = _RAND_1097[9:0];
  _RAND_1098 = {2{`RANDOM}};
  btb_274_target_address = _RAND_1098[63:0];
  _RAND_1099 = {1{`RANDOM}};
  btb_274_bht = _RAND_1099[1:0];
  _RAND_1100 = {1{`RANDOM}};
  btb_275_valid = _RAND_1100[0:0];
  _RAND_1101 = {1{`RANDOM}};
  btb_275_tag = _RAND_1101[9:0];
  _RAND_1102 = {2{`RANDOM}};
  btb_275_target_address = _RAND_1102[63:0];
  _RAND_1103 = {1{`RANDOM}};
  btb_275_bht = _RAND_1103[1:0];
  _RAND_1104 = {1{`RANDOM}};
  btb_276_valid = _RAND_1104[0:0];
  _RAND_1105 = {1{`RANDOM}};
  btb_276_tag = _RAND_1105[9:0];
  _RAND_1106 = {2{`RANDOM}};
  btb_276_target_address = _RAND_1106[63:0];
  _RAND_1107 = {1{`RANDOM}};
  btb_276_bht = _RAND_1107[1:0];
  _RAND_1108 = {1{`RANDOM}};
  btb_277_valid = _RAND_1108[0:0];
  _RAND_1109 = {1{`RANDOM}};
  btb_277_tag = _RAND_1109[9:0];
  _RAND_1110 = {2{`RANDOM}};
  btb_277_target_address = _RAND_1110[63:0];
  _RAND_1111 = {1{`RANDOM}};
  btb_277_bht = _RAND_1111[1:0];
  _RAND_1112 = {1{`RANDOM}};
  btb_278_valid = _RAND_1112[0:0];
  _RAND_1113 = {1{`RANDOM}};
  btb_278_tag = _RAND_1113[9:0];
  _RAND_1114 = {2{`RANDOM}};
  btb_278_target_address = _RAND_1114[63:0];
  _RAND_1115 = {1{`RANDOM}};
  btb_278_bht = _RAND_1115[1:0];
  _RAND_1116 = {1{`RANDOM}};
  btb_279_valid = _RAND_1116[0:0];
  _RAND_1117 = {1{`RANDOM}};
  btb_279_tag = _RAND_1117[9:0];
  _RAND_1118 = {2{`RANDOM}};
  btb_279_target_address = _RAND_1118[63:0];
  _RAND_1119 = {1{`RANDOM}};
  btb_279_bht = _RAND_1119[1:0];
  _RAND_1120 = {1{`RANDOM}};
  btb_280_valid = _RAND_1120[0:0];
  _RAND_1121 = {1{`RANDOM}};
  btb_280_tag = _RAND_1121[9:0];
  _RAND_1122 = {2{`RANDOM}};
  btb_280_target_address = _RAND_1122[63:0];
  _RAND_1123 = {1{`RANDOM}};
  btb_280_bht = _RAND_1123[1:0];
  _RAND_1124 = {1{`RANDOM}};
  btb_281_valid = _RAND_1124[0:0];
  _RAND_1125 = {1{`RANDOM}};
  btb_281_tag = _RAND_1125[9:0];
  _RAND_1126 = {2{`RANDOM}};
  btb_281_target_address = _RAND_1126[63:0];
  _RAND_1127 = {1{`RANDOM}};
  btb_281_bht = _RAND_1127[1:0];
  _RAND_1128 = {1{`RANDOM}};
  btb_282_valid = _RAND_1128[0:0];
  _RAND_1129 = {1{`RANDOM}};
  btb_282_tag = _RAND_1129[9:0];
  _RAND_1130 = {2{`RANDOM}};
  btb_282_target_address = _RAND_1130[63:0];
  _RAND_1131 = {1{`RANDOM}};
  btb_282_bht = _RAND_1131[1:0];
  _RAND_1132 = {1{`RANDOM}};
  btb_283_valid = _RAND_1132[0:0];
  _RAND_1133 = {1{`RANDOM}};
  btb_283_tag = _RAND_1133[9:0];
  _RAND_1134 = {2{`RANDOM}};
  btb_283_target_address = _RAND_1134[63:0];
  _RAND_1135 = {1{`RANDOM}};
  btb_283_bht = _RAND_1135[1:0];
  _RAND_1136 = {1{`RANDOM}};
  btb_284_valid = _RAND_1136[0:0];
  _RAND_1137 = {1{`RANDOM}};
  btb_284_tag = _RAND_1137[9:0];
  _RAND_1138 = {2{`RANDOM}};
  btb_284_target_address = _RAND_1138[63:0];
  _RAND_1139 = {1{`RANDOM}};
  btb_284_bht = _RAND_1139[1:0];
  _RAND_1140 = {1{`RANDOM}};
  btb_285_valid = _RAND_1140[0:0];
  _RAND_1141 = {1{`RANDOM}};
  btb_285_tag = _RAND_1141[9:0];
  _RAND_1142 = {2{`RANDOM}};
  btb_285_target_address = _RAND_1142[63:0];
  _RAND_1143 = {1{`RANDOM}};
  btb_285_bht = _RAND_1143[1:0];
  _RAND_1144 = {1{`RANDOM}};
  btb_286_valid = _RAND_1144[0:0];
  _RAND_1145 = {1{`RANDOM}};
  btb_286_tag = _RAND_1145[9:0];
  _RAND_1146 = {2{`RANDOM}};
  btb_286_target_address = _RAND_1146[63:0];
  _RAND_1147 = {1{`RANDOM}};
  btb_286_bht = _RAND_1147[1:0];
  _RAND_1148 = {1{`RANDOM}};
  btb_287_valid = _RAND_1148[0:0];
  _RAND_1149 = {1{`RANDOM}};
  btb_287_tag = _RAND_1149[9:0];
  _RAND_1150 = {2{`RANDOM}};
  btb_287_target_address = _RAND_1150[63:0];
  _RAND_1151 = {1{`RANDOM}};
  btb_287_bht = _RAND_1151[1:0];
  _RAND_1152 = {1{`RANDOM}};
  btb_288_valid = _RAND_1152[0:0];
  _RAND_1153 = {1{`RANDOM}};
  btb_288_tag = _RAND_1153[9:0];
  _RAND_1154 = {2{`RANDOM}};
  btb_288_target_address = _RAND_1154[63:0];
  _RAND_1155 = {1{`RANDOM}};
  btb_288_bht = _RAND_1155[1:0];
  _RAND_1156 = {1{`RANDOM}};
  btb_289_valid = _RAND_1156[0:0];
  _RAND_1157 = {1{`RANDOM}};
  btb_289_tag = _RAND_1157[9:0];
  _RAND_1158 = {2{`RANDOM}};
  btb_289_target_address = _RAND_1158[63:0];
  _RAND_1159 = {1{`RANDOM}};
  btb_289_bht = _RAND_1159[1:0];
  _RAND_1160 = {1{`RANDOM}};
  btb_290_valid = _RAND_1160[0:0];
  _RAND_1161 = {1{`RANDOM}};
  btb_290_tag = _RAND_1161[9:0];
  _RAND_1162 = {2{`RANDOM}};
  btb_290_target_address = _RAND_1162[63:0];
  _RAND_1163 = {1{`RANDOM}};
  btb_290_bht = _RAND_1163[1:0];
  _RAND_1164 = {1{`RANDOM}};
  btb_291_valid = _RAND_1164[0:0];
  _RAND_1165 = {1{`RANDOM}};
  btb_291_tag = _RAND_1165[9:0];
  _RAND_1166 = {2{`RANDOM}};
  btb_291_target_address = _RAND_1166[63:0];
  _RAND_1167 = {1{`RANDOM}};
  btb_291_bht = _RAND_1167[1:0];
  _RAND_1168 = {1{`RANDOM}};
  btb_292_valid = _RAND_1168[0:0];
  _RAND_1169 = {1{`RANDOM}};
  btb_292_tag = _RAND_1169[9:0];
  _RAND_1170 = {2{`RANDOM}};
  btb_292_target_address = _RAND_1170[63:0];
  _RAND_1171 = {1{`RANDOM}};
  btb_292_bht = _RAND_1171[1:0];
  _RAND_1172 = {1{`RANDOM}};
  btb_293_valid = _RAND_1172[0:0];
  _RAND_1173 = {1{`RANDOM}};
  btb_293_tag = _RAND_1173[9:0];
  _RAND_1174 = {2{`RANDOM}};
  btb_293_target_address = _RAND_1174[63:0];
  _RAND_1175 = {1{`RANDOM}};
  btb_293_bht = _RAND_1175[1:0];
  _RAND_1176 = {1{`RANDOM}};
  btb_294_valid = _RAND_1176[0:0];
  _RAND_1177 = {1{`RANDOM}};
  btb_294_tag = _RAND_1177[9:0];
  _RAND_1178 = {2{`RANDOM}};
  btb_294_target_address = _RAND_1178[63:0];
  _RAND_1179 = {1{`RANDOM}};
  btb_294_bht = _RAND_1179[1:0];
  _RAND_1180 = {1{`RANDOM}};
  btb_295_valid = _RAND_1180[0:0];
  _RAND_1181 = {1{`RANDOM}};
  btb_295_tag = _RAND_1181[9:0];
  _RAND_1182 = {2{`RANDOM}};
  btb_295_target_address = _RAND_1182[63:0];
  _RAND_1183 = {1{`RANDOM}};
  btb_295_bht = _RAND_1183[1:0];
  _RAND_1184 = {1{`RANDOM}};
  btb_296_valid = _RAND_1184[0:0];
  _RAND_1185 = {1{`RANDOM}};
  btb_296_tag = _RAND_1185[9:0];
  _RAND_1186 = {2{`RANDOM}};
  btb_296_target_address = _RAND_1186[63:0];
  _RAND_1187 = {1{`RANDOM}};
  btb_296_bht = _RAND_1187[1:0];
  _RAND_1188 = {1{`RANDOM}};
  btb_297_valid = _RAND_1188[0:0];
  _RAND_1189 = {1{`RANDOM}};
  btb_297_tag = _RAND_1189[9:0];
  _RAND_1190 = {2{`RANDOM}};
  btb_297_target_address = _RAND_1190[63:0];
  _RAND_1191 = {1{`RANDOM}};
  btb_297_bht = _RAND_1191[1:0];
  _RAND_1192 = {1{`RANDOM}};
  btb_298_valid = _RAND_1192[0:0];
  _RAND_1193 = {1{`RANDOM}};
  btb_298_tag = _RAND_1193[9:0];
  _RAND_1194 = {2{`RANDOM}};
  btb_298_target_address = _RAND_1194[63:0];
  _RAND_1195 = {1{`RANDOM}};
  btb_298_bht = _RAND_1195[1:0];
  _RAND_1196 = {1{`RANDOM}};
  btb_299_valid = _RAND_1196[0:0];
  _RAND_1197 = {1{`RANDOM}};
  btb_299_tag = _RAND_1197[9:0];
  _RAND_1198 = {2{`RANDOM}};
  btb_299_target_address = _RAND_1198[63:0];
  _RAND_1199 = {1{`RANDOM}};
  btb_299_bht = _RAND_1199[1:0];
  _RAND_1200 = {1{`RANDOM}};
  btb_300_valid = _RAND_1200[0:0];
  _RAND_1201 = {1{`RANDOM}};
  btb_300_tag = _RAND_1201[9:0];
  _RAND_1202 = {2{`RANDOM}};
  btb_300_target_address = _RAND_1202[63:0];
  _RAND_1203 = {1{`RANDOM}};
  btb_300_bht = _RAND_1203[1:0];
  _RAND_1204 = {1{`RANDOM}};
  btb_301_valid = _RAND_1204[0:0];
  _RAND_1205 = {1{`RANDOM}};
  btb_301_tag = _RAND_1205[9:0];
  _RAND_1206 = {2{`RANDOM}};
  btb_301_target_address = _RAND_1206[63:0];
  _RAND_1207 = {1{`RANDOM}};
  btb_301_bht = _RAND_1207[1:0];
  _RAND_1208 = {1{`RANDOM}};
  btb_302_valid = _RAND_1208[0:0];
  _RAND_1209 = {1{`RANDOM}};
  btb_302_tag = _RAND_1209[9:0];
  _RAND_1210 = {2{`RANDOM}};
  btb_302_target_address = _RAND_1210[63:0];
  _RAND_1211 = {1{`RANDOM}};
  btb_302_bht = _RAND_1211[1:0];
  _RAND_1212 = {1{`RANDOM}};
  btb_303_valid = _RAND_1212[0:0];
  _RAND_1213 = {1{`RANDOM}};
  btb_303_tag = _RAND_1213[9:0];
  _RAND_1214 = {2{`RANDOM}};
  btb_303_target_address = _RAND_1214[63:0];
  _RAND_1215 = {1{`RANDOM}};
  btb_303_bht = _RAND_1215[1:0];
  _RAND_1216 = {1{`RANDOM}};
  btb_304_valid = _RAND_1216[0:0];
  _RAND_1217 = {1{`RANDOM}};
  btb_304_tag = _RAND_1217[9:0];
  _RAND_1218 = {2{`RANDOM}};
  btb_304_target_address = _RAND_1218[63:0];
  _RAND_1219 = {1{`RANDOM}};
  btb_304_bht = _RAND_1219[1:0];
  _RAND_1220 = {1{`RANDOM}};
  btb_305_valid = _RAND_1220[0:0];
  _RAND_1221 = {1{`RANDOM}};
  btb_305_tag = _RAND_1221[9:0];
  _RAND_1222 = {2{`RANDOM}};
  btb_305_target_address = _RAND_1222[63:0];
  _RAND_1223 = {1{`RANDOM}};
  btb_305_bht = _RAND_1223[1:0];
  _RAND_1224 = {1{`RANDOM}};
  btb_306_valid = _RAND_1224[0:0];
  _RAND_1225 = {1{`RANDOM}};
  btb_306_tag = _RAND_1225[9:0];
  _RAND_1226 = {2{`RANDOM}};
  btb_306_target_address = _RAND_1226[63:0];
  _RAND_1227 = {1{`RANDOM}};
  btb_306_bht = _RAND_1227[1:0];
  _RAND_1228 = {1{`RANDOM}};
  btb_307_valid = _RAND_1228[0:0];
  _RAND_1229 = {1{`RANDOM}};
  btb_307_tag = _RAND_1229[9:0];
  _RAND_1230 = {2{`RANDOM}};
  btb_307_target_address = _RAND_1230[63:0];
  _RAND_1231 = {1{`RANDOM}};
  btb_307_bht = _RAND_1231[1:0];
  _RAND_1232 = {1{`RANDOM}};
  btb_308_valid = _RAND_1232[0:0];
  _RAND_1233 = {1{`RANDOM}};
  btb_308_tag = _RAND_1233[9:0];
  _RAND_1234 = {2{`RANDOM}};
  btb_308_target_address = _RAND_1234[63:0];
  _RAND_1235 = {1{`RANDOM}};
  btb_308_bht = _RAND_1235[1:0];
  _RAND_1236 = {1{`RANDOM}};
  btb_309_valid = _RAND_1236[0:0];
  _RAND_1237 = {1{`RANDOM}};
  btb_309_tag = _RAND_1237[9:0];
  _RAND_1238 = {2{`RANDOM}};
  btb_309_target_address = _RAND_1238[63:0];
  _RAND_1239 = {1{`RANDOM}};
  btb_309_bht = _RAND_1239[1:0];
  _RAND_1240 = {1{`RANDOM}};
  btb_310_valid = _RAND_1240[0:0];
  _RAND_1241 = {1{`RANDOM}};
  btb_310_tag = _RAND_1241[9:0];
  _RAND_1242 = {2{`RANDOM}};
  btb_310_target_address = _RAND_1242[63:0];
  _RAND_1243 = {1{`RANDOM}};
  btb_310_bht = _RAND_1243[1:0];
  _RAND_1244 = {1{`RANDOM}};
  btb_311_valid = _RAND_1244[0:0];
  _RAND_1245 = {1{`RANDOM}};
  btb_311_tag = _RAND_1245[9:0];
  _RAND_1246 = {2{`RANDOM}};
  btb_311_target_address = _RAND_1246[63:0];
  _RAND_1247 = {1{`RANDOM}};
  btb_311_bht = _RAND_1247[1:0];
  _RAND_1248 = {1{`RANDOM}};
  btb_312_valid = _RAND_1248[0:0];
  _RAND_1249 = {1{`RANDOM}};
  btb_312_tag = _RAND_1249[9:0];
  _RAND_1250 = {2{`RANDOM}};
  btb_312_target_address = _RAND_1250[63:0];
  _RAND_1251 = {1{`RANDOM}};
  btb_312_bht = _RAND_1251[1:0];
  _RAND_1252 = {1{`RANDOM}};
  btb_313_valid = _RAND_1252[0:0];
  _RAND_1253 = {1{`RANDOM}};
  btb_313_tag = _RAND_1253[9:0];
  _RAND_1254 = {2{`RANDOM}};
  btb_313_target_address = _RAND_1254[63:0];
  _RAND_1255 = {1{`RANDOM}};
  btb_313_bht = _RAND_1255[1:0];
  _RAND_1256 = {1{`RANDOM}};
  btb_314_valid = _RAND_1256[0:0];
  _RAND_1257 = {1{`RANDOM}};
  btb_314_tag = _RAND_1257[9:0];
  _RAND_1258 = {2{`RANDOM}};
  btb_314_target_address = _RAND_1258[63:0];
  _RAND_1259 = {1{`RANDOM}};
  btb_314_bht = _RAND_1259[1:0];
  _RAND_1260 = {1{`RANDOM}};
  btb_315_valid = _RAND_1260[0:0];
  _RAND_1261 = {1{`RANDOM}};
  btb_315_tag = _RAND_1261[9:0];
  _RAND_1262 = {2{`RANDOM}};
  btb_315_target_address = _RAND_1262[63:0];
  _RAND_1263 = {1{`RANDOM}};
  btb_315_bht = _RAND_1263[1:0];
  _RAND_1264 = {1{`RANDOM}};
  btb_316_valid = _RAND_1264[0:0];
  _RAND_1265 = {1{`RANDOM}};
  btb_316_tag = _RAND_1265[9:0];
  _RAND_1266 = {2{`RANDOM}};
  btb_316_target_address = _RAND_1266[63:0];
  _RAND_1267 = {1{`RANDOM}};
  btb_316_bht = _RAND_1267[1:0];
  _RAND_1268 = {1{`RANDOM}};
  btb_317_valid = _RAND_1268[0:0];
  _RAND_1269 = {1{`RANDOM}};
  btb_317_tag = _RAND_1269[9:0];
  _RAND_1270 = {2{`RANDOM}};
  btb_317_target_address = _RAND_1270[63:0];
  _RAND_1271 = {1{`RANDOM}};
  btb_317_bht = _RAND_1271[1:0];
  _RAND_1272 = {1{`RANDOM}};
  btb_318_valid = _RAND_1272[0:0];
  _RAND_1273 = {1{`RANDOM}};
  btb_318_tag = _RAND_1273[9:0];
  _RAND_1274 = {2{`RANDOM}};
  btb_318_target_address = _RAND_1274[63:0];
  _RAND_1275 = {1{`RANDOM}};
  btb_318_bht = _RAND_1275[1:0];
  _RAND_1276 = {1{`RANDOM}};
  btb_319_valid = _RAND_1276[0:0];
  _RAND_1277 = {1{`RANDOM}};
  btb_319_tag = _RAND_1277[9:0];
  _RAND_1278 = {2{`RANDOM}};
  btb_319_target_address = _RAND_1278[63:0];
  _RAND_1279 = {1{`RANDOM}};
  btb_319_bht = _RAND_1279[1:0];
  _RAND_1280 = {1{`RANDOM}};
  btb_320_valid = _RAND_1280[0:0];
  _RAND_1281 = {1{`RANDOM}};
  btb_320_tag = _RAND_1281[9:0];
  _RAND_1282 = {2{`RANDOM}};
  btb_320_target_address = _RAND_1282[63:0];
  _RAND_1283 = {1{`RANDOM}};
  btb_320_bht = _RAND_1283[1:0];
  _RAND_1284 = {1{`RANDOM}};
  btb_321_valid = _RAND_1284[0:0];
  _RAND_1285 = {1{`RANDOM}};
  btb_321_tag = _RAND_1285[9:0];
  _RAND_1286 = {2{`RANDOM}};
  btb_321_target_address = _RAND_1286[63:0];
  _RAND_1287 = {1{`RANDOM}};
  btb_321_bht = _RAND_1287[1:0];
  _RAND_1288 = {1{`RANDOM}};
  btb_322_valid = _RAND_1288[0:0];
  _RAND_1289 = {1{`RANDOM}};
  btb_322_tag = _RAND_1289[9:0];
  _RAND_1290 = {2{`RANDOM}};
  btb_322_target_address = _RAND_1290[63:0];
  _RAND_1291 = {1{`RANDOM}};
  btb_322_bht = _RAND_1291[1:0];
  _RAND_1292 = {1{`RANDOM}};
  btb_323_valid = _RAND_1292[0:0];
  _RAND_1293 = {1{`RANDOM}};
  btb_323_tag = _RAND_1293[9:0];
  _RAND_1294 = {2{`RANDOM}};
  btb_323_target_address = _RAND_1294[63:0];
  _RAND_1295 = {1{`RANDOM}};
  btb_323_bht = _RAND_1295[1:0];
  _RAND_1296 = {1{`RANDOM}};
  btb_324_valid = _RAND_1296[0:0];
  _RAND_1297 = {1{`RANDOM}};
  btb_324_tag = _RAND_1297[9:0];
  _RAND_1298 = {2{`RANDOM}};
  btb_324_target_address = _RAND_1298[63:0];
  _RAND_1299 = {1{`RANDOM}};
  btb_324_bht = _RAND_1299[1:0];
  _RAND_1300 = {1{`RANDOM}};
  btb_325_valid = _RAND_1300[0:0];
  _RAND_1301 = {1{`RANDOM}};
  btb_325_tag = _RAND_1301[9:0];
  _RAND_1302 = {2{`RANDOM}};
  btb_325_target_address = _RAND_1302[63:0];
  _RAND_1303 = {1{`RANDOM}};
  btb_325_bht = _RAND_1303[1:0];
  _RAND_1304 = {1{`RANDOM}};
  btb_326_valid = _RAND_1304[0:0];
  _RAND_1305 = {1{`RANDOM}};
  btb_326_tag = _RAND_1305[9:0];
  _RAND_1306 = {2{`RANDOM}};
  btb_326_target_address = _RAND_1306[63:0];
  _RAND_1307 = {1{`RANDOM}};
  btb_326_bht = _RAND_1307[1:0];
  _RAND_1308 = {1{`RANDOM}};
  btb_327_valid = _RAND_1308[0:0];
  _RAND_1309 = {1{`RANDOM}};
  btb_327_tag = _RAND_1309[9:0];
  _RAND_1310 = {2{`RANDOM}};
  btb_327_target_address = _RAND_1310[63:0];
  _RAND_1311 = {1{`RANDOM}};
  btb_327_bht = _RAND_1311[1:0];
  _RAND_1312 = {1{`RANDOM}};
  btb_328_valid = _RAND_1312[0:0];
  _RAND_1313 = {1{`RANDOM}};
  btb_328_tag = _RAND_1313[9:0];
  _RAND_1314 = {2{`RANDOM}};
  btb_328_target_address = _RAND_1314[63:0];
  _RAND_1315 = {1{`RANDOM}};
  btb_328_bht = _RAND_1315[1:0];
  _RAND_1316 = {1{`RANDOM}};
  btb_329_valid = _RAND_1316[0:0];
  _RAND_1317 = {1{`RANDOM}};
  btb_329_tag = _RAND_1317[9:0];
  _RAND_1318 = {2{`RANDOM}};
  btb_329_target_address = _RAND_1318[63:0];
  _RAND_1319 = {1{`RANDOM}};
  btb_329_bht = _RAND_1319[1:0];
  _RAND_1320 = {1{`RANDOM}};
  btb_330_valid = _RAND_1320[0:0];
  _RAND_1321 = {1{`RANDOM}};
  btb_330_tag = _RAND_1321[9:0];
  _RAND_1322 = {2{`RANDOM}};
  btb_330_target_address = _RAND_1322[63:0];
  _RAND_1323 = {1{`RANDOM}};
  btb_330_bht = _RAND_1323[1:0];
  _RAND_1324 = {1{`RANDOM}};
  btb_331_valid = _RAND_1324[0:0];
  _RAND_1325 = {1{`RANDOM}};
  btb_331_tag = _RAND_1325[9:0];
  _RAND_1326 = {2{`RANDOM}};
  btb_331_target_address = _RAND_1326[63:0];
  _RAND_1327 = {1{`RANDOM}};
  btb_331_bht = _RAND_1327[1:0];
  _RAND_1328 = {1{`RANDOM}};
  btb_332_valid = _RAND_1328[0:0];
  _RAND_1329 = {1{`RANDOM}};
  btb_332_tag = _RAND_1329[9:0];
  _RAND_1330 = {2{`RANDOM}};
  btb_332_target_address = _RAND_1330[63:0];
  _RAND_1331 = {1{`RANDOM}};
  btb_332_bht = _RAND_1331[1:0];
  _RAND_1332 = {1{`RANDOM}};
  btb_333_valid = _RAND_1332[0:0];
  _RAND_1333 = {1{`RANDOM}};
  btb_333_tag = _RAND_1333[9:0];
  _RAND_1334 = {2{`RANDOM}};
  btb_333_target_address = _RAND_1334[63:0];
  _RAND_1335 = {1{`RANDOM}};
  btb_333_bht = _RAND_1335[1:0];
  _RAND_1336 = {1{`RANDOM}};
  btb_334_valid = _RAND_1336[0:0];
  _RAND_1337 = {1{`RANDOM}};
  btb_334_tag = _RAND_1337[9:0];
  _RAND_1338 = {2{`RANDOM}};
  btb_334_target_address = _RAND_1338[63:0];
  _RAND_1339 = {1{`RANDOM}};
  btb_334_bht = _RAND_1339[1:0];
  _RAND_1340 = {1{`RANDOM}};
  btb_335_valid = _RAND_1340[0:0];
  _RAND_1341 = {1{`RANDOM}};
  btb_335_tag = _RAND_1341[9:0];
  _RAND_1342 = {2{`RANDOM}};
  btb_335_target_address = _RAND_1342[63:0];
  _RAND_1343 = {1{`RANDOM}};
  btb_335_bht = _RAND_1343[1:0];
  _RAND_1344 = {1{`RANDOM}};
  btb_336_valid = _RAND_1344[0:0];
  _RAND_1345 = {1{`RANDOM}};
  btb_336_tag = _RAND_1345[9:0];
  _RAND_1346 = {2{`RANDOM}};
  btb_336_target_address = _RAND_1346[63:0];
  _RAND_1347 = {1{`RANDOM}};
  btb_336_bht = _RAND_1347[1:0];
  _RAND_1348 = {1{`RANDOM}};
  btb_337_valid = _RAND_1348[0:0];
  _RAND_1349 = {1{`RANDOM}};
  btb_337_tag = _RAND_1349[9:0];
  _RAND_1350 = {2{`RANDOM}};
  btb_337_target_address = _RAND_1350[63:0];
  _RAND_1351 = {1{`RANDOM}};
  btb_337_bht = _RAND_1351[1:0];
  _RAND_1352 = {1{`RANDOM}};
  btb_338_valid = _RAND_1352[0:0];
  _RAND_1353 = {1{`RANDOM}};
  btb_338_tag = _RAND_1353[9:0];
  _RAND_1354 = {2{`RANDOM}};
  btb_338_target_address = _RAND_1354[63:0];
  _RAND_1355 = {1{`RANDOM}};
  btb_338_bht = _RAND_1355[1:0];
  _RAND_1356 = {1{`RANDOM}};
  btb_339_valid = _RAND_1356[0:0];
  _RAND_1357 = {1{`RANDOM}};
  btb_339_tag = _RAND_1357[9:0];
  _RAND_1358 = {2{`RANDOM}};
  btb_339_target_address = _RAND_1358[63:0];
  _RAND_1359 = {1{`RANDOM}};
  btb_339_bht = _RAND_1359[1:0];
  _RAND_1360 = {1{`RANDOM}};
  btb_340_valid = _RAND_1360[0:0];
  _RAND_1361 = {1{`RANDOM}};
  btb_340_tag = _RAND_1361[9:0];
  _RAND_1362 = {2{`RANDOM}};
  btb_340_target_address = _RAND_1362[63:0];
  _RAND_1363 = {1{`RANDOM}};
  btb_340_bht = _RAND_1363[1:0];
  _RAND_1364 = {1{`RANDOM}};
  btb_341_valid = _RAND_1364[0:0];
  _RAND_1365 = {1{`RANDOM}};
  btb_341_tag = _RAND_1365[9:0];
  _RAND_1366 = {2{`RANDOM}};
  btb_341_target_address = _RAND_1366[63:0];
  _RAND_1367 = {1{`RANDOM}};
  btb_341_bht = _RAND_1367[1:0];
  _RAND_1368 = {1{`RANDOM}};
  btb_342_valid = _RAND_1368[0:0];
  _RAND_1369 = {1{`RANDOM}};
  btb_342_tag = _RAND_1369[9:0];
  _RAND_1370 = {2{`RANDOM}};
  btb_342_target_address = _RAND_1370[63:0];
  _RAND_1371 = {1{`RANDOM}};
  btb_342_bht = _RAND_1371[1:0];
  _RAND_1372 = {1{`RANDOM}};
  btb_343_valid = _RAND_1372[0:0];
  _RAND_1373 = {1{`RANDOM}};
  btb_343_tag = _RAND_1373[9:0];
  _RAND_1374 = {2{`RANDOM}};
  btb_343_target_address = _RAND_1374[63:0];
  _RAND_1375 = {1{`RANDOM}};
  btb_343_bht = _RAND_1375[1:0];
  _RAND_1376 = {1{`RANDOM}};
  btb_344_valid = _RAND_1376[0:0];
  _RAND_1377 = {1{`RANDOM}};
  btb_344_tag = _RAND_1377[9:0];
  _RAND_1378 = {2{`RANDOM}};
  btb_344_target_address = _RAND_1378[63:0];
  _RAND_1379 = {1{`RANDOM}};
  btb_344_bht = _RAND_1379[1:0];
  _RAND_1380 = {1{`RANDOM}};
  btb_345_valid = _RAND_1380[0:0];
  _RAND_1381 = {1{`RANDOM}};
  btb_345_tag = _RAND_1381[9:0];
  _RAND_1382 = {2{`RANDOM}};
  btb_345_target_address = _RAND_1382[63:0];
  _RAND_1383 = {1{`RANDOM}};
  btb_345_bht = _RAND_1383[1:0];
  _RAND_1384 = {1{`RANDOM}};
  btb_346_valid = _RAND_1384[0:0];
  _RAND_1385 = {1{`RANDOM}};
  btb_346_tag = _RAND_1385[9:0];
  _RAND_1386 = {2{`RANDOM}};
  btb_346_target_address = _RAND_1386[63:0];
  _RAND_1387 = {1{`RANDOM}};
  btb_346_bht = _RAND_1387[1:0];
  _RAND_1388 = {1{`RANDOM}};
  btb_347_valid = _RAND_1388[0:0];
  _RAND_1389 = {1{`RANDOM}};
  btb_347_tag = _RAND_1389[9:0];
  _RAND_1390 = {2{`RANDOM}};
  btb_347_target_address = _RAND_1390[63:0];
  _RAND_1391 = {1{`RANDOM}};
  btb_347_bht = _RAND_1391[1:0];
  _RAND_1392 = {1{`RANDOM}};
  btb_348_valid = _RAND_1392[0:0];
  _RAND_1393 = {1{`RANDOM}};
  btb_348_tag = _RAND_1393[9:0];
  _RAND_1394 = {2{`RANDOM}};
  btb_348_target_address = _RAND_1394[63:0];
  _RAND_1395 = {1{`RANDOM}};
  btb_348_bht = _RAND_1395[1:0];
  _RAND_1396 = {1{`RANDOM}};
  btb_349_valid = _RAND_1396[0:0];
  _RAND_1397 = {1{`RANDOM}};
  btb_349_tag = _RAND_1397[9:0];
  _RAND_1398 = {2{`RANDOM}};
  btb_349_target_address = _RAND_1398[63:0];
  _RAND_1399 = {1{`RANDOM}};
  btb_349_bht = _RAND_1399[1:0];
  _RAND_1400 = {1{`RANDOM}};
  btb_350_valid = _RAND_1400[0:0];
  _RAND_1401 = {1{`RANDOM}};
  btb_350_tag = _RAND_1401[9:0];
  _RAND_1402 = {2{`RANDOM}};
  btb_350_target_address = _RAND_1402[63:0];
  _RAND_1403 = {1{`RANDOM}};
  btb_350_bht = _RAND_1403[1:0];
  _RAND_1404 = {1{`RANDOM}};
  btb_351_valid = _RAND_1404[0:0];
  _RAND_1405 = {1{`RANDOM}};
  btb_351_tag = _RAND_1405[9:0];
  _RAND_1406 = {2{`RANDOM}};
  btb_351_target_address = _RAND_1406[63:0];
  _RAND_1407 = {1{`RANDOM}};
  btb_351_bht = _RAND_1407[1:0];
  _RAND_1408 = {1{`RANDOM}};
  btb_352_valid = _RAND_1408[0:0];
  _RAND_1409 = {1{`RANDOM}};
  btb_352_tag = _RAND_1409[9:0];
  _RAND_1410 = {2{`RANDOM}};
  btb_352_target_address = _RAND_1410[63:0];
  _RAND_1411 = {1{`RANDOM}};
  btb_352_bht = _RAND_1411[1:0];
  _RAND_1412 = {1{`RANDOM}};
  btb_353_valid = _RAND_1412[0:0];
  _RAND_1413 = {1{`RANDOM}};
  btb_353_tag = _RAND_1413[9:0];
  _RAND_1414 = {2{`RANDOM}};
  btb_353_target_address = _RAND_1414[63:0];
  _RAND_1415 = {1{`RANDOM}};
  btb_353_bht = _RAND_1415[1:0];
  _RAND_1416 = {1{`RANDOM}};
  btb_354_valid = _RAND_1416[0:0];
  _RAND_1417 = {1{`RANDOM}};
  btb_354_tag = _RAND_1417[9:0];
  _RAND_1418 = {2{`RANDOM}};
  btb_354_target_address = _RAND_1418[63:0];
  _RAND_1419 = {1{`RANDOM}};
  btb_354_bht = _RAND_1419[1:0];
  _RAND_1420 = {1{`RANDOM}};
  btb_355_valid = _RAND_1420[0:0];
  _RAND_1421 = {1{`RANDOM}};
  btb_355_tag = _RAND_1421[9:0];
  _RAND_1422 = {2{`RANDOM}};
  btb_355_target_address = _RAND_1422[63:0];
  _RAND_1423 = {1{`RANDOM}};
  btb_355_bht = _RAND_1423[1:0];
  _RAND_1424 = {1{`RANDOM}};
  btb_356_valid = _RAND_1424[0:0];
  _RAND_1425 = {1{`RANDOM}};
  btb_356_tag = _RAND_1425[9:0];
  _RAND_1426 = {2{`RANDOM}};
  btb_356_target_address = _RAND_1426[63:0];
  _RAND_1427 = {1{`RANDOM}};
  btb_356_bht = _RAND_1427[1:0];
  _RAND_1428 = {1{`RANDOM}};
  btb_357_valid = _RAND_1428[0:0];
  _RAND_1429 = {1{`RANDOM}};
  btb_357_tag = _RAND_1429[9:0];
  _RAND_1430 = {2{`RANDOM}};
  btb_357_target_address = _RAND_1430[63:0];
  _RAND_1431 = {1{`RANDOM}};
  btb_357_bht = _RAND_1431[1:0];
  _RAND_1432 = {1{`RANDOM}};
  btb_358_valid = _RAND_1432[0:0];
  _RAND_1433 = {1{`RANDOM}};
  btb_358_tag = _RAND_1433[9:0];
  _RAND_1434 = {2{`RANDOM}};
  btb_358_target_address = _RAND_1434[63:0];
  _RAND_1435 = {1{`RANDOM}};
  btb_358_bht = _RAND_1435[1:0];
  _RAND_1436 = {1{`RANDOM}};
  btb_359_valid = _RAND_1436[0:0];
  _RAND_1437 = {1{`RANDOM}};
  btb_359_tag = _RAND_1437[9:0];
  _RAND_1438 = {2{`RANDOM}};
  btb_359_target_address = _RAND_1438[63:0];
  _RAND_1439 = {1{`RANDOM}};
  btb_359_bht = _RAND_1439[1:0];
  _RAND_1440 = {1{`RANDOM}};
  btb_360_valid = _RAND_1440[0:0];
  _RAND_1441 = {1{`RANDOM}};
  btb_360_tag = _RAND_1441[9:0];
  _RAND_1442 = {2{`RANDOM}};
  btb_360_target_address = _RAND_1442[63:0];
  _RAND_1443 = {1{`RANDOM}};
  btb_360_bht = _RAND_1443[1:0];
  _RAND_1444 = {1{`RANDOM}};
  btb_361_valid = _RAND_1444[0:0];
  _RAND_1445 = {1{`RANDOM}};
  btb_361_tag = _RAND_1445[9:0];
  _RAND_1446 = {2{`RANDOM}};
  btb_361_target_address = _RAND_1446[63:0];
  _RAND_1447 = {1{`RANDOM}};
  btb_361_bht = _RAND_1447[1:0];
  _RAND_1448 = {1{`RANDOM}};
  btb_362_valid = _RAND_1448[0:0];
  _RAND_1449 = {1{`RANDOM}};
  btb_362_tag = _RAND_1449[9:0];
  _RAND_1450 = {2{`RANDOM}};
  btb_362_target_address = _RAND_1450[63:0];
  _RAND_1451 = {1{`RANDOM}};
  btb_362_bht = _RAND_1451[1:0];
  _RAND_1452 = {1{`RANDOM}};
  btb_363_valid = _RAND_1452[0:0];
  _RAND_1453 = {1{`RANDOM}};
  btb_363_tag = _RAND_1453[9:0];
  _RAND_1454 = {2{`RANDOM}};
  btb_363_target_address = _RAND_1454[63:0];
  _RAND_1455 = {1{`RANDOM}};
  btb_363_bht = _RAND_1455[1:0];
  _RAND_1456 = {1{`RANDOM}};
  btb_364_valid = _RAND_1456[0:0];
  _RAND_1457 = {1{`RANDOM}};
  btb_364_tag = _RAND_1457[9:0];
  _RAND_1458 = {2{`RANDOM}};
  btb_364_target_address = _RAND_1458[63:0];
  _RAND_1459 = {1{`RANDOM}};
  btb_364_bht = _RAND_1459[1:0];
  _RAND_1460 = {1{`RANDOM}};
  btb_365_valid = _RAND_1460[0:0];
  _RAND_1461 = {1{`RANDOM}};
  btb_365_tag = _RAND_1461[9:0];
  _RAND_1462 = {2{`RANDOM}};
  btb_365_target_address = _RAND_1462[63:0];
  _RAND_1463 = {1{`RANDOM}};
  btb_365_bht = _RAND_1463[1:0];
  _RAND_1464 = {1{`RANDOM}};
  btb_366_valid = _RAND_1464[0:0];
  _RAND_1465 = {1{`RANDOM}};
  btb_366_tag = _RAND_1465[9:0];
  _RAND_1466 = {2{`RANDOM}};
  btb_366_target_address = _RAND_1466[63:0];
  _RAND_1467 = {1{`RANDOM}};
  btb_366_bht = _RAND_1467[1:0];
  _RAND_1468 = {1{`RANDOM}};
  btb_367_valid = _RAND_1468[0:0];
  _RAND_1469 = {1{`RANDOM}};
  btb_367_tag = _RAND_1469[9:0];
  _RAND_1470 = {2{`RANDOM}};
  btb_367_target_address = _RAND_1470[63:0];
  _RAND_1471 = {1{`RANDOM}};
  btb_367_bht = _RAND_1471[1:0];
  _RAND_1472 = {1{`RANDOM}};
  btb_368_valid = _RAND_1472[0:0];
  _RAND_1473 = {1{`RANDOM}};
  btb_368_tag = _RAND_1473[9:0];
  _RAND_1474 = {2{`RANDOM}};
  btb_368_target_address = _RAND_1474[63:0];
  _RAND_1475 = {1{`RANDOM}};
  btb_368_bht = _RAND_1475[1:0];
  _RAND_1476 = {1{`RANDOM}};
  btb_369_valid = _RAND_1476[0:0];
  _RAND_1477 = {1{`RANDOM}};
  btb_369_tag = _RAND_1477[9:0];
  _RAND_1478 = {2{`RANDOM}};
  btb_369_target_address = _RAND_1478[63:0];
  _RAND_1479 = {1{`RANDOM}};
  btb_369_bht = _RAND_1479[1:0];
  _RAND_1480 = {1{`RANDOM}};
  btb_370_valid = _RAND_1480[0:0];
  _RAND_1481 = {1{`RANDOM}};
  btb_370_tag = _RAND_1481[9:0];
  _RAND_1482 = {2{`RANDOM}};
  btb_370_target_address = _RAND_1482[63:0];
  _RAND_1483 = {1{`RANDOM}};
  btb_370_bht = _RAND_1483[1:0];
  _RAND_1484 = {1{`RANDOM}};
  btb_371_valid = _RAND_1484[0:0];
  _RAND_1485 = {1{`RANDOM}};
  btb_371_tag = _RAND_1485[9:0];
  _RAND_1486 = {2{`RANDOM}};
  btb_371_target_address = _RAND_1486[63:0];
  _RAND_1487 = {1{`RANDOM}};
  btb_371_bht = _RAND_1487[1:0];
  _RAND_1488 = {1{`RANDOM}};
  btb_372_valid = _RAND_1488[0:0];
  _RAND_1489 = {1{`RANDOM}};
  btb_372_tag = _RAND_1489[9:0];
  _RAND_1490 = {2{`RANDOM}};
  btb_372_target_address = _RAND_1490[63:0];
  _RAND_1491 = {1{`RANDOM}};
  btb_372_bht = _RAND_1491[1:0];
  _RAND_1492 = {1{`RANDOM}};
  btb_373_valid = _RAND_1492[0:0];
  _RAND_1493 = {1{`RANDOM}};
  btb_373_tag = _RAND_1493[9:0];
  _RAND_1494 = {2{`RANDOM}};
  btb_373_target_address = _RAND_1494[63:0];
  _RAND_1495 = {1{`RANDOM}};
  btb_373_bht = _RAND_1495[1:0];
  _RAND_1496 = {1{`RANDOM}};
  btb_374_valid = _RAND_1496[0:0];
  _RAND_1497 = {1{`RANDOM}};
  btb_374_tag = _RAND_1497[9:0];
  _RAND_1498 = {2{`RANDOM}};
  btb_374_target_address = _RAND_1498[63:0];
  _RAND_1499 = {1{`RANDOM}};
  btb_374_bht = _RAND_1499[1:0];
  _RAND_1500 = {1{`RANDOM}};
  btb_375_valid = _RAND_1500[0:0];
  _RAND_1501 = {1{`RANDOM}};
  btb_375_tag = _RAND_1501[9:0];
  _RAND_1502 = {2{`RANDOM}};
  btb_375_target_address = _RAND_1502[63:0];
  _RAND_1503 = {1{`RANDOM}};
  btb_375_bht = _RAND_1503[1:0];
  _RAND_1504 = {1{`RANDOM}};
  btb_376_valid = _RAND_1504[0:0];
  _RAND_1505 = {1{`RANDOM}};
  btb_376_tag = _RAND_1505[9:0];
  _RAND_1506 = {2{`RANDOM}};
  btb_376_target_address = _RAND_1506[63:0];
  _RAND_1507 = {1{`RANDOM}};
  btb_376_bht = _RAND_1507[1:0];
  _RAND_1508 = {1{`RANDOM}};
  btb_377_valid = _RAND_1508[0:0];
  _RAND_1509 = {1{`RANDOM}};
  btb_377_tag = _RAND_1509[9:0];
  _RAND_1510 = {2{`RANDOM}};
  btb_377_target_address = _RAND_1510[63:0];
  _RAND_1511 = {1{`RANDOM}};
  btb_377_bht = _RAND_1511[1:0];
  _RAND_1512 = {1{`RANDOM}};
  btb_378_valid = _RAND_1512[0:0];
  _RAND_1513 = {1{`RANDOM}};
  btb_378_tag = _RAND_1513[9:0];
  _RAND_1514 = {2{`RANDOM}};
  btb_378_target_address = _RAND_1514[63:0];
  _RAND_1515 = {1{`RANDOM}};
  btb_378_bht = _RAND_1515[1:0];
  _RAND_1516 = {1{`RANDOM}};
  btb_379_valid = _RAND_1516[0:0];
  _RAND_1517 = {1{`RANDOM}};
  btb_379_tag = _RAND_1517[9:0];
  _RAND_1518 = {2{`RANDOM}};
  btb_379_target_address = _RAND_1518[63:0];
  _RAND_1519 = {1{`RANDOM}};
  btb_379_bht = _RAND_1519[1:0];
  _RAND_1520 = {1{`RANDOM}};
  btb_380_valid = _RAND_1520[0:0];
  _RAND_1521 = {1{`RANDOM}};
  btb_380_tag = _RAND_1521[9:0];
  _RAND_1522 = {2{`RANDOM}};
  btb_380_target_address = _RAND_1522[63:0];
  _RAND_1523 = {1{`RANDOM}};
  btb_380_bht = _RAND_1523[1:0];
  _RAND_1524 = {1{`RANDOM}};
  btb_381_valid = _RAND_1524[0:0];
  _RAND_1525 = {1{`RANDOM}};
  btb_381_tag = _RAND_1525[9:0];
  _RAND_1526 = {2{`RANDOM}};
  btb_381_target_address = _RAND_1526[63:0];
  _RAND_1527 = {1{`RANDOM}};
  btb_381_bht = _RAND_1527[1:0];
  _RAND_1528 = {1{`RANDOM}};
  btb_382_valid = _RAND_1528[0:0];
  _RAND_1529 = {1{`RANDOM}};
  btb_382_tag = _RAND_1529[9:0];
  _RAND_1530 = {2{`RANDOM}};
  btb_382_target_address = _RAND_1530[63:0];
  _RAND_1531 = {1{`RANDOM}};
  btb_382_bht = _RAND_1531[1:0];
  _RAND_1532 = {1{`RANDOM}};
  btb_383_valid = _RAND_1532[0:0];
  _RAND_1533 = {1{`RANDOM}};
  btb_383_tag = _RAND_1533[9:0];
  _RAND_1534 = {2{`RANDOM}};
  btb_383_target_address = _RAND_1534[63:0];
  _RAND_1535 = {1{`RANDOM}};
  btb_383_bht = _RAND_1535[1:0];
  _RAND_1536 = {1{`RANDOM}};
  btb_384_valid = _RAND_1536[0:0];
  _RAND_1537 = {1{`RANDOM}};
  btb_384_tag = _RAND_1537[9:0];
  _RAND_1538 = {2{`RANDOM}};
  btb_384_target_address = _RAND_1538[63:0];
  _RAND_1539 = {1{`RANDOM}};
  btb_384_bht = _RAND_1539[1:0];
  _RAND_1540 = {1{`RANDOM}};
  btb_385_valid = _RAND_1540[0:0];
  _RAND_1541 = {1{`RANDOM}};
  btb_385_tag = _RAND_1541[9:0];
  _RAND_1542 = {2{`RANDOM}};
  btb_385_target_address = _RAND_1542[63:0];
  _RAND_1543 = {1{`RANDOM}};
  btb_385_bht = _RAND_1543[1:0];
  _RAND_1544 = {1{`RANDOM}};
  btb_386_valid = _RAND_1544[0:0];
  _RAND_1545 = {1{`RANDOM}};
  btb_386_tag = _RAND_1545[9:0];
  _RAND_1546 = {2{`RANDOM}};
  btb_386_target_address = _RAND_1546[63:0];
  _RAND_1547 = {1{`RANDOM}};
  btb_386_bht = _RAND_1547[1:0];
  _RAND_1548 = {1{`RANDOM}};
  btb_387_valid = _RAND_1548[0:0];
  _RAND_1549 = {1{`RANDOM}};
  btb_387_tag = _RAND_1549[9:0];
  _RAND_1550 = {2{`RANDOM}};
  btb_387_target_address = _RAND_1550[63:0];
  _RAND_1551 = {1{`RANDOM}};
  btb_387_bht = _RAND_1551[1:0];
  _RAND_1552 = {1{`RANDOM}};
  btb_388_valid = _RAND_1552[0:0];
  _RAND_1553 = {1{`RANDOM}};
  btb_388_tag = _RAND_1553[9:0];
  _RAND_1554 = {2{`RANDOM}};
  btb_388_target_address = _RAND_1554[63:0];
  _RAND_1555 = {1{`RANDOM}};
  btb_388_bht = _RAND_1555[1:0];
  _RAND_1556 = {1{`RANDOM}};
  btb_389_valid = _RAND_1556[0:0];
  _RAND_1557 = {1{`RANDOM}};
  btb_389_tag = _RAND_1557[9:0];
  _RAND_1558 = {2{`RANDOM}};
  btb_389_target_address = _RAND_1558[63:0];
  _RAND_1559 = {1{`RANDOM}};
  btb_389_bht = _RAND_1559[1:0];
  _RAND_1560 = {1{`RANDOM}};
  btb_390_valid = _RAND_1560[0:0];
  _RAND_1561 = {1{`RANDOM}};
  btb_390_tag = _RAND_1561[9:0];
  _RAND_1562 = {2{`RANDOM}};
  btb_390_target_address = _RAND_1562[63:0];
  _RAND_1563 = {1{`RANDOM}};
  btb_390_bht = _RAND_1563[1:0];
  _RAND_1564 = {1{`RANDOM}};
  btb_391_valid = _RAND_1564[0:0];
  _RAND_1565 = {1{`RANDOM}};
  btb_391_tag = _RAND_1565[9:0];
  _RAND_1566 = {2{`RANDOM}};
  btb_391_target_address = _RAND_1566[63:0];
  _RAND_1567 = {1{`RANDOM}};
  btb_391_bht = _RAND_1567[1:0];
  _RAND_1568 = {1{`RANDOM}};
  btb_392_valid = _RAND_1568[0:0];
  _RAND_1569 = {1{`RANDOM}};
  btb_392_tag = _RAND_1569[9:0];
  _RAND_1570 = {2{`RANDOM}};
  btb_392_target_address = _RAND_1570[63:0];
  _RAND_1571 = {1{`RANDOM}};
  btb_392_bht = _RAND_1571[1:0];
  _RAND_1572 = {1{`RANDOM}};
  btb_393_valid = _RAND_1572[0:0];
  _RAND_1573 = {1{`RANDOM}};
  btb_393_tag = _RAND_1573[9:0];
  _RAND_1574 = {2{`RANDOM}};
  btb_393_target_address = _RAND_1574[63:0];
  _RAND_1575 = {1{`RANDOM}};
  btb_393_bht = _RAND_1575[1:0];
  _RAND_1576 = {1{`RANDOM}};
  btb_394_valid = _RAND_1576[0:0];
  _RAND_1577 = {1{`RANDOM}};
  btb_394_tag = _RAND_1577[9:0];
  _RAND_1578 = {2{`RANDOM}};
  btb_394_target_address = _RAND_1578[63:0];
  _RAND_1579 = {1{`RANDOM}};
  btb_394_bht = _RAND_1579[1:0];
  _RAND_1580 = {1{`RANDOM}};
  btb_395_valid = _RAND_1580[0:0];
  _RAND_1581 = {1{`RANDOM}};
  btb_395_tag = _RAND_1581[9:0];
  _RAND_1582 = {2{`RANDOM}};
  btb_395_target_address = _RAND_1582[63:0];
  _RAND_1583 = {1{`RANDOM}};
  btb_395_bht = _RAND_1583[1:0];
  _RAND_1584 = {1{`RANDOM}};
  btb_396_valid = _RAND_1584[0:0];
  _RAND_1585 = {1{`RANDOM}};
  btb_396_tag = _RAND_1585[9:0];
  _RAND_1586 = {2{`RANDOM}};
  btb_396_target_address = _RAND_1586[63:0];
  _RAND_1587 = {1{`RANDOM}};
  btb_396_bht = _RAND_1587[1:0];
  _RAND_1588 = {1{`RANDOM}};
  btb_397_valid = _RAND_1588[0:0];
  _RAND_1589 = {1{`RANDOM}};
  btb_397_tag = _RAND_1589[9:0];
  _RAND_1590 = {2{`RANDOM}};
  btb_397_target_address = _RAND_1590[63:0];
  _RAND_1591 = {1{`RANDOM}};
  btb_397_bht = _RAND_1591[1:0];
  _RAND_1592 = {1{`RANDOM}};
  btb_398_valid = _RAND_1592[0:0];
  _RAND_1593 = {1{`RANDOM}};
  btb_398_tag = _RAND_1593[9:0];
  _RAND_1594 = {2{`RANDOM}};
  btb_398_target_address = _RAND_1594[63:0];
  _RAND_1595 = {1{`RANDOM}};
  btb_398_bht = _RAND_1595[1:0];
  _RAND_1596 = {1{`RANDOM}};
  btb_399_valid = _RAND_1596[0:0];
  _RAND_1597 = {1{`RANDOM}};
  btb_399_tag = _RAND_1597[9:0];
  _RAND_1598 = {2{`RANDOM}};
  btb_399_target_address = _RAND_1598[63:0];
  _RAND_1599 = {1{`RANDOM}};
  btb_399_bht = _RAND_1599[1:0];
  _RAND_1600 = {1{`RANDOM}};
  btb_400_valid = _RAND_1600[0:0];
  _RAND_1601 = {1{`RANDOM}};
  btb_400_tag = _RAND_1601[9:0];
  _RAND_1602 = {2{`RANDOM}};
  btb_400_target_address = _RAND_1602[63:0];
  _RAND_1603 = {1{`RANDOM}};
  btb_400_bht = _RAND_1603[1:0];
  _RAND_1604 = {1{`RANDOM}};
  btb_401_valid = _RAND_1604[0:0];
  _RAND_1605 = {1{`RANDOM}};
  btb_401_tag = _RAND_1605[9:0];
  _RAND_1606 = {2{`RANDOM}};
  btb_401_target_address = _RAND_1606[63:0];
  _RAND_1607 = {1{`RANDOM}};
  btb_401_bht = _RAND_1607[1:0];
  _RAND_1608 = {1{`RANDOM}};
  btb_402_valid = _RAND_1608[0:0];
  _RAND_1609 = {1{`RANDOM}};
  btb_402_tag = _RAND_1609[9:0];
  _RAND_1610 = {2{`RANDOM}};
  btb_402_target_address = _RAND_1610[63:0];
  _RAND_1611 = {1{`RANDOM}};
  btb_402_bht = _RAND_1611[1:0];
  _RAND_1612 = {1{`RANDOM}};
  btb_403_valid = _RAND_1612[0:0];
  _RAND_1613 = {1{`RANDOM}};
  btb_403_tag = _RAND_1613[9:0];
  _RAND_1614 = {2{`RANDOM}};
  btb_403_target_address = _RAND_1614[63:0];
  _RAND_1615 = {1{`RANDOM}};
  btb_403_bht = _RAND_1615[1:0];
  _RAND_1616 = {1{`RANDOM}};
  btb_404_valid = _RAND_1616[0:0];
  _RAND_1617 = {1{`RANDOM}};
  btb_404_tag = _RAND_1617[9:0];
  _RAND_1618 = {2{`RANDOM}};
  btb_404_target_address = _RAND_1618[63:0];
  _RAND_1619 = {1{`RANDOM}};
  btb_404_bht = _RAND_1619[1:0];
  _RAND_1620 = {1{`RANDOM}};
  btb_405_valid = _RAND_1620[0:0];
  _RAND_1621 = {1{`RANDOM}};
  btb_405_tag = _RAND_1621[9:0];
  _RAND_1622 = {2{`RANDOM}};
  btb_405_target_address = _RAND_1622[63:0];
  _RAND_1623 = {1{`RANDOM}};
  btb_405_bht = _RAND_1623[1:0];
  _RAND_1624 = {1{`RANDOM}};
  btb_406_valid = _RAND_1624[0:0];
  _RAND_1625 = {1{`RANDOM}};
  btb_406_tag = _RAND_1625[9:0];
  _RAND_1626 = {2{`RANDOM}};
  btb_406_target_address = _RAND_1626[63:0];
  _RAND_1627 = {1{`RANDOM}};
  btb_406_bht = _RAND_1627[1:0];
  _RAND_1628 = {1{`RANDOM}};
  btb_407_valid = _RAND_1628[0:0];
  _RAND_1629 = {1{`RANDOM}};
  btb_407_tag = _RAND_1629[9:0];
  _RAND_1630 = {2{`RANDOM}};
  btb_407_target_address = _RAND_1630[63:0];
  _RAND_1631 = {1{`RANDOM}};
  btb_407_bht = _RAND_1631[1:0];
  _RAND_1632 = {1{`RANDOM}};
  btb_408_valid = _RAND_1632[0:0];
  _RAND_1633 = {1{`RANDOM}};
  btb_408_tag = _RAND_1633[9:0];
  _RAND_1634 = {2{`RANDOM}};
  btb_408_target_address = _RAND_1634[63:0];
  _RAND_1635 = {1{`RANDOM}};
  btb_408_bht = _RAND_1635[1:0];
  _RAND_1636 = {1{`RANDOM}};
  btb_409_valid = _RAND_1636[0:0];
  _RAND_1637 = {1{`RANDOM}};
  btb_409_tag = _RAND_1637[9:0];
  _RAND_1638 = {2{`RANDOM}};
  btb_409_target_address = _RAND_1638[63:0];
  _RAND_1639 = {1{`RANDOM}};
  btb_409_bht = _RAND_1639[1:0];
  _RAND_1640 = {1{`RANDOM}};
  btb_410_valid = _RAND_1640[0:0];
  _RAND_1641 = {1{`RANDOM}};
  btb_410_tag = _RAND_1641[9:0];
  _RAND_1642 = {2{`RANDOM}};
  btb_410_target_address = _RAND_1642[63:0];
  _RAND_1643 = {1{`RANDOM}};
  btb_410_bht = _RAND_1643[1:0];
  _RAND_1644 = {1{`RANDOM}};
  btb_411_valid = _RAND_1644[0:0];
  _RAND_1645 = {1{`RANDOM}};
  btb_411_tag = _RAND_1645[9:0];
  _RAND_1646 = {2{`RANDOM}};
  btb_411_target_address = _RAND_1646[63:0];
  _RAND_1647 = {1{`RANDOM}};
  btb_411_bht = _RAND_1647[1:0];
  _RAND_1648 = {1{`RANDOM}};
  btb_412_valid = _RAND_1648[0:0];
  _RAND_1649 = {1{`RANDOM}};
  btb_412_tag = _RAND_1649[9:0];
  _RAND_1650 = {2{`RANDOM}};
  btb_412_target_address = _RAND_1650[63:0];
  _RAND_1651 = {1{`RANDOM}};
  btb_412_bht = _RAND_1651[1:0];
  _RAND_1652 = {1{`RANDOM}};
  btb_413_valid = _RAND_1652[0:0];
  _RAND_1653 = {1{`RANDOM}};
  btb_413_tag = _RAND_1653[9:0];
  _RAND_1654 = {2{`RANDOM}};
  btb_413_target_address = _RAND_1654[63:0];
  _RAND_1655 = {1{`RANDOM}};
  btb_413_bht = _RAND_1655[1:0];
  _RAND_1656 = {1{`RANDOM}};
  btb_414_valid = _RAND_1656[0:0];
  _RAND_1657 = {1{`RANDOM}};
  btb_414_tag = _RAND_1657[9:0];
  _RAND_1658 = {2{`RANDOM}};
  btb_414_target_address = _RAND_1658[63:0];
  _RAND_1659 = {1{`RANDOM}};
  btb_414_bht = _RAND_1659[1:0];
  _RAND_1660 = {1{`RANDOM}};
  btb_415_valid = _RAND_1660[0:0];
  _RAND_1661 = {1{`RANDOM}};
  btb_415_tag = _RAND_1661[9:0];
  _RAND_1662 = {2{`RANDOM}};
  btb_415_target_address = _RAND_1662[63:0];
  _RAND_1663 = {1{`RANDOM}};
  btb_415_bht = _RAND_1663[1:0];
  _RAND_1664 = {1{`RANDOM}};
  btb_416_valid = _RAND_1664[0:0];
  _RAND_1665 = {1{`RANDOM}};
  btb_416_tag = _RAND_1665[9:0];
  _RAND_1666 = {2{`RANDOM}};
  btb_416_target_address = _RAND_1666[63:0];
  _RAND_1667 = {1{`RANDOM}};
  btb_416_bht = _RAND_1667[1:0];
  _RAND_1668 = {1{`RANDOM}};
  btb_417_valid = _RAND_1668[0:0];
  _RAND_1669 = {1{`RANDOM}};
  btb_417_tag = _RAND_1669[9:0];
  _RAND_1670 = {2{`RANDOM}};
  btb_417_target_address = _RAND_1670[63:0];
  _RAND_1671 = {1{`RANDOM}};
  btb_417_bht = _RAND_1671[1:0];
  _RAND_1672 = {1{`RANDOM}};
  btb_418_valid = _RAND_1672[0:0];
  _RAND_1673 = {1{`RANDOM}};
  btb_418_tag = _RAND_1673[9:0];
  _RAND_1674 = {2{`RANDOM}};
  btb_418_target_address = _RAND_1674[63:0];
  _RAND_1675 = {1{`RANDOM}};
  btb_418_bht = _RAND_1675[1:0];
  _RAND_1676 = {1{`RANDOM}};
  btb_419_valid = _RAND_1676[0:0];
  _RAND_1677 = {1{`RANDOM}};
  btb_419_tag = _RAND_1677[9:0];
  _RAND_1678 = {2{`RANDOM}};
  btb_419_target_address = _RAND_1678[63:0];
  _RAND_1679 = {1{`RANDOM}};
  btb_419_bht = _RAND_1679[1:0];
  _RAND_1680 = {1{`RANDOM}};
  btb_420_valid = _RAND_1680[0:0];
  _RAND_1681 = {1{`RANDOM}};
  btb_420_tag = _RAND_1681[9:0];
  _RAND_1682 = {2{`RANDOM}};
  btb_420_target_address = _RAND_1682[63:0];
  _RAND_1683 = {1{`RANDOM}};
  btb_420_bht = _RAND_1683[1:0];
  _RAND_1684 = {1{`RANDOM}};
  btb_421_valid = _RAND_1684[0:0];
  _RAND_1685 = {1{`RANDOM}};
  btb_421_tag = _RAND_1685[9:0];
  _RAND_1686 = {2{`RANDOM}};
  btb_421_target_address = _RAND_1686[63:0];
  _RAND_1687 = {1{`RANDOM}};
  btb_421_bht = _RAND_1687[1:0];
  _RAND_1688 = {1{`RANDOM}};
  btb_422_valid = _RAND_1688[0:0];
  _RAND_1689 = {1{`RANDOM}};
  btb_422_tag = _RAND_1689[9:0];
  _RAND_1690 = {2{`RANDOM}};
  btb_422_target_address = _RAND_1690[63:0];
  _RAND_1691 = {1{`RANDOM}};
  btb_422_bht = _RAND_1691[1:0];
  _RAND_1692 = {1{`RANDOM}};
  btb_423_valid = _RAND_1692[0:0];
  _RAND_1693 = {1{`RANDOM}};
  btb_423_tag = _RAND_1693[9:0];
  _RAND_1694 = {2{`RANDOM}};
  btb_423_target_address = _RAND_1694[63:0];
  _RAND_1695 = {1{`RANDOM}};
  btb_423_bht = _RAND_1695[1:0];
  _RAND_1696 = {1{`RANDOM}};
  btb_424_valid = _RAND_1696[0:0];
  _RAND_1697 = {1{`RANDOM}};
  btb_424_tag = _RAND_1697[9:0];
  _RAND_1698 = {2{`RANDOM}};
  btb_424_target_address = _RAND_1698[63:0];
  _RAND_1699 = {1{`RANDOM}};
  btb_424_bht = _RAND_1699[1:0];
  _RAND_1700 = {1{`RANDOM}};
  btb_425_valid = _RAND_1700[0:0];
  _RAND_1701 = {1{`RANDOM}};
  btb_425_tag = _RAND_1701[9:0];
  _RAND_1702 = {2{`RANDOM}};
  btb_425_target_address = _RAND_1702[63:0];
  _RAND_1703 = {1{`RANDOM}};
  btb_425_bht = _RAND_1703[1:0];
  _RAND_1704 = {1{`RANDOM}};
  btb_426_valid = _RAND_1704[0:0];
  _RAND_1705 = {1{`RANDOM}};
  btb_426_tag = _RAND_1705[9:0];
  _RAND_1706 = {2{`RANDOM}};
  btb_426_target_address = _RAND_1706[63:0];
  _RAND_1707 = {1{`RANDOM}};
  btb_426_bht = _RAND_1707[1:0];
  _RAND_1708 = {1{`RANDOM}};
  btb_427_valid = _RAND_1708[0:0];
  _RAND_1709 = {1{`RANDOM}};
  btb_427_tag = _RAND_1709[9:0];
  _RAND_1710 = {2{`RANDOM}};
  btb_427_target_address = _RAND_1710[63:0];
  _RAND_1711 = {1{`RANDOM}};
  btb_427_bht = _RAND_1711[1:0];
  _RAND_1712 = {1{`RANDOM}};
  btb_428_valid = _RAND_1712[0:0];
  _RAND_1713 = {1{`RANDOM}};
  btb_428_tag = _RAND_1713[9:0];
  _RAND_1714 = {2{`RANDOM}};
  btb_428_target_address = _RAND_1714[63:0];
  _RAND_1715 = {1{`RANDOM}};
  btb_428_bht = _RAND_1715[1:0];
  _RAND_1716 = {1{`RANDOM}};
  btb_429_valid = _RAND_1716[0:0];
  _RAND_1717 = {1{`RANDOM}};
  btb_429_tag = _RAND_1717[9:0];
  _RAND_1718 = {2{`RANDOM}};
  btb_429_target_address = _RAND_1718[63:0];
  _RAND_1719 = {1{`RANDOM}};
  btb_429_bht = _RAND_1719[1:0];
  _RAND_1720 = {1{`RANDOM}};
  btb_430_valid = _RAND_1720[0:0];
  _RAND_1721 = {1{`RANDOM}};
  btb_430_tag = _RAND_1721[9:0];
  _RAND_1722 = {2{`RANDOM}};
  btb_430_target_address = _RAND_1722[63:0];
  _RAND_1723 = {1{`RANDOM}};
  btb_430_bht = _RAND_1723[1:0];
  _RAND_1724 = {1{`RANDOM}};
  btb_431_valid = _RAND_1724[0:0];
  _RAND_1725 = {1{`RANDOM}};
  btb_431_tag = _RAND_1725[9:0];
  _RAND_1726 = {2{`RANDOM}};
  btb_431_target_address = _RAND_1726[63:0];
  _RAND_1727 = {1{`RANDOM}};
  btb_431_bht = _RAND_1727[1:0];
  _RAND_1728 = {1{`RANDOM}};
  btb_432_valid = _RAND_1728[0:0];
  _RAND_1729 = {1{`RANDOM}};
  btb_432_tag = _RAND_1729[9:0];
  _RAND_1730 = {2{`RANDOM}};
  btb_432_target_address = _RAND_1730[63:0];
  _RAND_1731 = {1{`RANDOM}};
  btb_432_bht = _RAND_1731[1:0];
  _RAND_1732 = {1{`RANDOM}};
  btb_433_valid = _RAND_1732[0:0];
  _RAND_1733 = {1{`RANDOM}};
  btb_433_tag = _RAND_1733[9:0];
  _RAND_1734 = {2{`RANDOM}};
  btb_433_target_address = _RAND_1734[63:0];
  _RAND_1735 = {1{`RANDOM}};
  btb_433_bht = _RAND_1735[1:0];
  _RAND_1736 = {1{`RANDOM}};
  btb_434_valid = _RAND_1736[0:0];
  _RAND_1737 = {1{`RANDOM}};
  btb_434_tag = _RAND_1737[9:0];
  _RAND_1738 = {2{`RANDOM}};
  btb_434_target_address = _RAND_1738[63:0];
  _RAND_1739 = {1{`RANDOM}};
  btb_434_bht = _RAND_1739[1:0];
  _RAND_1740 = {1{`RANDOM}};
  btb_435_valid = _RAND_1740[0:0];
  _RAND_1741 = {1{`RANDOM}};
  btb_435_tag = _RAND_1741[9:0];
  _RAND_1742 = {2{`RANDOM}};
  btb_435_target_address = _RAND_1742[63:0];
  _RAND_1743 = {1{`RANDOM}};
  btb_435_bht = _RAND_1743[1:0];
  _RAND_1744 = {1{`RANDOM}};
  btb_436_valid = _RAND_1744[0:0];
  _RAND_1745 = {1{`RANDOM}};
  btb_436_tag = _RAND_1745[9:0];
  _RAND_1746 = {2{`RANDOM}};
  btb_436_target_address = _RAND_1746[63:0];
  _RAND_1747 = {1{`RANDOM}};
  btb_436_bht = _RAND_1747[1:0];
  _RAND_1748 = {1{`RANDOM}};
  btb_437_valid = _RAND_1748[0:0];
  _RAND_1749 = {1{`RANDOM}};
  btb_437_tag = _RAND_1749[9:0];
  _RAND_1750 = {2{`RANDOM}};
  btb_437_target_address = _RAND_1750[63:0];
  _RAND_1751 = {1{`RANDOM}};
  btb_437_bht = _RAND_1751[1:0];
  _RAND_1752 = {1{`RANDOM}};
  btb_438_valid = _RAND_1752[0:0];
  _RAND_1753 = {1{`RANDOM}};
  btb_438_tag = _RAND_1753[9:0];
  _RAND_1754 = {2{`RANDOM}};
  btb_438_target_address = _RAND_1754[63:0];
  _RAND_1755 = {1{`RANDOM}};
  btb_438_bht = _RAND_1755[1:0];
  _RAND_1756 = {1{`RANDOM}};
  btb_439_valid = _RAND_1756[0:0];
  _RAND_1757 = {1{`RANDOM}};
  btb_439_tag = _RAND_1757[9:0];
  _RAND_1758 = {2{`RANDOM}};
  btb_439_target_address = _RAND_1758[63:0];
  _RAND_1759 = {1{`RANDOM}};
  btb_439_bht = _RAND_1759[1:0];
  _RAND_1760 = {1{`RANDOM}};
  btb_440_valid = _RAND_1760[0:0];
  _RAND_1761 = {1{`RANDOM}};
  btb_440_tag = _RAND_1761[9:0];
  _RAND_1762 = {2{`RANDOM}};
  btb_440_target_address = _RAND_1762[63:0];
  _RAND_1763 = {1{`RANDOM}};
  btb_440_bht = _RAND_1763[1:0];
  _RAND_1764 = {1{`RANDOM}};
  btb_441_valid = _RAND_1764[0:0];
  _RAND_1765 = {1{`RANDOM}};
  btb_441_tag = _RAND_1765[9:0];
  _RAND_1766 = {2{`RANDOM}};
  btb_441_target_address = _RAND_1766[63:0];
  _RAND_1767 = {1{`RANDOM}};
  btb_441_bht = _RAND_1767[1:0];
  _RAND_1768 = {1{`RANDOM}};
  btb_442_valid = _RAND_1768[0:0];
  _RAND_1769 = {1{`RANDOM}};
  btb_442_tag = _RAND_1769[9:0];
  _RAND_1770 = {2{`RANDOM}};
  btb_442_target_address = _RAND_1770[63:0];
  _RAND_1771 = {1{`RANDOM}};
  btb_442_bht = _RAND_1771[1:0];
  _RAND_1772 = {1{`RANDOM}};
  btb_443_valid = _RAND_1772[0:0];
  _RAND_1773 = {1{`RANDOM}};
  btb_443_tag = _RAND_1773[9:0];
  _RAND_1774 = {2{`RANDOM}};
  btb_443_target_address = _RAND_1774[63:0];
  _RAND_1775 = {1{`RANDOM}};
  btb_443_bht = _RAND_1775[1:0];
  _RAND_1776 = {1{`RANDOM}};
  btb_444_valid = _RAND_1776[0:0];
  _RAND_1777 = {1{`RANDOM}};
  btb_444_tag = _RAND_1777[9:0];
  _RAND_1778 = {2{`RANDOM}};
  btb_444_target_address = _RAND_1778[63:0];
  _RAND_1779 = {1{`RANDOM}};
  btb_444_bht = _RAND_1779[1:0];
  _RAND_1780 = {1{`RANDOM}};
  btb_445_valid = _RAND_1780[0:0];
  _RAND_1781 = {1{`RANDOM}};
  btb_445_tag = _RAND_1781[9:0];
  _RAND_1782 = {2{`RANDOM}};
  btb_445_target_address = _RAND_1782[63:0];
  _RAND_1783 = {1{`RANDOM}};
  btb_445_bht = _RAND_1783[1:0];
  _RAND_1784 = {1{`RANDOM}};
  btb_446_valid = _RAND_1784[0:0];
  _RAND_1785 = {1{`RANDOM}};
  btb_446_tag = _RAND_1785[9:0];
  _RAND_1786 = {2{`RANDOM}};
  btb_446_target_address = _RAND_1786[63:0];
  _RAND_1787 = {1{`RANDOM}};
  btb_446_bht = _RAND_1787[1:0];
  _RAND_1788 = {1{`RANDOM}};
  btb_447_valid = _RAND_1788[0:0];
  _RAND_1789 = {1{`RANDOM}};
  btb_447_tag = _RAND_1789[9:0];
  _RAND_1790 = {2{`RANDOM}};
  btb_447_target_address = _RAND_1790[63:0];
  _RAND_1791 = {1{`RANDOM}};
  btb_447_bht = _RAND_1791[1:0];
  _RAND_1792 = {1{`RANDOM}};
  btb_448_valid = _RAND_1792[0:0];
  _RAND_1793 = {1{`RANDOM}};
  btb_448_tag = _RAND_1793[9:0];
  _RAND_1794 = {2{`RANDOM}};
  btb_448_target_address = _RAND_1794[63:0];
  _RAND_1795 = {1{`RANDOM}};
  btb_448_bht = _RAND_1795[1:0];
  _RAND_1796 = {1{`RANDOM}};
  btb_449_valid = _RAND_1796[0:0];
  _RAND_1797 = {1{`RANDOM}};
  btb_449_tag = _RAND_1797[9:0];
  _RAND_1798 = {2{`RANDOM}};
  btb_449_target_address = _RAND_1798[63:0];
  _RAND_1799 = {1{`RANDOM}};
  btb_449_bht = _RAND_1799[1:0];
  _RAND_1800 = {1{`RANDOM}};
  btb_450_valid = _RAND_1800[0:0];
  _RAND_1801 = {1{`RANDOM}};
  btb_450_tag = _RAND_1801[9:0];
  _RAND_1802 = {2{`RANDOM}};
  btb_450_target_address = _RAND_1802[63:0];
  _RAND_1803 = {1{`RANDOM}};
  btb_450_bht = _RAND_1803[1:0];
  _RAND_1804 = {1{`RANDOM}};
  btb_451_valid = _RAND_1804[0:0];
  _RAND_1805 = {1{`RANDOM}};
  btb_451_tag = _RAND_1805[9:0];
  _RAND_1806 = {2{`RANDOM}};
  btb_451_target_address = _RAND_1806[63:0];
  _RAND_1807 = {1{`RANDOM}};
  btb_451_bht = _RAND_1807[1:0];
  _RAND_1808 = {1{`RANDOM}};
  btb_452_valid = _RAND_1808[0:0];
  _RAND_1809 = {1{`RANDOM}};
  btb_452_tag = _RAND_1809[9:0];
  _RAND_1810 = {2{`RANDOM}};
  btb_452_target_address = _RAND_1810[63:0];
  _RAND_1811 = {1{`RANDOM}};
  btb_452_bht = _RAND_1811[1:0];
  _RAND_1812 = {1{`RANDOM}};
  btb_453_valid = _RAND_1812[0:0];
  _RAND_1813 = {1{`RANDOM}};
  btb_453_tag = _RAND_1813[9:0];
  _RAND_1814 = {2{`RANDOM}};
  btb_453_target_address = _RAND_1814[63:0];
  _RAND_1815 = {1{`RANDOM}};
  btb_453_bht = _RAND_1815[1:0];
  _RAND_1816 = {1{`RANDOM}};
  btb_454_valid = _RAND_1816[0:0];
  _RAND_1817 = {1{`RANDOM}};
  btb_454_tag = _RAND_1817[9:0];
  _RAND_1818 = {2{`RANDOM}};
  btb_454_target_address = _RAND_1818[63:0];
  _RAND_1819 = {1{`RANDOM}};
  btb_454_bht = _RAND_1819[1:0];
  _RAND_1820 = {1{`RANDOM}};
  btb_455_valid = _RAND_1820[0:0];
  _RAND_1821 = {1{`RANDOM}};
  btb_455_tag = _RAND_1821[9:0];
  _RAND_1822 = {2{`RANDOM}};
  btb_455_target_address = _RAND_1822[63:0];
  _RAND_1823 = {1{`RANDOM}};
  btb_455_bht = _RAND_1823[1:0];
  _RAND_1824 = {1{`RANDOM}};
  btb_456_valid = _RAND_1824[0:0];
  _RAND_1825 = {1{`RANDOM}};
  btb_456_tag = _RAND_1825[9:0];
  _RAND_1826 = {2{`RANDOM}};
  btb_456_target_address = _RAND_1826[63:0];
  _RAND_1827 = {1{`RANDOM}};
  btb_456_bht = _RAND_1827[1:0];
  _RAND_1828 = {1{`RANDOM}};
  btb_457_valid = _RAND_1828[0:0];
  _RAND_1829 = {1{`RANDOM}};
  btb_457_tag = _RAND_1829[9:0];
  _RAND_1830 = {2{`RANDOM}};
  btb_457_target_address = _RAND_1830[63:0];
  _RAND_1831 = {1{`RANDOM}};
  btb_457_bht = _RAND_1831[1:0];
  _RAND_1832 = {1{`RANDOM}};
  btb_458_valid = _RAND_1832[0:0];
  _RAND_1833 = {1{`RANDOM}};
  btb_458_tag = _RAND_1833[9:0];
  _RAND_1834 = {2{`RANDOM}};
  btb_458_target_address = _RAND_1834[63:0];
  _RAND_1835 = {1{`RANDOM}};
  btb_458_bht = _RAND_1835[1:0];
  _RAND_1836 = {1{`RANDOM}};
  btb_459_valid = _RAND_1836[0:0];
  _RAND_1837 = {1{`RANDOM}};
  btb_459_tag = _RAND_1837[9:0];
  _RAND_1838 = {2{`RANDOM}};
  btb_459_target_address = _RAND_1838[63:0];
  _RAND_1839 = {1{`RANDOM}};
  btb_459_bht = _RAND_1839[1:0];
  _RAND_1840 = {1{`RANDOM}};
  btb_460_valid = _RAND_1840[0:0];
  _RAND_1841 = {1{`RANDOM}};
  btb_460_tag = _RAND_1841[9:0];
  _RAND_1842 = {2{`RANDOM}};
  btb_460_target_address = _RAND_1842[63:0];
  _RAND_1843 = {1{`RANDOM}};
  btb_460_bht = _RAND_1843[1:0];
  _RAND_1844 = {1{`RANDOM}};
  btb_461_valid = _RAND_1844[0:0];
  _RAND_1845 = {1{`RANDOM}};
  btb_461_tag = _RAND_1845[9:0];
  _RAND_1846 = {2{`RANDOM}};
  btb_461_target_address = _RAND_1846[63:0];
  _RAND_1847 = {1{`RANDOM}};
  btb_461_bht = _RAND_1847[1:0];
  _RAND_1848 = {1{`RANDOM}};
  btb_462_valid = _RAND_1848[0:0];
  _RAND_1849 = {1{`RANDOM}};
  btb_462_tag = _RAND_1849[9:0];
  _RAND_1850 = {2{`RANDOM}};
  btb_462_target_address = _RAND_1850[63:0];
  _RAND_1851 = {1{`RANDOM}};
  btb_462_bht = _RAND_1851[1:0];
  _RAND_1852 = {1{`RANDOM}};
  btb_463_valid = _RAND_1852[0:0];
  _RAND_1853 = {1{`RANDOM}};
  btb_463_tag = _RAND_1853[9:0];
  _RAND_1854 = {2{`RANDOM}};
  btb_463_target_address = _RAND_1854[63:0];
  _RAND_1855 = {1{`RANDOM}};
  btb_463_bht = _RAND_1855[1:0];
  _RAND_1856 = {1{`RANDOM}};
  btb_464_valid = _RAND_1856[0:0];
  _RAND_1857 = {1{`RANDOM}};
  btb_464_tag = _RAND_1857[9:0];
  _RAND_1858 = {2{`RANDOM}};
  btb_464_target_address = _RAND_1858[63:0];
  _RAND_1859 = {1{`RANDOM}};
  btb_464_bht = _RAND_1859[1:0];
  _RAND_1860 = {1{`RANDOM}};
  btb_465_valid = _RAND_1860[0:0];
  _RAND_1861 = {1{`RANDOM}};
  btb_465_tag = _RAND_1861[9:0];
  _RAND_1862 = {2{`RANDOM}};
  btb_465_target_address = _RAND_1862[63:0];
  _RAND_1863 = {1{`RANDOM}};
  btb_465_bht = _RAND_1863[1:0];
  _RAND_1864 = {1{`RANDOM}};
  btb_466_valid = _RAND_1864[0:0];
  _RAND_1865 = {1{`RANDOM}};
  btb_466_tag = _RAND_1865[9:0];
  _RAND_1866 = {2{`RANDOM}};
  btb_466_target_address = _RAND_1866[63:0];
  _RAND_1867 = {1{`RANDOM}};
  btb_466_bht = _RAND_1867[1:0];
  _RAND_1868 = {1{`RANDOM}};
  btb_467_valid = _RAND_1868[0:0];
  _RAND_1869 = {1{`RANDOM}};
  btb_467_tag = _RAND_1869[9:0];
  _RAND_1870 = {2{`RANDOM}};
  btb_467_target_address = _RAND_1870[63:0];
  _RAND_1871 = {1{`RANDOM}};
  btb_467_bht = _RAND_1871[1:0];
  _RAND_1872 = {1{`RANDOM}};
  btb_468_valid = _RAND_1872[0:0];
  _RAND_1873 = {1{`RANDOM}};
  btb_468_tag = _RAND_1873[9:0];
  _RAND_1874 = {2{`RANDOM}};
  btb_468_target_address = _RAND_1874[63:0];
  _RAND_1875 = {1{`RANDOM}};
  btb_468_bht = _RAND_1875[1:0];
  _RAND_1876 = {1{`RANDOM}};
  btb_469_valid = _RAND_1876[0:0];
  _RAND_1877 = {1{`RANDOM}};
  btb_469_tag = _RAND_1877[9:0];
  _RAND_1878 = {2{`RANDOM}};
  btb_469_target_address = _RAND_1878[63:0];
  _RAND_1879 = {1{`RANDOM}};
  btb_469_bht = _RAND_1879[1:0];
  _RAND_1880 = {1{`RANDOM}};
  btb_470_valid = _RAND_1880[0:0];
  _RAND_1881 = {1{`RANDOM}};
  btb_470_tag = _RAND_1881[9:0];
  _RAND_1882 = {2{`RANDOM}};
  btb_470_target_address = _RAND_1882[63:0];
  _RAND_1883 = {1{`RANDOM}};
  btb_470_bht = _RAND_1883[1:0];
  _RAND_1884 = {1{`RANDOM}};
  btb_471_valid = _RAND_1884[0:0];
  _RAND_1885 = {1{`RANDOM}};
  btb_471_tag = _RAND_1885[9:0];
  _RAND_1886 = {2{`RANDOM}};
  btb_471_target_address = _RAND_1886[63:0];
  _RAND_1887 = {1{`RANDOM}};
  btb_471_bht = _RAND_1887[1:0];
  _RAND_1888 = {1{`RANDOM}};
  btb_472_valid = _RAND_1888[0:0];
  _RAND_1889 = {1{`RANDOM}};
  btb_472_tag = _RAND_1889[9:0];
  _RAND_1890 = {2{`RANDOM}};
  btb_472_target_address = _RAND_1890[63:0];
  _RAND_1891 = {1{`RANDOM}};
  btb_472_bht = _RAND_1891[1:0];
  _RAND_1892 = {1{`RANDOM}};
  btb_473_valid = _RAND_1892[0:0];
  _RAND_1893 = {1{`RANDOM}};
  btb_473_tag = _RAND_1893[9:0];
  _RAND_1894 = {2{`RANDOM}};
  btb_473_target_address = _RAND_1894[63:0];
  _RAND_1895 = {1{`RANDOM}};
  btb_473_bht = _RAND_1895[1:0];
  _RAND_1896 = {1{`RANDOM}};
  btb_474_valid = _RAND_1896[0:0];
  _RAND_1897 = {1{`RANDOM}};
  btb_474_tag = _RAND_1897[9:0];
  _RAND_1898 = {2{`RANDOM}};
  btb_474_target_address = _RAND_1898[63:0];
  _RAND_1899 = {1{`RANDOM}};
  btb_474_bht = _RAND_1899[1:0];
  _RAND_1900 = {1{`RANDOM}};
  btb_475_valid = _RAND_1900[0:0];
  _RAND_1901 = {1{`RANDOM}};
  btb_475_tag = _RAND_1901[9:0];
  _RAND_1902 = {2{`RANDOM}};
  btb_475_target_address = _RAND_1902[63:0];
  _RAND_1903 = {1{`RANDOM}};
  btb_475_bht = _RAND_1903[1:0];
  _RAND_1904 = {1{`RANDOM}};
  btb_476_valid = _RAND_1904[0:0];
  _RAND_1905 = {1{`RANDOM}};
  btb_476_tag = _RAND_1905[9:0];
  _RAND_1906 = {2{`RANDOM}};
  btb_476_target_address = _RAND_1906[63:0];
  _RAND_1907 = {1{`RANDOM}};
  btb_476_bht = _RAND_1907[1:0];
  _RAND_1908 = {1{`RANDOM}};
  btb_477_valid = _RAND_1908[0:0];
  _RAND_1909 = {1{`RANDOM}};
  btb_477_tag = _RAND_1909[9:0];
  _RAND_1910 = {2{`RANDOM}};
  btb_477_target_address = _RAND_1910[63:0];
  _RAND_1911 = {1{`RANDOM}};
  btb_477_bht = _RAND_1911[1:0];
  _RAND_1912 = {1{`RANDOM}};
  btb_478_valid = _RAND_1912[0:0];
  _RAND_1913 = {1{`RANDOM}};
  btb_478_tag = _RAND_1913[9:0];
  _RAND_1914 = {2{`RANDOM}};
  btb_478_target_address = _RAND_1914[63:0];
  _RAND_1915 = {1{`RANDOM}};
  btb_478_bht = _RAND_1915[1:0];
  _RAND_1916 = {1{`RANDOM}};
  btb_479_valid = _RAND_1916[0:0];
  _RAND_1917 = {1{`RANDOM}};
  btb_479_tag = _RAND_1917[9:0];
  _RAND_1918 = {2{`RANDOM}};
  btb_479_target_address = _RAND_1918[63:0];
  _RAND_1919 = {1{`RANDOM}};
  btb_479_bht = _RAND_1919[1:0];
  _RAND_1920 = {1{`RANDOM}};
  btb_480_valid = _RAND_1920[0:0];
  _RAND_1921 = {1{`RANDOM}};
  btb_480_tag = _RAND_1921[9:0];
  _RAND_1922 = {2{`RANDOM}};
  btb_480_target_address = _RAND_1922[63:0];
  _RAND_1923 = {1{`RANDOM}};
  btb_480_bht = _RAND_1923[1:0];
  _RAND_1924 = {1{`RANDOM}};
  btb_481_valid = _RAND_1924[0:0];
  _RAND_1925 = {1{`RANDOM}};
  btb_481_tag = _RAND_1925[9:0];
  _RAND_1926 = {2{`RANDOM}};
  btb_481_target_address = _RAND_1926[63:0];
  _RAND_1927 = {1{`RANDOM}};
  btb_481_bht = _RAND_1927[1:0];
  _RAND_1928 = {1{`RANDOM}};
  btb_482_valid = _RAND_1928[0:0];
  _RAND_1929 = {1{`RANDOM}};
  btb_482_tag = _RAND_1929[9:0];
  _RAND_1930 = {2{`RANDOM}};
  btb_482_target_address = _RAND_1930[63:0];
  _RAND_1931 = {1{`RANDOM}};
  btb_482_bht = _RAND_1931[1:0];
  _RAND_1932 = {1{`RANDOM}};
  btb_483_valid = _RAND_1932[0:0];
  _RAND_1933 = {1{`RANDOM}};
  btb_483_tag = _RAND_1933[9:0];
  _RAND_1934 = {2{`RANDOM}};
  btb_483_target_address = _RAND_1934[63:0];
  _RAND_1935 = {1{`RANDOM}};
  btb_483_bht = _RAND_1935[1:0];
  _RAND_1936 = {1{`RANDOM}};
  btb_484_valid = _RAND_1936[0:0];
  _RAND_1937 = {1{`RANDOM}};
  btb_484_tag = _RAND_1937[9:0];
  _RAND_1938 = {2{`RANDOM}};
  btb_484_target_address = _RAND_1938[63:0];
  _RAND_1939 = {1{`RANDOM}};
  btb_484_bht = _RAND_1939[1:0];
  _RAND_1940 = {1{`RANDOM}};
  btb_485_valid = _RAND_1940[0:0];
  _RAND_1941 = {1{`RANDOM}};
  btb_485_tag = _RAND_1941[9:0];
  _RAND_1942 = {2{`RANDOM}};
  btb_485_target_address = _RAND_1942[63:0];
  _RAND_1943 = {1{`RANDOM}};
  btb_485_bht = _RAND_1943[1:0];
  _RAND_1944 = {1{`RANDOM}};
  btb_486_valid = _RAND_1944[0:0];
  _RAND_1945 = {1{`RANDOM}};
  btb_486_tag = _RAND_1945[9:0];
  _RAND_1946 = {2{`RANDOM}};
  btb_486_target_address = _RAND_1946[63:0];
  _RAND_1947 = {1{`RANDOM}};
  btb_486_bht = _RAND_1947[1:0];
  _RAND_1948 = {1{`RANDOM}};
  btb_487_valid = _RAND_1948[0:0];
  _RAND_1949 = {1{`RANDOM}};
  btb_487_tag = _RAND_1949[9:0];
  _RAND_1950 = {2{`RANDOM}};
  btb_487_target_address = _RAND_1950[63:0];
  _RAND_1951 = {1{`RANDOM}};
  btb_487_bht = _RAND_1951[1:0];
  _RAND_1952 = {1{`RANDOM}};
  btb_488_valid = _RAND_1952[0:0];
  _RAND_1953 = {1{`RANDOM}};
  btb_488_tag = _RAND_1953[9:0];
  _RAND_1954 = {2{`RANDOM}};
  btb_488_target_address = _RAND_1954[63:0];
  _RAND_1955 = {1{`RANDOM}};
  btb_488_bht = _RAND_1955[1:0];
  _RAND_1956 = {1{`RANDOM}};
  btb_489_valid = _RAND_1956[0:0];
  _RAND_1957 = {1{`RANDOM}};
  btb_489_tag = _RAND_1957[9:0];
  _RAND_1958 = {2{`RANDOM}};
  btb_489_target_address = _RAND_1958[63:0];
  _RAND_1959 = {1{`RANDOM}};
  btb_489_bht = _RAND_1959[1:0];
  _RAND_1960 = {1{`RANDOM}};
  btb_490_valid = _RAND_1960[0:0];
  _RAND_1961 = {1{`RANDOM}};
  btb_490_tag = _RAND_1961[9:0];
  _RAND_1962 = {2{`RANDOM}};
  btb_490_target_address = _RAND_1962[63:0];
  _RAND_1963 = {1{`RANDOM}};
  btb_490_bht = _RAND_1963[1:0];
  _RAND_1964 = {1{`RANDOM}};
  btb_491_valid = _RAND_1964[0:0];
  _RAND_1965 = {1{`RANDOM}};
  btb_491_tag = _RAND_1965[9:0];
  _RAND_1966 = {2{`RANDOM}};
  btb_491_target_address = _RAND_1966[63:0];
  _RAND_1967 = {1{`RANDOM}};
  btb_491_bht = _RAND_1967[1:0];
  _RAND_1968 = {1{`RANDOM}};
  btb_492_valid = _RAND_1968[0:0];
  _RAND_1969 = {1{`RANDOM}};
  btb_492_tag = _RAND_1969[9:0];
  _RAND_1970 = {2{`RANDOM}};
  btb_492_target_address = _RAND_1970[63:0];
  _RAND_1971 = {1{`RANDOM}};
  btb_492_bht = _RAND_1971[1:0];
  _RAND_1972 = {1{`RANDOM}};
  btb_493_valid = _RAND_1972[0:0];
  _RAND_1973 = {1{`RANDOM}};
  btb_493_tag = _RAND_1973[9:0];
  _RAND_1974 = {2{`RANDOM}};
  btb_493_target_address = _RAND_1974[63:0];
  _RAND_1975 = {1{`RANDOM}};
  btb_493_bht = _RAND_1975[1:0];
  _RAND_1976 = {1{`RANDOM}};
  btb_494_valid = _RAND_1976[0:0];
  _RAND_1977 = {1{`RANDOM}};
  btb_494_tag = _RAND_1977[9:0];
  _RAND_1978 = {2{`RANDOM}};
  btb_494_target_address = _RAND_1978[63:0];
  _RAND_1979 = {1{`RANDOM}};
  btb_494_bht = _RAND_1979[1:0];
  _RAND_1980 = {1{`RANDOM}};
  btb_495_valid = _RAND_1980[0:0];
  _RAND_1981 = {1{`RANDOM}};
  btb_495_tag = _RAND_1981[9:0];
  _RAND_1982 = {2{`RANDOM}};
  btb_495_target_address = _RAND_1982[63:0];
  _RAND_1983 = {1{`RANDOM}};
  btb_495_bht = _RAND_1983[1:0];
  _RAND_1984 = {1{`RANDOM}};
  btb_496_valid = _RAND_1984[0:0];
  _RAND_1985 = {1{`RANDOM}};
  btb_496_tag = _RAND_1985[9:0];
  _RAND_1986 = {2{`RANDOM}};
  btb_496_target_address = _RAND_1986[63:0];
  _RAND_1987 = {1{`RANDOM}};
  btb_496_bht = _RAND_1987[1:0];
  _RAND_1988 = {1{`RANDOM}};
  btb_497_valid = _RAND_1988[0:0];
  _RAND_1989 = {1{`RANDOM}};
  btb_497_tag = _RAND_1989[9:0];
  _RAND_1990 = {2{`RANDOM}};
  btb_497_target_address = _RAND_1990[63:0];
  _RAND_1991 = {1{`RANDOM}};
  btb_497_bht = _RAND_1991[1:0];
  _RAND_1992 = {1{`RANDOM}};
  btb_498_valid = _RAND_1992[0:0];
  _RAND_1993 = {1{`RANDOM}};
  btb_498_tag = _RAND_1993[9:0];
  _RAND_1994 = {2{`RANDOM}};
  btb_498_target_address = _RAND_1994[63:0];
  _RAND_1995 = {1{`RANDOM}};
  btb_498_bht = _RAND_1995[1:0];
  _RAND_1996 = {1{`RANDOM}};
  btb_499_valid = _RAND_1996[0:0];
  _RAND_1997 = {1{`RANDOM}};
  btb_499_tag = _RAND_1997[9:0];
  _RAND_1998 = {2{`RANDOM}};
  btb_499_target_address = _RAND_1998[63:0];
  _RAND_1999 = {1{`RANDOM}};
  btb_499_bht = _RAND_1999[1:0];
  _RAND_2000 = {1{`RANDOM}};
  btb_500_valid = _RAND_2000[0:0];
  _RAND_2001 = {1{`RANDOM}};
  btb_500_tag = _RAND_2001[9:0];
  _RAND_2002 = {2{`RANDOM}};
  btb_500_target_address = _RAND_2002[63:0];
  _RAND_2003 = {1{`RANDOM}};
  btb_500_bht = _RAND_2003[1:0];
  _RAND_2004 = {1{`RANDOM}};
  btb_501_valid = _RAND_2004[0:0];
  _RAND_2005 = {1{`RANDOM}};
  btb_501_tag = _RAND_2005[9:0];
  _RAND_2006 = {2{`RANDOM}};
  btb_501_target_address = _RAND_2006[63:0];
  _RAND_2007 = {1{`RANDOM}};
  btb_501_bht = _RAND_2007[1:0];
  _RAND_2008 = {1{`RANDOM}};
  btb_502_valid = _RAND_2008[0:0];
  _RAND_2009 = {1{`RANDOM}};
  btb_502_tag = _RAND_2009[9:0];
  _RAND_2010 = {2{`RANDOM}};
  btb_502_target_address = _RAND_2010[63:0];
  _RAND_2011 = {1{`RANDOM}};
  btb_502_bht = _RAND_2011[1:0];
  _RAND_2012 = {1{`RANDOM}};
  btb_503_valid = _RAND_2012[0:0];
  _RAND_2013 = {1{`RANDOM}};
  btb_503_tag = _RAND_2013[9:0];
  _RAND_2014 = {2{`RANDOM}};
  btb_503_target_address = _RAND_2014[63:0];
  _RAND_2015 = {1{`RANDOM}};
  btb_503_bht = _RAND_2015[1:0];
  _RAND_2016 = {1{`RANDOM}};
  btb_504_valid = _RAND_2016[0:0];
  _RAND_2017 = {1{`RANDOM}};
  btb_504_tag = _RAND_2017[9:0];
  _RAND_2018 = {2{`RANDOM}};
  btb_504_target_address = _RAND_2018[63:0];
  _RAND_2019 = {1{`RANDOM}};
  btb_504_bht = _RAND_2019[1:0];
  _RAND_2020 = {1{`RANDOM}};
  btb_505_valid = _RAND_2020[0:0];
  _RAND_2021 = {1{`RANDOM}};
  btb_505_tag = _RAND_2021[9:0];
  _RAND_2022 = {2{`RANDOM}};
  btb_505_target_address = _RAND_2022[63:0];
  _RAND_2023 = {1{`RANDOM}};
  btb_505_bht = _RAND_2023[1:0];
  _RAND_2024 = {1{`RANDOM}};
  btb_506_valid = _RAND_2024[0:0];
  _RAND_2025 = {1{`RANDOM}};
  btb_506_tag = _RAND_2025[9:0];
  _RAND_2026 = {2{`RANDOM}};
  btb_506_target_address = _RAND_2026[63:0];
  _RAND_2027 = {1{`RANDOM}};
  btb_506_bht = _RAND_2027[1:0];
  _RAND_2028 = {1{`RANDOM}};
  btb_507_valid = _RAND_2028[0:0];
  _RAND_2029 = {1{`RANDOM}};
  btb_507_tag = _RAND_2029[9:0];
  _RAND_2030 = {2{`RANDOM}};
  btb_507_target_address = _RAND_2030[63:0];
  _RAND_2031 = {1{`RANDOM}};
  btb_507_bht = _RAND_2031[1:0];
  _RAND_2032 = {1{`RANDOM}};
  btb_508_valid = _RAND_2032[0:0];
  _RAND_2033 = {1{`RANDOM}};
  btb_508_tag = _RAND_2033[9:0];
  _RAND_2034 = {2{`RANDOM}};
  btb_508_target_address = _RAND_2034[63:0];
  _RAND_2035 = {1{`RANDOM}};
  btb_508_bht = _RAND_2035[1:0];
  _RAND_2036 = {1{`RANDOM}};
  btb_509_valid = _RAND_2036[0:0];
  _RAND_2037 = {1{`RANDOM}};
  btb_509_tag = _RAND_2037[9:0];
  _RAND_2038 = {2{`RANDOM}};
  btb_509_target_address = _RAND_2038[63:0];
  _RAND_2039 = {1{`RANDOM}};
  btb_509_bht = _RAND_2039[1:0];
  _RAND_2040 = {1{`RANDOM}};
  btb_510_valid = _RAND_2040[0:0];
  _RAND_2041 = {1{`RANDOM}};
  btb_510_tag = _RAND_2041[9:0];
  _RAND_2042 = {2{`RANDOM}};
  btb_510_target_address = _RAND_2042[63:0];
  _RAND_2043 = {1{`RANDOM}};
  btb_510_bht = _RAND_2043[1:0];
  _RAND_2044 = {1{`RANDOM}};
  btb_511_valid = _RAND_2044[0:0];
  _RAND_2045 = {1{`RANDOM}};
  btb_511_tag = _RAND_2045[9:0];
  _RAND_2046 = {2{`RANDOM}};
  btb_511_target_address = _RAND_2046[63:0];
  _RAND_2047 = {1{`RANDOM}};
  btb_511_bht = _RAND_2047[1:0];
  _RAND_2048 = {1{`RANDOM}};
  btb_victim_ptr = _RAND_2048[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
